
  // General control and status                                                  
  input                                         sys__pe0__allSynchronized     ;
  output                                        pe0__sys__thisSynchronized    ;
  output                                        pe0__sys__ready               ;
  output                                        pe0__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe1__allSynchronized     ;
  output                                        pe1__sys__thisSynchronized    ;
  output                                        pe1__sys__ready               ;
  output                                        pe1__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe2__allSynchronized     ;
  output                                        pe2__sys__thisSynchronized    ;
  output                                        pe2__sys__ready               ;
  output                                        pe2__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe3__allSynchronized     ;
  output                                        pe3__sys__thisSynchronized    ;
  output                                        pe3__sys__ready               ;
  output                                        pe3__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe4__allSynchronized     ;
  output                                        pe4__sys__thisSynchronized    ;
  output                                        pe4__sys__ready               ;
  output                                        pe4__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe5__allSynchronized     ;
  output                                        pe5__sys__thisSynchronized    ;
  output                                        pe5__sys__ready               ;
  output                                        pe5__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe6__allSynchronized     ;
  output                                        pe6__sys__thisSynchronized    ;
  output                                        pe6__sys__ready               ;
  output                                        pe6__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe7__allSynchronized     ;
  output                                        pe7__sys__thisSynchronized    ;
  output                                        pe7__sys__ready               ;
  output                                        pe7__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe8__allSynchronized     ;
  output                                        pe8__sys__thisSynchronized    ;
  output                                        pe8__sys__ready               ;
  output                                        pe8__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe9__allSynchronized     ;
  output                                        pe9__sys__thisSynchronized    ;
  output                                        pe9__sys__ready               ;
  output                                        pe9__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe10__allSynchronized     ;
  output                                        pe10__sys__thisSynchronized    ;
  output                                        pe10__sys__ready               ;
  output                                        pe10__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe11__allSynchronized     ;
  output                                        pe11__sys__thisSynchronized    ;
  output                                        pe11__sys__ready               ;
  output                                        pe11__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe12__allSynchronized     ;
  output                                        pe12__sys__thisSynchronized    ;
  output                                        pe12__sys__ready               ;
  output                                        pe12__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe13__allSynchronized     ;
  output                                        pe13__sys__thisSynchronized    ;
  output                                        pe13__sys__ready               ;
  output                                        pe13__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe14__allSynchronized     ;
  output                                        pe14__sys__thisSynchronized    ;
  output                                        pe14__sys__ready               ;
  output                                        pe14__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe15__allSynchronized     ;
  output                                        pe15__sys__thisSynchronized    ;
  output                                        pe15__sys__ready               ;
  output                                        pe15__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe16__allSynchronized     ;
  output                                        pe16__sys__thisSynchronized    ;
  output                                        pe16__sys__ready               ;
  output                                        pe16__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe17__allSynchronized     ;
  output                                        pe17__sys__thisSynchronized    ;
  output                                        pe17__sys__ready               ;
  output                                        pe17__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe18__allSynchronized     ;
  output                                        pe18__sys__thisSynchronized    ;
  output                                        pe18__sys__ready               ;
  output                                        pe18__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe19__allSynchronized     ;
  output                                        pe19__sys__thisSynchronized    ;
  output                                        pe19__sys__ready               ;
  output                                        pe19__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe20__allSynchronized     ;
  output                                        pe20__sys__thisSynchronized    ;
  output                                        pe20__sys__ready               ;
  output                                        pe20__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe21__allSynchronized     ;
  output                                        pe21__sys__thisSynchronized    ;
  output                                        pe21__sys__ready               ;
  output                                        pe21__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe22__allSynchronized     ;
  output                                        pe22__sys__thisSynchronized    ;
  output                                        pe22__sys__ready               ;
  output                                        pe22__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe23__allSynchronized     ;
  output                                        pe23__sys__thisSynchronized    ;
  output                                        pe23__sys__ready               ;
  output                                        pe23__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe24__allSynchronized     ;
  output                                        pe24__sys__thisSynchronized    ;
  output                                        pe24__sys__ready               ;
  output                                        pe24__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe25__allSynchronized     ;
  output                                        pe25__sys__thisSynchronized    ;
  output                                        pe25__sys__ready               ;
  output                                        pe25__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe26__allSynchronized     ;
  output                                        pe26__sys__thisSynchronized    ;
  output                                        pe26__sys__ready               ;
  output                                        pe26__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe27__allSynchronized     ;
  output                                        pe27__sys__thisSynchronized    ;
  output                                        pe27__sys__ready               ;
  output                                        pe27__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe28__allSynchronized     ;
  output                                        pe28__sys__thisSynchronized    ;
  output                                        pe28__sys__ready               ;
  output                                        pe28__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe29__allSynchronized     ;
  output                                        pe29__sys__thisSynchronized    ;
  output                                        pe29__sys__ready               ;
  output                                        pe29__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe30__allSynchronized     ;
  output                                        pe30__sys__thisSynchronized    ;
  output                                        pe30__sys__ready               ;
  output                                        pe30__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe31__allSynchronized     ;
  output                                        pe31__sys__thisSynchronized    ;
  output                                        pe31__sys__ready               ;
  output                                        pe31__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe32__allSynchronized     ;
  output                                        pe32__sys__thisSynchronized    ;
  output                                        pe32__sys__ready               ;
  output                                        pe32__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe33__allSynchronized     ;
  output                                        pe33__sys__thisSynchronized    ;
  output                                        pe33__sys__ready               ;
  output                                        pe33__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe34__allSynchronized     ;
  output                                        pe34__sys__thisSynchronized    ;
  output                                        pe34__sys__ready               ;
  output                                        pe34__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe35__allSynchronized     ;
  output                                        pe35__sys__thisSynchronized    ;
  output                                        pe35__sys__ready               ;
  output                                        pe35__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe36__allSynchronized     ;
  output                                        pe36__sys__thisSynchronized    ;
  output                                        pe36__sys__ready               ;
  output                                        pe36__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe37__allSynchronized     ;
  output                                        pe37__sys__thisSynchronized    ;
  output                                        pe37__sys__ready               ;
  output                                        pe37__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe38__allSynchronized     ;
  output                                        pe38__sys__thisSynchronized    ;
  output                                        pe38__sys__ready               ;
  output                                        pe38__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe39__allSynchronized     ;
  output                                        pe39__sys__thisSynchronized    ;
  output                                        pe39__sys__ready               ;
  output                                        pe39__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe40__allSynchronized     ;
  output                                        pe40__sys__thisSynchronized    ;
  output                                        pe40__sys__ready               ;
  output                                        pe40__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe41__allSynchronized     ;
  output                                        pe41__sys__thisSynchronized    ;
  output                                        pe41__sys__ready               ;
  output                                        pe41__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe42__allSynchronized     ;
  output                                        pe42__sys__thisSynchronized    ;
  output                                        pe42__sys__ready               ;
  output                                        pe42__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe43__allSynchronized     ;
  output                                        pe43__sys__thisSynchronized    ;
  output                                        pe43__sys__ready               ;
  output                                        pe43__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe44__allSynchronized     ;
  output                                        pe44__sys__thisSynchronized    ;
  output                                        pe44__sys__ready               ;
  output                                        pe44__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe45__allSynchronized     ;
  output                                        pe45__sys__thisSynchronized    ;
  output                                        pe45__sys__ready               ;
  output                                        pe45__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe46__allSynchronized     ;
  output                                        pe46__sys__thisSynchronized    ;
  output                                        pe46__sys__ready               ;
  output                                        pe46__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe47__allSynchronized     ;
  output                                        pe47__sys__thisSynchronized    ;
  output                                        pe47__sys__ready               ;
  output                                        pe47__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe48__allSynchronized     ;
  output                                        pe48__sys__thisSynchronized    ;
  output                                        pe48__sys__ready               ;
  output                                        pe48__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe49__allSynchronized     ;
  output                                        pe49__sys__thisSynchronized    ;
  output                                        pe49__sys__ready               ;
  output                                        pe49__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe50__allSynchronized     ;
  output                                        pe50__sys__thisSynchronized    ;
  output                                        pe50__sys__ready               ;
  output                                        pe50__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe51__allSynchronized     ;
  output                                        pe51__sys__thisSynchronized    ;
  output                                        pe51__sys__ready               ;
  output                                        pe51__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe52__allSynchronized     ;
  output                                        pe52__sys__thisSynchronized    ;
  output                                        pe52__sys__ready               ;
  output                                        pe52__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe53__allSynchronized     ;
  output                                        pe53__sys__thisSynchronized    ;
  output                                        pe53__sys__ready               ;
  output                                        pe53__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe54__allSynchronized     ;
  output                                        pe54__sys__thisSynchronized    ;
  output                                        pe54__sys__ready               ;
  output                                        pe54__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe55__allSynchronized     ;
  output                                        pe55__sys__thisSynchronized    ;
  output                                        pe55__sys__ready               ;
  output                                        pe55__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe56__allSynchronized     ;
  output                                        pe56__sys__thisSynchronized    ;
  output                                        pe56__sys__ready               ;
  output                                        pe56__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe57__allSynchronized     ;
  output                                        pe57__sys__thisSynchronized    ;
  output                                        pe57__sys__ready               ;
  output                                        pe57__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe58__allSynchronized     ;
  output                                        pe58__sys__thisSynchronized    ;
  output                                        pe58__sys__ready               ;
  output                                        pe58__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe59__allSynchronized     ;
  output                                        pe59__sys__thisSynchronized    ;
  output                                        pe59__sys__ready               ;
  output                                        pe59__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe60__allSynchronized     ;
  output                                        pe60__sys__thisSynchronized    ;
  output                                        pe60__sys__ready               ;
  output                                        pe60__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe61__allSynchronized     ;
  output                                        pe61__sys__thisSynchronized    ;
  output                                        pe61__sys__ready               ;
  output                                        pe61__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe62__allSynchronized     ;
  output                                        pe62__sys__thisSynchronized    ;
  output                                        pe62__sys__ready               ;
  output                                        pe62__sys__complete            ;
  // General control and status                                                  
  input                                         sys__pe63__allSynchronized     ;
  output                                        pe63__sys__thisSynchronized    ;
  output                                        pe63__sys__ready               ;
  output                                        pe63__sys__complete            ;