
  // General control and status                                                   
  output                                        mgr0__sys__allSynchronized     ;
  input                                         sys__mgr0__thisSynchronized    ;
  input                                         sys__mgr0__ready               ;
  input                                         sys__mgr0__complete            ;
  // General control and status                                                   
  output                                        mgr1__sys__allSynchronized     ;
  input                                         sys__mgr1__thisSynchronized    ;
  input                                         sys__mgr1__ready               ;
  input                                         sys__mgr1__complete            ;
  // General control and status                                                   
  output                                        mgr2__sys__allSynchronized     ;
  input                                         sys__mgr2__thisSynchronized    ;
  input                                         sys__mgr2__ready               ;
  input                                         sys__mgr2__complete            ;
  // General control and status                                                   
  output                                        mgr3__sys__allSynchronized     ;
  input                                         sys__mgr3__thisSynchronized    ;
  input                                         sys__mgr3__ready               ;
  input                                         sys__mgr3__complete            ;