
    // Lane 0                 
    std__pe0__lane0_strm0_cntl        = 'd0         ;
    std__pe0__lane0_strm0_data        = 'h1234_5678 ;
    std__pe0__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe0__lane0_strm1_cntl        = 'd0         ;
    std__pe0__lane0_strm1_data        = 'h1234_5678 ;
    std__pe0__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe0__lane1_strm0_cntl        = 'd0         ;
    std__pe0__lane1_strm0_data        = 'h1234_5678 ;
    std__pe0__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe0__lane1_strm1_cntl        = 'd0         ;
    std__pe0__lane1_strm1_data        = 'h1234_5678 ;
    std__pe0__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe0__lane2_strm0_cntl        = 'd0         ;
    std__pe0__lane2_strm0_data        = 'h1234_5678 ;
    std__pe0__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe0__lane2_strm1_cntl        = 'd0         ;
    std__pe0__lane2_strm1_data        = 'h1234_5678 ;
    std__pe0__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe0__lane3_strm0_cntl        = 'd0         ;
    std__pe0__lane3_strm0_data        = 'h1234_5678 ;
    std__pe0__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe0__lane3_strm1_cntl        = 'd0         ;
    std__pe0__lane3_strm1_data        = 'h1234_5678 ;
    std__pe0__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe0__lane4_strm0_cntl        = 'd0         ;
    std__pe0__lane4_strm0_data        = 'h1234_5678 ;
    std__pe0__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe0__lane4_strm1_cntl        = 'd0         ;
    std__pe0__lane4_strm1_data        = 'h1234_5678 ;
    std__pe0__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe0__lane5_strm0_cntl        = 'd0         ;
    std__pe0__lane5_strm0_data        = 'h1234_5678 ;
    std__pe0__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe0__lane5_strm1_cntl        = 'd0         ;
    std__pe0__lane5_strm1_data        = 'h1234_5678 ;
    std__pe0__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe0__lane6_strm0_cntl        = 'd0         ;
    std__pe0__lane6_strm0_data        = 'h1234_5678 ;
    std__pe0__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe0__lane6_strm1_cntl        = 'd0         ;
    std__pe0__lane6_strm1_data        = 'h1234_5678 ;
    std__pe0__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe0__lane7_strm0_cntl        = 'd0         ;
    std__pe0__lane7_strm0_data        = 'h1234_5678 ;
    std__pe0__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe0__lane7_strm1_cntl        = 'd0         ;
    std__pe0__lane7_strm1_data        = 'h1234_5678 ;
    std__pe0__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe0__lane8_strm0_cntl        = 'd0         ;
    std__pe0__lane8_strm0_data        = 'h1234_5678 ;
    std__pe0__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe0__lane8_strm1_cntl        = 'd0         ;
    std__pe0__lane8_strm1_data        = 'h1234_5678 ;
    std__pe0__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe0__lane9_strm0_cntl        = 'd0         ;
    std__pe0__lane9_strm0_data        = 'h1234_5678 ;
    std__pe0__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe0__lane9_strm1_cntl        = 'd0         ;
    std__pe0__lane9_strm1_data        = 'h1234_5678 ;
    std__pe0__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe0__lane10_strm0_cntl        = 'd0         ;
    std__pe0__lane10_strm0_data        = 'h1234_5678 ;
    std__pe0__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe0__lane10_strm1_cntl        = 'd0         ;
    std__pe0__lane10_strm1_data        = 'h1234_5678 ;
    std__pe0__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe0__lane11_strm0_cntl        = 'd0         ;
    std__pe0__lane11_strm0_data        = 'h1234_5678 ;
    std__pe0__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe0__lane11_strm1_cntl        = 'd0         ;
    std__pe0__lane11_strm1_data        = 'h1234_5678 ;
    std__pe0__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe0__lane12_strm0_cntl        = 'd0         ;
    std__pe0__lane12_strm0_data        = 'h1234_5678 ;
    std__pe0__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe0__lane12_strm1_cntl        = 'd0         ;
    std__pe0__lane12_strm1_data        = 'h1234_5678 ;
    std__pe0__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe0__lane13_strm0_cntl        = 'd0         ;
    std__pe0__lane13_strm0_data        = 'h1234_5678 ;
    std__pe0__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe0__lane13_strm1_cntl        = 'd0         ;
    std__pe0__lane13_strm1_data        = 'h1234_5678 ;
    std__pe0__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe0__lane14_strm0_cntl        = 'd0         ;
    std__pe0__lane14_strm0_data        = 'h1234_5678 ;
    std__pe0__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe0__lane14_strm1_cntl        = 'd0         ;
    std__pe0__lane14_strm1_data        = 'h1234_5678 ;
    std__pe0__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe0__lane15_strm0_cntl        = 'd0         ;
    std__pe0__lane15_strm0_data        = 'h1234_5678 ;
    std__pe0__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe0__lane15_strm1_cntl        = 'd0         ;
    std__pe0__lane15_strm1_data        = 'h1234_5678 ;
    std__pe0__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe0__lane16_strm0_cntl        = 'd0         ;
    std__pe0__lane16_strm0_data        = 'h1234_5678 ;
    std__pe0__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe0__lane16_strm1_cntl        = 'd0         ;
    std__pe0__lane16_strm1_data        = 'h1234_5678 ;
    std__pe0__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe0__lane17_strm0_cntl        = 'd0         ;
    std__pe0__lane17_strm0_data        = 'h1234_5678 ;
    std__pe0__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe0__lane17_strm1_cntl        = 'd0         ;
    std__pe0__lane17_strm1_data        = 'h1234_5678 ;
    std__pe0__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe0__lane18_strm0_cntl        = 'd0         ;
    std__pe0__lane18_strm0_data        = 'h1234_5678 ;
    std__pe0__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe0__lane18_strm1_cntl        = 'd0         ;
    std__pe0__lane18_strm1_data        = 'h1234_5678 ;
    std__pe0__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe0__lane19_strm0_cntl        = 'd0         ;
    std__pe0__lane19_strm0_data        = 'h1234_5678 ;
    std__pe0__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe0__lane19_strm1_cntl        = 'd0         ;
    std__pe0__lane19_strm1_data        = 'h1234_5678 ;
    std__pe0__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe0__lane20_strm0_cntl        = 'd0         ;
    std__pe0__lane20_strm0_data        = 'h1234_5678 ;
    std__pe0__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe0__lane20_strm1_cntl        = 'd0         ;
    std__pe0__lane20_strm1_data        = 'h1234_5678 ;
    std__pe0__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe0__lane21_strm0_cntl        = 'd0         ;
    std__pe0__lane21_strm0_data        = 'h1234_5678 ;
    std__pe0__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe0__lane21_strm1_cntl        = 'd0         ;
    std__pe0__lane21_strm1_data        = 'h1234_5678 ;
    std__pe0__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe0__lane22_strm0_cntl        = 'd0         ;
    std__pe0__lane22_strm0_data        = 'h1234_5678 ;
    std__pe0__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe0__lane22_strm1_cntl        = 'd0         ;
    std__pe0__lane22_strm1_data        = 'h1234_5678 ;
    std__pe0__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe0__lane23_strm0_cntl        = 'd0         ;
    std__pe0__lane23_strm0_data        = 'h1234_5678 ;
    std__pe0__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe0__lane23_strm1_cntl        = 'd0         ;
    std__pe0__lane23_strm1_data        = 'h1234_5678 ;
    std__pe0__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe0__lane24_strm0_cntl        = 'd0         ;
    std__pe0__lane24_strm0_data        = 'h1234_5678 ;
    std__pe0__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe0__lane24_strm1_cntl        = 'd0         ;
    std__pe0__lane24_strm1_data        = 'h1234_5678 ;
    std__pe0__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe0__lane25_strm0_cntl        = 'd0         ;
    std__pe0__lane25_strm0_data        = 'h1234_5678 ;
    std__pe0__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe0__lane25_strm1_cntl        = 'd0         ;
    std__pe0__lane25_strm1_data        = 'h1234_5678 ;
    std__pe0__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe0__lane26_strm0_cntl        = 'd0         ;
    std__pe0__lane26_strm0_data        = 'h1234_5678 ;
    std__pe0__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe0__lane26_strm1_cntl        = 'd0         ;
    std__pe0__lane26_strm1_data        = 'h1234_5678 ;
    std__pe0__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe0__lane27_strm0_cntl        = 'd0         ;
    std__pe0__lane27_strm0_data        = 'h1234_5678 ;
    std__pe0__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe0__lane27_strm1_cntl        = 'd0         ;
    std__pe0__lane27_strm1_data        = 'h1234_5678 ;
    std__pe0__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe0__lane28_strm0_cntl        = 'd0         ;
    std__pe0__lane28_strm0_data        = 'h1234_5678 ;
    std__pe0__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe0__lane28_strm1_cntl        = 'd0         ;
    std__pe0__lane28_strm1_data        = 'h1234_5678 ;
    std__pe0__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe0__lane29_strm0_cntl        = 'd0         ;
    std__pe0__lane29_strm0_data        = 'h1234_5678 ;
    std__pe0__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe0__lane29_strm1_cntl        = 'd0         ;
    std__pe0__lane29_strm1_data        = 'h1234_5678 ;
    std__pe0__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe0__lane30_strm0_cntl        = 'd0         ;
    std__pe0__lane30_strm0_data        = 'h1234_5678 ;
    std__pe0__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe0__lane30_strm1_cntl        = 'd0         ;
    std__pe0__lane30_strm1_data        = 'h1234_5678 ;
    std__pe0__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe0__lane31_strm0_cntl        = 'd0         ;
    std__pe0__lane31_strm0_data        = 'h1234_5678 ;
    std__pe0__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe0__lane31_strm1_cntl        = 'd0         ;
    std__pe0__lane31_strm1_data        = 'h1234_5678 ;
    std__pe0__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe1__lane0_strm0_cntl        = 'd0         ;
    std__pe1__lane0_strm0_data        = 'h1234_5678 ;
    std__pe1__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe1__lane0_strm1_cntl        = 'd0         ;
    std__pe1__lane0_strm1_data        = 'h1234_5678 ;
    std__pe1__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe1__lane1_strm0_cntl        = 'd0         ;
    std__pe1__lane1_strm0_data        = 'h1234_5678 ;
    std__pe1__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe1__lane1_strm1_cntl        = 'd0         ;
    std__pe1__lane1_strm1_data        = 'h1234_5678 ;
    std__pe1__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe1__lane2_strm0_cntl        = 'd0         ;
    std__pe1__lane2_strm0_data        = 'h1234_5678 ;
    std__pe1__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe1__lane2_strm1_cntl        = 'd0         ;
    std__pe1__lane2_strm1_data        = 'h1234_5678 ;
    std__pe1__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe1__lane3_strm0_cntl        = 'd0         ;
    std__pe1__lane3_strm0_data        = 'h1234_5678 ;
    std__pe1__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe1__lane3_strm1_cntl        = 'd0         ;
    std__pe1__lane3_strm1_data        = 'h1234_5678 ;
    std__pe1__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe1__lane4_strm0_cntl        = 'd0         ;
    std__pe1__lane4_strm0_data        = 'h1234_5678 ;
    std__pe1__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe1__lane4_strm1_cntl        = 'd0         ;
    std__pe1__lane4_strm1_data        = 'h1234_5678 ;
    std__pe1__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe1__lane5_strm0_cntl        = 'd0         ;
    std__pe1__lane5_strm0_data        = 'h1234_5678 ;
    std__pe1__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe1__lane5_strm1_cntl        = 'd0         ;
    std__pe1__lane5_strm1_data        = 'h1234_5678 ;
    std__pe1__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe1__lane6_strm0_cntl        = 'd0         ;
    std__pe1__lane6_strm0_data        = 'h1234_5678 ;
    std__pe1__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe1__lane6_strm1_cntl        = 'd0         ;
    std__pe1__lane6_strm1_data        = 'h1234_5678 ;
    std__pe1__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe1__lane7_strm0_cntl        = 'd0         ;
    std__pe1__lane7_strm0_data        = 'h1234_5678 ;
    std__pe1__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe1__lane7_strm1_cntl        = 'd0         ;
    std__pe1__lane7_strm1_data        = 'h1234_5678 ;
    std__pe1__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe1__lane8_strm0_cntl        = 'd0         ;
    std__pe1__lane8_strm0_data        = 'h1234_5678 ;
    std__pe1__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe1__lane8_strm1_cntl        = 'd0         ;
    std__pe1__lane8_strm1_data        = 'h1234_5678 ;
    std__pe1__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe1__lane9_strm0_cntl        = 'd0         ;
    std__pe1__lane9_strm0_data        = 'h1234_5678 ;
    std__pe1__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe1__lane9_strm1_cntl        = 'd0         ;
    std__pe1__lane9_strm1_data        = 'h1234_5678 ;
    std__pe1__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe1__lane10_strm0_cntl        = 'd0         ;
    std__pe1__lane10_strm0_data        = 'h1234_5678 ;
    std__pe1__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe1__lane10_strm1_cntl        = 'd0         ;
    std__pe1__lane10_strm1_data        = 'h1234_5678 ;
    std__pe1__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe1__lane11_strm0_cntl        = 'd0         ;
    std__pe1__lane11_strm0_data        = 'h1234_5678 ;
    std__pe1__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe1__lane11_strm1_cntl        = 'd0         ;
    std__pe1__lane11_strm1_data        = 'h1234_5678 ;
    std__pe1__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe1__lane12_strm0_cntl        = 'd0         ;
    std__pe1__lane12_strm0_data        = 'h1234_5678 ;
    std__pe1__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe1__lane12_strm1_cntl        = 'd0         ;
    std__pe1__lane12_strm1_data        = 'h1234_5678 ;
    std__pe1__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe1__lane13_strm0_cntl        = 'd0         ;
    std__pe1__lane13_strm0_data        = 'h1234_5678 ;
    std__pe1__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe1__lane13_strm1_cntl        = 'd0         ;
    std__pe1__lane13_strm1_data        = 'h1234_5678 ;
    std__pe1__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe1__lane14_strm0_cntl        = 'd0         ;
    std__pe1__lane14_strm0_data        = 'h1234_5678 ;
    std__pe1__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe1__lane14_strm1_cntl        = 'd0         ;
    std__pe1__lane14_strm1_data        = 'h1234_5678 ;
    std__pe1__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe1__lane15_strm0_cntl        = 'd0         ;
    std__pe1__lane15_strm0_data        = 'h1234_5678 ;
    std__pe1__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe1__lane15_strm1_cntl        = 'd0         ;
    std__pe1__lane15_strm1_data        = 'h1234_5678 ;
    std__pe1__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe1__lane16_strm0_cntl        = 'd0         ;
    std__pe1__lane16_strm0_data        = 'h1234_5678 ;
    std__pe1__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe1__lane16_strm1_cntl        = 'd0         ;
    std__pe1__lane16_strm1_data        = 'h1234_5678 ;
    std__pe1__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe1__lane17_strm0_cntl        = 'd0         ;
    std__pe1__lane17_strm0_data        = 'h1234_5678 ;
    std__pe1__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe1__lane17_strm1_cntl        = 'd0         ;
    std__pe1__lane17_strm1_data        = 'h1234_5678 ;
    std__pe1__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe1__lane18_strm0_cntl        = 'd0         ;
    std__pe1__lane18_strm0_data        = 'h1234_5678 ;
    std__pe1__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe1__lane18_strm1_cntl        = 'd0         ;
    std__pe1__lane18_strm1_data        = 'h1234_5678 ;
    std__pe1__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe1__lane19_strm0_cntl        = 'd0         ;
    std__pe1__lane19_strm0_data        = 'h1234_5678 ;
    std__pe1__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe1__lane19_strm1_cntl        = 'd0         ;
    std__pe1__lane19_strm1_data        = 'h1234_5678 ;
    std__pe1__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe1__lane20_strm0_cntl        = 'd0         ;
    std__pe1__lane20_strm0_data        = 'h1234_5678 ;
    std__pe1__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe1__lane20_strm1_cntl        = 'd0         ;
    std__pe1__lane20_strm1_data        = 'h1234_5678 ;
    std__pe1__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe1__lane21_strm0_cntl        = 'd0         ;
    std__pe1__lane21_strm0_data        = 'h1234_5678 ;
    std__pe1__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe1__lane21_strm1_cntl        = 'd0         ;
    std__pe1__lane21_strm1_data        = 'h1234_5678 ;
    std__pe1__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe1__lane22_strm0_cntl        = 'd0         ;
    std__pe1__lane22_strm0_data        = 'h1234_5678 ;
    std__pe1__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe1__lane22_strm1_cntl        = 'd0         ;
    std__pe1__lane22_strm1_data        = 'h1234_5678 ;
    std__pe1__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe1__lane23_strm0_cntl        = 'd0         ;
    std__pe1__lane23_strm0_data        = 'h1234_5678 ;
    std__pe1__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe1__lane23_strm1_cntl        = 'd0         ;
    std__pe1__lane23_strm1_data        = 'h1234_5678 ;
    std__pe1__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe1__lane24_strm0_cntl        = 'd0         ;
    std__pe1__lane24_strm0_data        = 'h1234_5678 ;
    std__pe1__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe1__lane24_strm1_cntl        = 'd0         ;
    std__pe1__lane24_strm1_data        = 'h1234_5678 ;
    std__pe1__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe1__lane25_strm0_cntl        = 'd0         ;
    std__pe1__lane25_strm0_data        = 'h1234_5678 ;
    std__pe1__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe1__lane25_strm1_cntl        = 'd0         ;
    std__pe1__lane25_strm1_data        = 'h1234_5678 ;
    std__pe1__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe1__lane26_strm0_cntl        = 'd0         ;
    std__pe1__lane26_strm0_data        = 'h1234_5678 ;
    std__pe1__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe1__lane26_strm1_cntl        = 'd0         ;
    std__pe1__lane26_strm1_data        = 'h1234_5678 ;
    std__pe1__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe1__lane27_strm0_cntl        = 'd0         ;
    std__pe1__lane27_strm0_data        = 'h1234_5678 ;
    std__pe1__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe1__lane27_strm1_cntl        = 'd0         ;
    std__pe1__lane27_strm1_data        = 'h1234_5678 ;
    std__pe1__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe1__lane28_strm0_cntl        = 'd0         ;
    std__pe1__lane28_strm0_data        = 'h1234_5678 ;
    std__pe1__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe1__lane28_strm1_cntl        = 'd0         ;
    std__pe1__lane28_strm1_data        = 'h1234_5678 ;
    std__pe1__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe1__lane29_strm0_cntl        = 'd0         ;
    std__pe1__lane29_strm0_data        = 'h1234_5678 ;
    std__pe1__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe1__lane29_strm1_cntl        = 'd0         ;
    std__pe1__lane29_strm1_data        = 'h1234_5678 ;
    std__pe1__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe1__lane30_strm0_cntl        = 'd0         ;
    std__pe1__lane30_strm0_data        = 'h1234_5678 ;
    std__pe1__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe1__lane30_strm1_cntl        = 'd0         ;
    std__pe1__lane30_strm1_data        = 'h1234_5678 ;
    std__pe1__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe1__lane31_strm0_cntl        = 'd0         ;
    std__pe1__lane31_strm0_data        = 'h1234_5678 ;
    std__pe1__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe1__lane31_strm1_cntl        = 'd0         ;
    std__pe1__lane31_strm1_data        = 'h1234_5678 ;
    std__pe1__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe2__lane0_strm0_cntl        = 'd0         ;
    std__pe2__lane0_strm0_data        = 'h1234_5678 ;
    std__pe2__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe2__lane0_strm1_cntl        = 'd0         ;
    std__pe2__lane0_strm1_data        = 'h1234_5678 ;
    std__pe2__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe2__lane1_strm0_cntl        = 'd0         ;
    std__pe2__lane1_strm0_data        = 'h1234_5678 ;
    std__pe2__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe2__lane1_strm1_cntl        = 'd0         ;
    std__pe2__lane1_strm1_data        = 'h1234_5678 ;
    std__pe2__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe2__lane2_strm0_cntl        = 'd0         ;
    std__pe2__lane2_strm0_data        = 'h1234_5678 ;
    std__pe2__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe2__lane2_strm1_cntl        = 'd0         ;
    std__pe2__lane2_strm1_data        = 'h1234_5678 ;
    std__pe2__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe2__lane3_strm0_cntl        = 'd0         ;
    std__pe2__lane3_strm0_data        = 'h1234_5678 ;
    std__pe2__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe2__lane3_strm1_cntl        = 'd0         ;
    std__pe2__lane3_strm1_data        = 'h1234_5678 ;
    std__pe2__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe2__lane4_strm0_cntl        = 'd0         ;
    std__pe2__lane4_strm0_data        = 'h1234_5678 ;
    std__pe2__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe2__lane4_strm1_cntl        = 'd0         ;
    std__pe2__lane4_strm1_data        = 'h1234_5678 ;
    std__pe2__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe2__lane5_strm0_cntl        = 'd0         ;
    std__pe2__lane5_strm0_data        = 'h1234_5678 ;
    std__pe2__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe2__lane5_strm1_cntl        = 'd0         ;
    std__pe2__lane5_strm1_data        = 'h1234_5678 ;
    std__pe2__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe2__lane6_strm0_cntl        = 'd0         ;
    std__pe2__lane6_strm0_data        = 'h1234_5678 ;
    std__pe2__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe2__lane6_strm1_cntl        = 'd0         ;
    std__pe2__lane6_strm1_data        = 'h1234_5678 ;
    std__pe2__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe2__lane7_strm0_cntl        = 'd0         ;
    std__pe2__lane7_strm0_data        = 'h1234_5678 ;
    std__pe2__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe2__lane7_strm1_cntl        = 'd0         ;
    std__pe2__lane7_strm1_data        = 'h1234_5678 ;
    std__pe2__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe2__lane8_strm0_cntl        = 'd0         ;
    std__pe2__lane8_strm0_data        = 'h1234_5678 ;
    std__pe2__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe2__lane8_strm1_cntl        = 'd0         ;
    std__pe2__lane8_strm1_data        = 'h1234_5678 ;
    std__pe2__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe2__lane9_strm0_cntl        = 'd0         ;
    std__pe2__lane9_strm0_data        = 'h1234_5678 ;
    std__pe2__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe2__lane9_strm1_cntl        = 'd0         ;
    std__pe2__lane9_strm1_data        = 'h1234_5678 ;
    std__pe2__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe2__lane10_strm0_cntl        = 'd0         ;
    std__pe2__lane10_strm0_data        = 'h1234_5678 ;
    std__pe2__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe2__lane10_strm1_cntl        = 'd0         ;
    std__pe2__lane10_strm1_data        = 'h1234_5678 ;
    std__pe2__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe2__lane11_strm0_cntl        = 'd0         ;
    std__pe2__lane11_strm0_data        = 'h1234_5678 ;
    std__pe2__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe2__lane11_strm1_cntl        = 'd0         ;
    std__pe2__lane11_strm1_data        = 'h1234_5678 ;
    std__pe2__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe2__lane12_strm0_cntl        = 'd0         ;
    std__pe2__lane12_strm0_data        = 'h1234_5678 ;
    std__pe2__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe2__lane12_strm1_cntl        = 'd0         ;
    std__pe2__lane12_strm1_data        = 'h1234_5678 ;
    std__pe2__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe2__lane13_strm0_cntl        = 'd0         ;
    std__pe2__lane13_strm0_data        = 'h1234_5678 ;
    std__pe2__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe2__lane13_strm1_cntl        = 'd0         ;
    std__pe2__lane13_strm1_data        = 'h1234_5678 ;
    std__pe2__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe2__lane14_strm0_cntl        = 'd0         ;
    std__pe2__lane14_strm0_data        = 'h1234_5678 ;
    std__pe2__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe2__lane14_strm1_cntl        = 'd0         ;
    std__pe2__lane14_strm1_data        = 'h1234_5678 ;
    std__pe2__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe2__lane15_strm0_cntl        = 'd0         ;
    std__pe2__lane15_strm0_data        = 'h1234_5678 ;
    std__pe2__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe2__lane15_strm1_cntl        = 'd0         ;
    std__pe2__lane15_strm1_data        = 'h1234_5678 ;
    std__pe2__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe2__lane16_strm0_cntl        = 'd0         ;
    std__pe2__lane16_strm0_data        = 'h1234_5678 ;
    std__pe2__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe2__lane16_strm1_cntl        = 'd0         ;
    std__pe2__lane16_strm1_data        = 'h1234_5678 ;
    std__pe2__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe2__lane17_strm0_cntl        = 'd0         ;
    std__pe2__lane17_strm0_data        = 'h1234_5678 ;
    std__pe2__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe2__lane17_strm1_cntl        = 'd0         ;
    std__pe2__lane17_strm1_data        = 'h1234_5678 ;
    std__pe2__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe2__lane18_strm0_cntl        = 'd0         ;
    std__pe2__lane18_strm0_data        = 'h1234_5678 ;
    std__pe2__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe2__lane18_strm1_cntl        = 'd0         ;
    std__pe2__lane18_strm1_data        = 'h1234_5678 ;
    std__pe2__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe2__lane19_strm0_cntl        = 'd0         ;
    std__pe2__lane19_strm0_data        = 'h1234_5678 ;
    std__pe2__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe2__lane19_strm1_cntl        = 'd0         ;
    std__pe2__lane19_strm1_data        = 'h1234_5678 ;
    std__pe2__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe2__lane20_strm0_cntl        = 'd0         ;
    std__pe2__lane20_strm0_data        = 'h1234_5678 ;
    std__pe2__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe2__lane20_strm1_cntl        = 'd0         ;
    std__pe2__lane20_strm1_data        = 'h1234_5678 ;
    std__pe2__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe2__lane21_strm0_cntl        = 'd0         ;
    std__pe2__lane21_strm0_data        = 'h1234_5678 ;
    std__pe2__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe2__lane21_strm1_cntl        = 'd0         ;
    std__pe2__lane21_strm1_data        = 'h1234_5678 ;
    std__pe2__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe2__lane22_strm0_cntl        = 'd0         ;
    std__pe2__lane22_strm0_data        = 'h1234_5678 ;
    std__pe2__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe2__lane22_strm1_cntl        = 'd0         ;
    std__pe2__lane22_strm1_data        = 'h1234_5678 ;
    std__pe2__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe2__lane23_strm0_cntl        = 'd0         ;
    std__pe2__lane23_strm0_data        = 'h1234_5678 ;
    std__pe2__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe2__lane23_strm1_cntl        = 'd0         ;
    std__pe2__lane23_strm1_data        = 'h1234_5678 ;
    std__pe2__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe2__lane24_strm0_cntl        = 'd0         ;
    std__pe2__lane24_strm0_data        = 'h1234_5678 ;
    std__pe2__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe2__lane24_strm1_cntl        = 'd0         ;
    std__pe2__lane24_strm1_data        = 'h1234_5678 ;
    std__pe2__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe2__lane25_strm0_cntl        = 'd0         ;
    std__pe2__lane25_strm0_data        = 'h1234_5678 ;
    std__pe2__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe2__lane25_strm1_cntl        = 'd0         ;
    std__pe2__lane25_strm1_data        = 'h1234_5678 ;
    std__pe2__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe2__lane26_strm0_cntl        = 'd0         ;
    std__pe2__lane26_strm0_data        = 'h1234_5678 ;
    std__pe2__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe2__lane26_strm1_cntl        = 'd0         ;
    std__pe2__lane26_strm1_data        = 'h1234_5678 ;
    std__pe2__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe2__lane27_strm0_cntl        = 'd0         ;
    std__pe2__lane27_strm0_data        = 'h1234_5678 ;
    std__pe2__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe2__lane27_strm1_cntl        = 'd0         ;
    std__pe2__lane27_strm1_data        = 'h1234_5678 ;
    std__pe2__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe2__lane28_strm0_cntl        = 'd0         ;
    std__pe2__lane28_strm0_data        = 'h1234_5678 ;
    std__pe2__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe2__lane28_strm1_cntl        = 'd0         ;
    std__pe2__lane28_strm1_data        = 'h1234_5678 ;
    std__pe2__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe2__lane29_strm0_cntl        = 'd0         ;
    std__pe2__lane29_strm0_data        = 'h1234_5678 ;
    std__pe2__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe2__lane29_strm1_cntl        = 'd0         ;
    std__pe2__lane29_strm1_data        = 'h1234_5678 ;
    std__pe2__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe2__lane30_strm0_cntl        = 'd0         ;
    std__pe2__lane30_strm0_data        = 'h1234_5678 ;
    std__pe2__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe2__lane30_strm1_cntl        = 'd0         ;
    std__pe2__lane30_strm1_data        = 'h1234_5678 ;
    std__pe2__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe2__lane31_strm0_cntl        = 'd0         ;
    std__pe2__lane31_strm0_data        = 'h1234_5678 ;
    std__pe2__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe2__lane31_strm1_cntl        = 'd0         ;
    std__pe2__lane31_strm1_data        = 'h1234_5678 ;
    std__pe2__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe3__lane0_strm0_cntl        = 'd0         ;
    std__pe3__lane0_strm0_data        = 'h1234_5678 ;
    std__pe3__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe3__lane0_strm1_cntl        = 'd0         ;
    std__pe3__lane0_strm1_data        = 'h1234_5678 ;
    std__pe3__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe3__lane1_strm0_cntl        = 'd0         ;
    std__pe3__lane1_strm0_data        = 'h1234_5678 ;
    std__pe3__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe3__lane1_strm1_cntl        = 'd0         ;
    std__pe3__lane1_strm1_data        = 'h1234_5678 ;
    std__pe3__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe3__lane2_strm0_cntl        = 'd0         ;
    std__pe3__lane2_strm0_data        = 'h1234_5678 ;
    std__pe3__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe3__lane2_strm1_cntl        = 'd0         ;
    std__pe3__lane2_strm1_data        = 'h1234_5678 ;
    std__pe3__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe3__lane3_strm0_cntl        = 'd0         ;
    std__pe3__lane3_strm0_data        = 'h1234_5678 ;
    std__pe3__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe3__lane3_strm1_cntl        = 'd0         ;
    std__pe3__lane3_strm1_data        = 'h1234_5678 ;
    std__pe3__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe3__lane4_strm0_cntl        = 'd0         ;
    std__pe3__lane4_strm0_data        = 'h1234_5678 ;
    std__pe3__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe3__lane4_strm1_cntl        = 'd0         ;
    std__pe3__lane4_strm1_data        = 'h1234_5678 ;
    std__pe3__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe3__lane5_strm0_cntl        = 'd0         ;
    std__pe3__lane5_strm0_data        = 'h1234_5678 ;
    std__pe3__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe3__lane5_strm1_cntl        = 'd0         ;
    std__pe3__lane5_strm1_data        = 'h1234_5678 ;
    std__pe3__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe3__lane6_strm0_cntl        = 'd0         ;
    std__pe3__lane6_strm0_data        = 'h1234_5678 ;
    std__pe3__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe3__lane6_strm1_cntl        = 'd0         ;
    std__pe3__lane6_strm1_data        = 'h1234_5678 ;
    std__pe3__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe3__lane7_strm0_cntl        = 'd0         ;
    std__pe3__lane7_strm0_data        = 'h1234_5678 ;
    std__pe3__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe3__lane7_strm1_cntl        = 'd0         ;
    std__pe3__lane7_strm1_data        = 'h1234_5678 ;
    std__pe3__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe3__lane8_strm0_cntl        = 'd0         ;
    std__pe3__lane8_strm0_data        = 'h1234_5678 ;
    std__pe3__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe3__lane8_strm1_cntl        = 'd0         ;
    std__pe3__lane8_strm1_data        = 'h1234_5678 ;
    std__pe3__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe3__lane9_strm0_cntl        = 'd0         ;
    std__pe3__lane9_strm0_data        = 'h1234_5678 ;
    std__pe3__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe3__lane9_strm1_cntl        = 'd0         ;
    std__pe3__lane9_strm1_data        = 'h1234_5678 ;
    std__pe3__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe3__lane10_strm0_cntl        = 'd0         ;
    std__pe3__lane10_strm0_data        = 'h1234_5678 ;
    std__pe3__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe3__lane10_strm1_cntl        = 'd0         ;
    std__pe3__lane10_strm1_data        = 'h1234_5678 ;
    std__pe3__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe3__lane11_strm0_cntl        = 'd0         ;
    std__pe3__lane11_strm0_data        = 'h1234_5678 ;
    std__pe3__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe3__lane11_strm1_cntl        = 'd0         ;
    std__pe3__lane11_strm1_data        = 'h1234_5678 ;
    std__pe3__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe3__lane12_strm0_cntl        = 'd0         ;
    std__pe3__lane12_strm0_data        = 'h1234_5678 ;
    std__pe3__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe3__lane12_strm1_cntl        = 'd0         ;
    std__pe3__lane12_strm1_data        = 'h1234_5678 ;
    std__pe3__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe3__lane13_strm0_cntl        = 'd0         ;
    std__pe3__lane13_strm0_data        = 'h1234_5678 ;
    std__pe3__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe3__lane13_strm1_cntl        = 'd0         ;
    std__pe3__lane13_strm1_data        = 'h1234_5678 ;
    std__pe3__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe3__lane14_strm0_cntl        = 'd0         ;
    std__pe3__lane14_strm0_data        = 'h1234_5678 ;
    std__pe3__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe3__lane14_strm1_cntl        = 'd0         ;
    std__pe3__lane14_strm1_data        = 'h1234_5678 ;
    std__pe3__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe3__lane15_strm0_cntl        = 'd0         ;
    std__pe3__lane15_strm0_data        = 'h1234_5678 ;
    std__pe3__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe3__lane15_strm1_cntl        = 'd0         ;
    std__pe3__lane15_strm1_data        = 'h1234_5678 ;
    std__pe3__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe3__lane16_strm0_cntl        = 'd0         ;
    std__pe3__lane16_strm0_data        = 'h1234_5678 ;
    std__pe3__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe3__lane16_strm1_cntl        = 'd0         ;
    std__pe3__lane16_strm1_data        = 'h1234_5678 ;
    std__pe3__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe3__lane17_strm0_cntl        = 'd0         ;
    std__pe3__lane17_strm0_data        = 'h1234_5678 ;
    std__pe3__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe3__lane17_strm1_cntl        = 'd0         ;
    std__pe3__lane17_strm1_data        = 'h1234_5678 ;
    std__pe3__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe3__lane18_strm0_cntl        = 'd0         ;
    std__pe3__lane18_strm0_data        = 'h1234_5678 ;
    std__pe3__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe3__lane18_strm1_cntl        = 'd0         ;
    std__pe3__lane18_strm1_data        = 'h1234_5678 ;
    std__pe3__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe3__lane19_strm0_cntl        = 'd0         ;
    std__pe3__lane19_strm0_data        = 'h1234_5678 ;
    std__pe3__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe3__lane19_strm1_cntl        = 'd0         ;
    std__pe3__lane19_strm1_data        = 'h1234_5678 ;
    std__pe3__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe3__lane20_strm0_cntl        = 'd0         ;
    std__pe3__lane20_strm0_data        = 'h1234_5678 ;
    std__pe3__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe3__lane20_strm1_cntl        = 'd0         ;
    std__pe3__lane20_strm1_data        = 'h1234_5678 ;
    std__pe3__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe3__lane21_strm0_cntl        = 'd0         ;
    std__pe3__lane21_strm0_data        = 'h1234_5678 ;
    std__pe3__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe3__lane21_strm1_cntl        = 'd0         ;
    std__pe3__lane21_strm1_data        = 'h1234_5678 ;
    std__pe3__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe3__lane22_strm0_cntl        = 'd0         ;
    std__pe3__lane22_strm0_data        = 'h1234_5678 ;
    std__pe3__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe3__lane22_strm1_cntl        = 'd0         ;
    std__pe3__lane22_strm1_data        = 'h1234_5678 ;
    std__pe3__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe3__lane23_strm0_cntl        = 'd0         ;
    std__pe3__lane23_strm0_data        = 'h1234_5678 ;
    std__pe3__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe3__lane23_strm1_cntl        = 'd0         ;
    std__pe3__lane23_strm1_data        = 'h1234_5678 ;
    std__pe3__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe3__lane24_strm0_cntl        = 'd0         ;
    std__pe3__lane24_strm0_data        = 'h1234_5678 ;
    std__pe3__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe3__lane24_strm1_cntl        = 'd0         ;
    std__pe3__lane24_strm1_data        = 'h1234_5678 ;
    std__pe3__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe3__lane25_strm0_cntl        = 'd0         ;
    std__pe3__lane25_strm0_data        = 'h1234_5678 ;
    std__pe3__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe3__lane25_strm1_cntl        = 'd0         ;
    std__pe3__lane25_strm1_data        = 'h1234_5678 ;
    std__pe3__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe3__lane26_strm0_cntl        = 'd0         ;
    std__pe3__lane26_strm0_data        = 'h1234_5678 ;
    std__pe3__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe3__lane26_strm1_cntl        = 'd0         ;
    std__pe3__lane26_strm1_data        = 'h1234_5678 ;
    std__pe3__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe3__lane27_strm0_cntl        = 'd0         ;
    std__pe3__lane27_strm0_data        = 'h1234_5678 ;
    std__pe3__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe3__lane27_strm1_cntl        = 'd0         ;
    std__pe3__lane27_strm1_data        = 'h1234_5678 ;
    std__pe3__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe3__lane28_strm0_cntl        = 'd0         ;
    std__pe3__lane28_strm0_data        = 'h1234_5678 ;
    std__pe3__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe3__lane28_strm1_cntl        = 'd0         ;
    std__pe3__lane28_strm1_data        = 'h1234_5678 ;
    std__pe3__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe3__lane29_strm0_cntl        = 'd0         ;
    std__pe3__lane29_strm0_data        = 'h1234_5678 ;
    std__pe3__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe3__lane29_strm1_cntl        = 'd0         ;
    std__pe3__lane29_strm1_data        = 'h1234_5678 ;
    std__pe3__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe3__lane30_strm0_cntl        = 'd0         ;
    std__pe3__lane30_strm0_data        = 'h1234_5678 ;
    std__pe3__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe3__lane30_strm1_cntl        = 'd0         ;
    std__pe3__lane30_strm1_data        = 'h1234_5678 ;
    std__pe3__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe3__lane31_strm0_cntl        = 'd0         ;
    std__pe3__lane31_strm0_data        = 'h1234_5678 ;
    std__pe3__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe3__lane31_strm1_cntl        = 'd0         ;
    std__pe3__lane31_strm1_data        = 'h1234_5678 ;
    std__pe3__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe4__lane0_strm0_cntl        = 'd0         ;
    std__pe4__lane0_strm0_data        = 'h1234_5678 ;
    std__pe4__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe4__lane0_strm1_cntl        = 'd0         ;
    std__pe4__lane0_strm1_data        = 'h1234_5678 ;
    std__pe4__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe4__lane1_strm0_cntl        = 'd0         ;
    std__pe4__lane1_strm0_data        = 'h1234_5678 ;
    std__pe4__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe4__lane1_strm1_cntl        = 'd0         ;
    std__pe4__lane1_strm1_data        = 'h1234_5678 ;
    std__pe4__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe4__lane2_strm0_cntl        = 'd0         ;
    std__pe4__lane2_strm0_data        = 'h1234_5678 ;
    std__pe4__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe4__lane2_strm1_cntl        = 'd0         ;
    std__pe4__lane2_strm1_data        = 'h1234_5678 ;
    std__pe4__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe4__lane3_strm0_cntl        = 'd0         ;
    std__pe4__lane3_strm0_data        = 'h1234_5678 ;
    std__pe4__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe4__lane3_strm1_cntl        = 'd0         ;
    std__pe4__lane3_strm1_data        = 'h1234_5678 ;
    std__pe4__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe4__lane4_strm0_cntl        = 'd0         ;
    std__pe4__lane4_strm0_data        = 'h1234_5678 ;
    std__pe4__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe4__lane4_strm1_cntl        = 'd0         ;
    std__pe4__lane4_strm1_data        = 'h1234_5678 ;
    std__pe4__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe4__lane5_strm0_cntl        = 'd0         ;
    std__pe4__lane5_strm0_data        = 'h1234_5678 ;
    std__pe4__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe4__lane5_strm1_cntl        = 'd0         ;
    std__pe4__lane5_strm1_data        = 'h1234_5678 ;
    std__pe4__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe4__lane6_strm0_cntl        = 'd0         ;
    std__pe4__lane6_strm0_data        = 'h1234_5678 ;
    std__pe4__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe4__lane6_strm1_cntl        = 'd0         ;
    std__pe4__lane6_strm1_data        = 'h1234_5678 ;
    std__pe4__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe4__lane7_strm0_cntl        = 'd0         ;
    std__pe4__lane7_strm0_data        = 'h1234_5678 ;
    std__pe4__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe4__lane7_strm1_cntl        = 'd0         ;
    std__pe4__lane7_strm1_data        = 'h1234_5678 ;
    std__pe4__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe4__lane8_strm0_cntl        = 'd0         ;
    std__pe4__lane8_strm0_data        = 'h1234_5678 ;
    std__pe4__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe4__lane8_strm1_cntl        = 'd0         ;
    std__pe4__lane8_strm1_data        = 'h1234_5678 ;
    std__pe4__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe4__lane9_strm0_cntl        = 'd0         ;
    std__pe4__lane9_strm0_data        = 'h1234_5678 ;
    std__pe4__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe4__lane9_strm1_cntl        = 'd0         ;
    std__pe4__lane9_strm1_data        = 'h1234_5678 ;
    std__pe4__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe4__lane10_strm0_cntl        = 'd0         ;
    std__pe4__lane10_strm0_data        = 'h1234_5678 ;
    std__pe4__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe4__lane10_strm1_cntl        = 'd0         ;
    std__pe4__lane10_strm1_data        = 'h1234_5678 ;
    std__pe4__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe4__lane11_strm0_cntl        = 'd0         ;
    std__pe4__lane11_strm0_data        = 'h1234_5678 ;
    std__pe4__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe4__lane11_strm1_cntl        = 'd0         ;
    std__pe4__lane11_strm1_data        = 'h1234_5678 ;
    std__pe4__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe4__lane12_strm0_cntl        = 'd0         ;
    std__pe4__lane12_strm0_data        = 'h1234_5678 ;
    std__pe4__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe4__lane12_strm1_cntl        = 'd0         ;
    std__pe4__lane12_strm1_data        = 'h1234_5678 ;
    std__pe4__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe4__lane13_strm0_cntl        = 'd0         ;
    std__pe4__lane13_strm0_data        = 'h1234_5678 ;
    std__pe4__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe4__lane13_strm1_cntl        = 'd0         ;
    std__pe4__lane13_strm1_data        = 'h1234_5678 ;
    std__pe4__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe4__lane14_strm0_cntl        = 'd0         ;
    std__pe4__lane14_strm0_data        = 'h1234_5678 ;
    std__pe4__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe4__lane14_strm1_cntl        = 'd0         ;
    std__pe4__lane14_strm1_data        = 'h1234_5678 ;
    std__pe4__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe4__lane15_strm0_cntl        = 'd0         ;
    std__pe4__lane15_strm0_data        = 'h1234_5678 ;
    std__pe4__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe4__lane15_strm1_cntl        = 'd0         ;
    std__pe4__lane15_strm1_data        = 'h1234_5678 ;
    std__pe4__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe4__lane16_strm0_cntl        = 'd0         ;
    std__pe4__lane16_strm0_data        = 'h1234_5678 ;
    std__pe4__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe4__lane16_strm1_cntl        = 'd0         ;
    std__pe4__lane16_strm1_data        = 'h1234_5678 ;
    std__pe4__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe4__lane17_strm0_cntl        = 'd0         ;
    std__pe4__lane17_strm0_data        = 'h1234_5678 ;
    std__pe4__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe4__lane17_strm1_cntl        = 'd0         ;
    std__pe4__lane17_strm1_data        = 'h1234_5678 ;
    std__pe4__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe4__lane18_strm0_cntl        = 'd0         ;
    std__pe4__lane18_strm0_data        = 'h1234_5678 ;
    std__pe4__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe4__lane18_strm1_cntl        = 'd0         ;
    std__pe4__lane18_strm1_data        = 'h1234_5678 ;
    std__pe4__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe4__lane19_strm0_cntl        = 'd0         ;
    std__pe4__lane19_strm0_data        = 'h1234_5678 ;
    std__pe4__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe4__lane19_strm1_cntl        = 'd0         ;
    std__pe4__lane19_strm1_data        = 'h1234_5678 ;
    std__pe4__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe4__lane20_strm0_cntl        = 'd0         ;
    std__pe4__lane20_strm0_data        = 'h1234_5678 ;
    std__pe4__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe4__lane20_strm1_cntl        = 'd0         ;
    std__pe4__lane20_strm1_data        = 'h1234_5678 ;
    std__pe4__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe4__lane21_strm0_cntl        = 'd0         ;
    std__pe4__lane21_strm0_data        = 'h1234_5678 ;
    std__pe4__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe4__lane21_strm1_cntl        = 'd0         ;
    std__pe4__lane21_strm1_data        = 'h1234_5678 ;
    std__pe4__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe4__lane22_strm0_cntl        = 'd0         ;
    std__pe4__lane22_strm0_data        = 'h1234_5678 ;
    std__pe4__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe4__lane22_strm1_cntl        = 'd0         ;
    std__pe4__lane22_strm1_data        = 'h1234_5678 ;
    std__pe4__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe4__lane23_strm0_cntl        = 'd0         ;
    std__pe4__lane23_strm0_data        = 'h1234_5678 ;
    std__pe4__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe4__lane23_strm1_cntl        = 'd0         ;
    std__pe4__lane23_strm1_data        = 'h1234_5678 ;
    std__pe4__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe4__lane24_strm0_cntl        = 'd0         ;
    std__pe4__lane24_strm0_data        = 'h1234_5678 ;
    std__pe4__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe4__lane24_strm1_cntl        = 'd0         ;
    std__pe4__lane24_strm1_data        = 'h1234_5678 ;
    std__pe4__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe4__lane25_strm0_cntl        = 'd0         ;
    std__pe4__lane25_strm0_data        = 'h1234_5678 ;
    std__pe4__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe4__lane25_strm1_cntl        = 'd0         ;
    std__pe4__lane25_strm1_data        = 'h1234_5678 ;
    std__pe4__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe4__lane26_strm0_cntl        = 'd0         ;
    std__pe4__lane26_strm0_data        = 'h1234_5678 ;
    std__pe4__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe4__lane26_strm1_cntl        = 'd0         ;
    std__pe4__lane26_strm1_data        = 'h1234_5678 ;
    std__pe4__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe4__lane27_strm0_cntl        = 'd0         ;
    std__pe4__lane27_strm0_data        = 'h1234_5678 ;
    std__pe4__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe4__lane27_strm1_cntl        = 'd0         ;
    std__pe4__lane27_strm1_data        = 'h1234_5678 ;
    std__pe4__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe4__lane28_strm0_cntl        = 'd0         ;
    std__pe4__lane28_strm0_data        = 'h1234_5678 ;
    std__pe4__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe4__lane28_strm1_cntl        = 'd0         ;
    std__pe4__lane28_strm1_data        = 'h1234_5678 ;
    std__pe4__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe4__lane29_strm0_cntl        = 'd0         ;
    std__pe4__lane29_strm0_data        = 'h1234_5678 ;
    std__pe4__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe4__lane29_strm1_cntl        = 'd0         ;
    std__pe4__lane29_strm1_data        = 'h1234_5678 ;
    std__pe4__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe4__lane30_strm0_cntl        = 'd0         ;
    std__pe4__lane30_strm0_data        = 'h1234_5678 ;
    std__pe4__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe4__lane30_strm1_cntl        = 'd0         ;
    std__pe4__lane30_strm1_data        = 'h1234_5678 ;
    std__pe4__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe4__lane31_strm0_cntl        = 'd0         ;
    std__pe4__lane31_strm0_data        = 'h1234_5678 ;
    std__pe4__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe4__lane31_strm1_cntl        = 'd0         ;
    std__pe4__lane31_strm1_data        = 'h1234_5678 ;
    std__pe4__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe5__lane0_strm0_cntl        = 'd0         ;
    std__pe5__lane0_strm0_data        = 'h1234_5678 ;
    std__pe5__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe5__lane0_strm1_cntl        = 'd0         ;
    std__pe5__lane0_strm1_data        = 'h1234_5678 ;
    std__pe5__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe5__lane1_strm0_cntl        = 'd0         ;
    std__pe5__lane1_strm0_data        = 'h1234_5678 ;
    std__pe5__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe5__lane1_strm1_cntl        = 'd0         ;
    std__pe5__lane1_strm1_data        = 'h1234_5678 ;
    std__pe5__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe5__lane2_strm0_cntl        = 'd0         ;
    std__pe5__lane2_strm0_data        = 'h1234_5678 ;
    std__pe5__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe5__lane2_strm1_cntl        = 'd0         ;
    std__pe5__lane2_strm1_data        = 'h1234_5678 ;
    std__pe5__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe5__lane3_strm0_cntl        = 'd0         ;
    std__pe5__lane3_strm0_data        = 'h1234_5678 ;
    std__pe5__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe5__lane3_strm1_cntl        = 'd0         ;
    std__pe5__lane3_strm1_data        = 'h1234_5678 ;
    std__pe5__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe5__lane4_strm0_cntl        = 'd0         ;
    std__pe5__lane4_strm0_data        = 'h1234_5678 ;
    std__pe5__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe5__lane4_strm1_cntl        = 'd0         ;
    std__pe5__lane4_strm1_data        = 'h1234_5678 ;
    std__pe5__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe5__lane5_strm0_cntl        = 'd0         ;
    std__pe5__lane5_strm0_data        = 'h1234_5678 ;
    std__pe5__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe5__lane5_strm1_cntl        = 'd0         ;
    std__pe5__lane5_strm1_data        = 'h1234_5678 ;
    std__pe5__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe5__lane6_strm0_cntl        = 'd0         ;
    std__pe5__lane6_strm0_data        = 'h1234_5678 ;
    std__pe5__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe5__lane6_strm1_cntl        = 'd0         ;
    std__pe5__lane6_strm1_data        = 'h1234_5678 ;
    std__pe5__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe5__lane7_strm0_cntl        = 'd0         ;
    std__pe5__lane7_strm0_data        = 'h1234_5678 ;
    std__pe5__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe5__lane7_strm1_cntl        = 'd0         ;
    std__pe5__lane7_strm1_data        = 'h1234_5678 ;
    std__pe5__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe5__lane8_strm0_cntl        = 'd0         ;
    std__pe5__lane8_strm0_data        = 'h1234_5678 ;
    std__pe5__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe5__lane8_strm1_cntl        = 'd0         ;
    std__pe5__lane8_strm1_data        = 'h1234_5678 ;
    std__pe5__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe5__lane9_strm0_cntl        = 'd0         ;
    std__pe5__lane9_strm0_data        = 'h1234_5678 ;
    std__pe5__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe5__lane9_strm1_cntl        = 'd0         ;
    std__pe5__lane9_strm1_data        = 'h1234_5678 ;
    std__pe5__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe5__lane10_strm0_cntl        = 'd0         ;
    std__pe5__lane10_strm0_data        = 'h1234_5678 ;
    std__pe5__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe5__lane10_strm1_cntl        = 'd0         ;
    std__pe5__lane10_strm1_data        = 'h1234_5678 ;
    std__pe5__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe5__lane11_strm0_cntl        = 'd0         ;
    std__pe5__lane11_strm0_data        = 'h1234_5678 ;
    std__pe5__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe5__lane11_strm1_cntl        = 'd0         ;
    std__pe5__lane11_strm1_data        = 'h1234_5678 ;
    std__pe5__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe5__lane12_strm0_cntl        = 'd0         ;
    std__pe5__lane12_strm0_data        = 'h1234_5678 ;
    std__pe5__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe5__lane12_strm1_cntl        = 'd0         ;
    std__pe5__lane12_strm1_data        = 'h1234_5678 ;
    std__pe5__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe5__lane13_strm0_cntl        = 'd0         ;
    std__pe5__lane13_strm0_data        = 'h1234_5678 ;
    std__pe5__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe5__lane13_strm1_cntl        = 'd0         ;
    std__pe5__lane13_strm1_data        = 'h1234_5678 ;
    std__pe5__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe5__lane14_strm0_cntl        = 'd0         ;
    std__pe5__lane14_strm0_data        = 'h1234_5678 ;
    std__pe5__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe5__lane14_strm1_cntl        = 'd0         ;
    std__pe5__lane14_strm1_data        = 'h1234_5678 ;
    std__pe5__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe5__lane15_strm0_cntl        = 'd0         ;
    std__pe5__lane15_strm0_data        = 'h1234_5678 ;
    std__pe5__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe5__lane15_strm1_cntl        = 'd0         ;
    std__pe5__lane15_strm1_data        = 'h1234_5678 ;
    std__pe5__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe5__lane16_strm0_cntl        = 'd0         ;
    std__pe5__lane16_strm0_data        = 'h1234_5678 ;
    std__pe5__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe5__lane16_strm1_cntl        = 'd0         ;
    std__pe5__lane16_strm1_data        = 'h1234_5678 ;
    std__pe5__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe5__lane17_strm0_cntl        = 'd0         ;
    std__pe5__lane17_strm0_data        = 'h1234_5678 ;
    std__pe5__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe5__lane17_strm1_cntl        = 'd0         ;
    std__pe5__lane17_strm1_data        = 'h1234_5678 ;
    std__pe5__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe5__lane18_strm0_cntl        = 'd0         ;
    std__pe5__lane18_strm0_data        = 'h1234_5678 ;
    std__pe5__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe5__lane18_strm1_cntl        = 'd0         ;
    std__pe5__lane18_strm1_data        = 'h1234_5678 ;
    std__pe5__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe5__lane19_strm0_cntl        = 'd0         ;
    std__pe5__lane19_strm0_data        = 'h1234_5678 ;
    std__pe5__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe5__lane19_strm1_cntl        = 'd0         ;
    std__pe5__lane19_strm1_data        = 'h1234_5678 ;
    std__pe5__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe5__lane20_strm0_cntl        = 'd0         ;
    std__pe5__lane20_strm0_data        = 'h1234_5678 ;
    std__pe5__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe5__lane20_strm1_cntl        = 'd0         ;
    std__pe5__lane20_strm1_data        = 'h1234_5678 ;
    std__pe5__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe5__lane21_strm0_cntl        = 'd0         ;
    std__pe5__lane21_strm0_data        = 'h1234_5678 ;
    std__pe5__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe5__lane21_strm1_cntl        = 'd0         ;
    std__pe5__lane21_strm1_data        = 'h1234_5678 ;
    std__pe5__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe5__lane22_strm0_cntl        = 'd0         ;
    std__pe5__lane22_strm0_data        = 'h1234_5678 ;
    std__pe5__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe5__lane22_strm1_cntl        = 'd0         ;
    std__pe5__lane22_strm1_data        = 'h1234_5678 ;
    std__pe5__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe5__lane23_strm0_cntl        = 'd0         ;
    std__pe5__lane23_strm0_data        = 'h1234_5678 ;
    std__pe5__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe5__lane23_strm1_cntl        = 'd0         ;
    std__pe5__lane23_strm1_data        = 'h1234_5678 ;
    std__pe5__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe5__lane24_strm0_cntl        = 'd0         ;
    std__pe5__lane24_strm0_data        = 'h1234_5678 ;
    std__pe5__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe5__lane24_strm1_cntl        = 'd0         ;
    std__pe5__lane24_strm1_data        = 'h1234_5678 ;
    std__pe5__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe5__lane25_strm0_cntl        = 'd0         ;
    std__pe5__lane25_strm0_data        = 'h1234_5678 ;
    std__pe5__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe5__lane25_strm1_cntl        = 'd0         ;
    std__pe5__lane25_strm1_data        = 'h1234_5678 ;
    std__pe5__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe5__lane26_strm0_cntl        = 'd0         ;
    std__pe5__lane26_strm0_data        = 'h1234_5678 ;
    std__pe5__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe5__lane26_strm1_cntl        = 'd0         ;
    std__pe5__lane26_strm1_data        = 'h1234_5678 ;
    std__pe5__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe5__lane27_strm0_cntl        = 'd0         ;
    std__pe5__lane27_strm0_data        = 'h1234_5678 ;
    std__pe5__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe5__lane27_strm1_cntl        = 'd0         ;
    std__pe5__lane27_strm1_data        = 'h1234_5678 ;
    std__pe5__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe5__lane28_strm0_cntl        = 'd0         ;
    std__pe5__lane28_strm0_data        = 'h1234_5678 ;
    std__pe5__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe5__lane28_strm1_cntl        = 'd0         ;
    std__pe5__lane28_strm1_data        = 'h1234_5678 ;
    std__pe5__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe5__lane29_strm0_cntl        = 'd0         ;
    std__pe5__lane29_strm0_data        = 'h1234_5678 ;
    std__pe5__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe5__lane29_strm1_cntl        = 'd0         ;
    std__pe5__lane29_strm1_data        = 'h1234_5678 ;
    std__pe5__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe5__lane30_strm0_cntl        = 'd0         ;
    std__pe5__lane30_strm0_data        = 'h1234_5678 ;
    std__pe5__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe5__lane30_strm1_cntl        = 'd0         ;
    std__pe5__lane30_strm1_data        = 'h1234_5678 ;
    std__pe5__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe5__lane31_strm0_cntl        = 'd0         ;
    std__pe5__lane31_strm0_data        = 'h1234_5678 ;
    std__pe5__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe5__lane31_strm1_cntl        = 'd0         ;
    std__pe5__lane31_strm1_data        = 'h1234_5678 ;
    std__pe5__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe6__lane0_strm0_cntl        = 'd0         ;
    std__pe6__lane0_strm0_data        = 'h1234_5678 ;
    std__pe6__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe6__lane0_strm1_cntl        = 'd0         ;
    std__pe6__lane0_strm1_data        = 'h1234_5678 ;
    std__pe6__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe6__lane1_strm0_cntl        = 'd0         ;
    std__pe6__lane1_strm0_data        = 'h1234_5678 ;
    std__pe6__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe6__lane1_strm1_cntl        = 'd0         ;
    std__pe6__lane1_strm1_data        = 'h1234_5678 ;
    std__pe6__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe6__lane2_strm0_cntl        = 'd0         ;
    std__pe6__lane2_strm0_data        = 'h1234_5678 ;
    std__pe6__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe6__lane2_strm1_cntl        = 'd0         ;
    std__pe6__lane2_strm1_data        = 'h1234_5678 ;
    std__pe6__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe6__lane3_strm0_cntl        = 'd0         ;
    std__pe6__lane3_strm0_data        = 'h1234_5678 ;
    std__pe6__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe6__lane3_strm1_cntl        = 'd0         ;
    std__pe6__lane3_strm1_data        = 'h1234_5678 ;
    std__pe6__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe6__lane4_strm0_cntl        = 'd0         ;
    std__pe6__lane4_strm0_data        = 'h1234_5678 ;
    std__pe6__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe6__lane4_strm1_cntl        = 'd0         ;
    std__pe6__lane4_strm1_data        = 'h1234_5678 ;
    std__pe6__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe6__lane5_strm0_cntl        = 'd0         ;
    std__pe6__lane5_strm0_data        = 'h1234_5678 ;
    std__pe6__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe6__lane5_strm1_cntl        = 'd0         ;
    std__pe6__lane5_strm1_data        = 'h1234_5678 ;
    std__pe6__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe6__lane6_strm0_cntl        = 'd0         ;
    std__pe6__lane6_strm0_data        = 'h1234_5678 ;
    std__pe6__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe6__lane6_strm1_cntl        = 'd0         ;
    std__pe6__lane6_strm1_data        = 'h1234_5678 ;
    std__pe6__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe6__lane7_strm0_cntl        = 'd0         ;
    std__pe6__lane7_strm0_data        = 'h1234_5678 ;
    std__pe6__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe6__lane7_strm1_cntl        = 'd0         ;
    std__pe6__lane7_strm1_data        = 'h1234_5678 ;
    std__pe6__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe6__lane8_strm0_cntl        = 'd0         ;
    std__pe6__lane8_strm0_data        = 'h1234_5678 ;
    std__pe6__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe6__lane8_strm1_cntl        = 'd0         ;
    std__pe6__lane8_strm1_data        = 'h1234_5678 ;
    std__pe6__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe6__lane9_strm0_cntl        = 'd0         ;
    std__pe6__lane9_strm0_data        = 'h1234_5678 ;
    std__pe6__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe6__lane9_strm1_cntl        = 'd0         ;
    std__pe6__lane9_strm1_data        = 'h1234_5678 ;
    std__pe6__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe6__lane10_strm0_cntl        = 'd0         ;
    std__pe6__lane10_strm0_data        = 'h1234_5678 ;
    std__pe6__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe6__lane10_strm1_cntl        = 'd0         ;
    std__pe6__lane10_strm1_data        = 'h1234_5678 ;
    std__pe6__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe6__lane11_strm0_cntl        = 'd0         ;
    std__pe6__lane11_strm0_data        = 'h1234_5678 ;
    std__pe6__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe6__lane11_strm1_cntl        = 'd0         ;
    std__pe6__lane11_strm1_data        = 'h1234_5678 ;
    std__pe6__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe6__lane12_strm0_cntl        = 'd0         ;
    std__pe6__lane12_strm0_data        = 'h1234_5678 ;
    std__pe6__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe6__lane12_strm1_cntl        = 'd0         ;
    std__pe6__lane12_strm1_data        = 'h1234_5678 ;
    std__pe6__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe6__lane13_strm0_cntl        = 'd0         ;
    std__pe6__lane13_strm0_data        = 'h1234_5678 ;
    std__pe6__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe6__lane13_strm1_cntl        = 'd0         ;
    std__pe6__lane13_strm1_data        = 'h1234_5678 ;
    std__pe6__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe6__lane14_strm0_cntl        = 'd0         ;
    std__pe6__lane14_strm0_data        = 'h1234_5678 ;
    std__pe6__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe6__lane14_strm1_cntl        = 'd0         ;
    std__pe6__lane14_strm1_data        = 'h1234_5678 ;
    std__pe6__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe6__lane15_strm0_cntl        = 'd0         ;
    std__pe6__lane15_strm0_data        = 'h1234_5678 ;
    std__pe6__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe6__lane15_strm1_cntl        = 'd0         ;
    std__pe6__lane15_strm1_data        = 'h1234_5678 ;
    std__pe6__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe6__lane16_strm0_cntl        = 'd0         ;
    std__pe6__lane16_strm0_data        = 'h1234_5678 ;
    std__pe6__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe6__lane16_strm1_cntl        = 'd0         ;
    std__pe6__lane16_strm1_data        = 'h1234_5678 ;
    std__pe6__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe6__lane17_strm0_cntl        = 'd0         ;
    std__pe6__lane17_strm0_data        = 'h1234_5678 ;
    std__pe6__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe6__lane17_strm1_cntl        = 'd0         ;
    std__pe6__lane17_strm1_data        = 'h1234_5678 ;
    std__pe6__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe6__lane18_strm0_cntl        = 'd0         ;
    std__pe6__lane18_strm0_data        = 'h1234_5678 ;
    std__pe6__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe6__lane18_strm1_cntl        = 'd0         ;
    std__pe6__lane18_strm1_data        = 'h1234_5678 ;
    std__pe6__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe6__lane19_strm0_cntl        = 'd0         ;
    std__pe6__lane19_strm0_data        = 'h1234_5678 ;
    std__pe6__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe6__lane19_strm1_cntl        = 'd0         ;
    std__pe6__lane19_strm1_data        = 'h1234_5678 ;
    std__pe6__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe6__lane20_strm0_cntl        = 'd0         ;
    std__pe6__lane20_strm0_data        = 'h1234_5678 ;
    std__pe6__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe6__lane20_strm1_cntl        = 'd0         ;
    std__pe6__lane20_strm1_data        = 'h1234_5678 ;
    std__pe6__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe6__lane21_strm0_cntl        = 'd0         ;
    std__pe6__lane21_strm0_data        = 'h1234_5678 ;
    std__pe6__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe6__lane21_strm1_cntl        = 'd0         ;
    std__pe6__lane21_strm1_data        = 'h1234_5678 ;
    std__pe6__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe6__lane22_strm0_cntl        = 'd0         ;
    std__pe6__lane22_strm0_data        = 'h1234_5678 ;
    std__pe6__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe6__lane22_strm1_cntl        = 'd0         ;
    std__pe6__lane22_strm1_data        = 'h1234_5678 ;
    std__pe6__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe6__lane23_strm0_cntl        = 'd0         ;
    std__pe6__lane23_strm0_data        = 'h1234_5678 ;
    std__pe6__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe6__lane23_strm1_cntl        = 'd0         ;
    std__pe6__lane23_strm1_data        = 'h1234_5678 ;
    std__pe6__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe6__lane24_strm0_cntl        = 'd0         ;
    std__pe6__lane24_strm0_data        = 'h1234_5678 ;
    std__pe6__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe6__lane24_strm1_cntl        = 'd0         ;
    std__pe6__lane24_strm1_data        = 'h1234_5678 ;
    std__pe6__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe6__lane25_strm0_cntl        = 'd0         ;
    std__pe6__lane25_strm0_data        = 'h1234_5678 ;
    std__pe6__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe6__lane25_strm1_cntl        = 'd0         ;
    std__pe6__lane25_strm1_data        = 'h1234_5678 ;
    std__pe6__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe6__lane26_strm0_cntl        = 'd0         ;
    std__pe6__lane26_strm0_data        = 'h1234_5678 ;
    std__pe6__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe6__lane26_strm1_cntl        = 'd0         ;
    std__pe6__lane26_strm1_data        = 'h1234_5678 ;
    std__pe6__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe6__lane27_strm0_cntl        = 'd0         ;
    std__pe6__lane27_strm0_data        = 'h1234_5678 ;
    std__pe6__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe6__lane27_strm1_cntl        = 'd0         ;
    std__pe6__lane27_strm1_data        = 'h1234_5678 ;
    std__pe6__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe6__lane28_strm0_cntl        = 'd0         ;
    std__pe6__lane28_strm0_data        = 'h1234_5678 ;
    std__pe6__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe6__lane28_strm1_cntl        = 'd0         ;
    std__pe6__lane28_strm1_data        = 'h1234_5678 ;
    std__pe6__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe6__lane29_strm0_cntl        = 'd0         ;
    std__pe6__lane29_strm0_data        = 'h1234_5678 ;
    std__pe6__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe6__lane29_strm1_cntl        = 'd0         ;
    std__pe6__lane29_strm1_data        = 'h1234_5678 ;
    std__pe6__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe6__lane30_strm0_cntl        = 'd0         ;
    std__pe6__lane30_strm0_data        = 'h1234_5678 ;
    std__pe6__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe6__lane30_strm1_cntl        = 'd0         ;
    std__pe6__lane30_strm1_data        = 'h1234_5678 ;
    std__pe6__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe6__lane31_strm0_cntl        = 'd0         ;
    std__pe6__lane31_strm0_data        = 'h1234_5678 ;
    std__pe6__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe6__lane31_strm1_cntl        = 'd0         ;
    std__pe6__lane31_strm1_data        = 'h1234_5678 ;
    std__pe6__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe7__lane0_strm0_cntl        = 'd0         ;
    std__pe7__lane0_strm0_data        = 'h1234_5678 ;
    std__pe7__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe7__lane0_strm1_cntl        = 'd0         ;
    std__pe7__lane0_strm1_data        = 'h1234_5678 ;
    std__pe7__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe7__lane1_strm0_cntl        = 'd0         ;
    std__pe7__lane1_strm0_data        = 'h1234_5678 ;
    std__pe7__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe7__lane1_strm1_cntl        = 'd0         ;
    std__pe7__lane1_strm1_data        = 'h1234_5678 ;
    std__pe7__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe7__lane2_strm0_cntl        = 'd0         ;
    std__pe7__lane2_strm0_data        = 'h1234_5678 ;
    std__pe7__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe7__lane2_strm1_cntl        = 'd0         ;
    std__pe7__lane2_strm1_data        = 'h1234_5678 ;
    std__pe7__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe7__lane3_strm0_cntl        = 'd0         ;
    std__pe7__lane3_strm0_data        = 'h1234_5678 ;
    std__pe7__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe7__lane3_strm1_cntl        = 'd0         ;
    std__pe7__lane3_strm1_data        = 'h1234_5678 ;
    std__pe7__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe7__lane4_strm0_cntl        = 'd0         ;
    std__pe7__lane4_strm0_data        = 'h1234_5678 ;
    std__pe7__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe7__lane4_strm1_cntl        = 'd0         ;
    std__pe7__lane4_strm1_data        = 'h1234_5678 ;
    std__pe7__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe7__lane5_strm0_cntl        = 'd0         ;
    std__pe7__lane5_strm0_data        = 'h1234_5678 ;
    std__pe7__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe7__lane5_strm1_cntl        = 'd0         ;
    std__pe7__lane5_strm1_data        = 'h1234_5678 ;
    std__pe7__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe7__lane6_strm0_cntl        = 'd0         ;
    std__pe7__lane6_strm0_data        = 'h1234_5678 ;
    std__pe7__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe7__lane6_strm1_cntl        = 'd0         ;
    std__pe7__lane6_strm1_data        = 'h1234_5678 ;
    std__pe7__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe7__lane7_strm0_cntl        = 'd0         ;
    std__pe7__lane7_strm0_data        = 'h1234_5678 ;
    std__pe7__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe7__lane7_strm1_cntl        = 'd0         ;
    std__pe7__lane7_strm1_data        = 'h1234_5678 ;
    std__pe7__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe7__lane8_strm0_cntl        = 'd0         ;
    std__pe7__lane8_strm0_data        = 'h1234_5678 ;
    std__pe7__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe7__lane8_strm1_cntl        = 'd0         ;
    std__pe7__lane8_strm1_data        = 'h1234_5678 ;
    std__pe7__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe7__lane9_strm0_cntl        = 'd0         ;
    std__pe7__lane9_strm0_data        = 'h1234_5678 ;
    std__pe7__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe7__lane9_strm1_cntl        = 'd0         ;
    std__pe7__lane9_strm1_data        = 'h1234_5678 ;
    std__pe7__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe7__lane10_strm0_cntl        = 'd0         ;
    std__pe7__lane10_strm0_data        = 'h1234_5678 ;
    std__pe7__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe7__lane10_strm1_cntl        = 'd0         ;
    std__pe7__lane10_strm1_data        = 'h1234_5678 ;
    std__pe7__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe7__lane11_strm0_cntl        = 'd0         ;
    std__pe7__lane11_strm0_data        = 'h1234_5678 ;
    std__pe7__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe7__lane11_strm1_cntl        = 'd0         ;
    std__pe7__lane11_strm1_data        = 'h1234_5678 ;
    std__pe7__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe7__lane12_strm0_cntl        = 'd0         ;
    std__pe7__lane12_strm0_data        = 'h1234_5678 ;
    std__pe7__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe7__lane12_strm1_cntl        = 'd0         ;
    std__pe7__lane12_strm1_data        = 'h1234_5678 ;
    std__pe7__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe7__lane13_strm0_cntl        = 'd0         ;
    std__pe7__lane13_strm0_data        = 'h1234_5678 ;
    std__pe7__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe7__lane13_strm1_cntl        = 'd0         ;
    std__pe7__lane13_strm1_data        = 'h1234_5678 ;
    std__pe7__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe7__lane14_strm0_cntl        = 'd0         ;
    std__pe7__lane14_strm0_data        = 'h1234_5678 ;
    std__pe7__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe7__lane14_strm1_cntl        = 'd0         ;
    std__pe7__lane14_strm1_data        = 'h1234_5678 ;
    std__pe7__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe7__lane15_strm0_cntl        = 'd0         ;
    std__pe7__lane15_strm0_data        = 'h1234_5678 ;
    std__pe7__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe7__lane15_strm1_cntl        = 'd0         ;
    std__pe7__lane15_strm1_data        = 'h1234_5678 ;
    std__pe7__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe7__lane16_strm0_cntl        = 'd0         ;
    std__pe7__lane16_strm0_data        = 'h1234_5678 ;
    std__pe7__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe7__lane16_strm1_cntl        = 'd0         ;
    std__pe7__lane16_strm1_data        = 'h1234_5678 ;
    std__pe7__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe7__lane17_strm0_cntl        = 'd0         ;
    std__pe7__lane17_strm0_data        = 'h1234_5678 ;
    std__pe7__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe7__lane17_strm1_cntl        = 'd0         ;
    std__pe7__lane17_strm1_data        = 'h1234_5678 ;
    std__pe7__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe7__lane18_strm0_cntl        = 'd0         ;
    std__pe7__lane18_strm0_data        = 'h1234_5678 ;
    std__pe7__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe7__lane18_strm1_cntl        = 'd0         ;
    std__pe7__lane18_strm1_data        = 'h1234_5678 ;
    std__pe7__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe7__lane19_strm0_cntl        = 'd0         ;
    std__pe7__lane19_strm0_data        = 'h1234_5678 ;
    std__pe7__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe7__lane19_strm1_cntl        = 'd0         ;
    std__pe7__lane19_strm1_data        = 'h1234_5678 ;
    std__pe7__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe7__lane20_strm0_cntl        = 'd0         ;
    std__pe7__lane20_strm0_data        = 'h1234_5678 ;
    std__pe7__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe7__lane20_strm1_cntl        = 'd0         ;
    std__pe7__lane20_strm1_data        = 'h1234_5678 ;
    std__pe7__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe7__lane21_strm0_cntl        = 'd0         ;
    std__pe7__lane21_strm0_data        = 'h1234_5678 ;
    std__pe7__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe7__lane21_strm1_cntl        = 'd0         ;
    std__pe7__lane21_strm1_data        = 'h1234_5678 ;
    std__pe7__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe7__lane22_strm0_cntl        = 'd0         ;
    std__pe7__lane22_strm0_data        = 'h1234_5678 ;
    std__pe7__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe7__lane22_strm1_cntl        = 'd0         ;
    std__pe7__lane22_strm1_data        = 'h1234_5678 ;
    std__pe7__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe7__lane23_strm0_cntl        = 'd0         ;
    std__pe7__lane23_strm0_data        = 'h1234_5678 ;
    std__pe7__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe7__lane23_strm1_cntl        = 'd0         ;
    std__pe7__lane23_strm1_data        = 'h1234_5678 ;
    std__pe7__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe7__lane24_strm0_cntl        = 'd0         ;
    std__pe7__lane24_strm0_data        = 'h1234_5678 ;
    std__pe7__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe7__lane24_strm1_cntl        = 'd0         ;
    std__pe7__lane24_strm1_data        = 'h1234_5678 ;
    std__pe7__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe7__lane25_strm0_cntl        = 'd0         ;
    std__pe7__lane25_strm0_data        = 'h1234_5678 ;
    std__pe7__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe7__lane25_strm1_cntl        = 'd0         ;
    std__pe7__lane25_strm1_data        = 'h1234_5678 ;
    std__pe7__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe7__lane26_strm0_cntl        = 'd0         ;
    std__pe7__lane26_strm0_data        = 'h1234_5678 ;
    std__pe7__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe7__lane26_strm1_cntl        = 'd0         ;
    std__pe7__lane26_strm1_data        = 'h1234_5678 ;
    std__pe7__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe7__lane27_strm0_cntl        = 'd0         ;
    std__pe7__lane27_strm0_data        = 'h1234_5678 ;
    std__pe7__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe7__lane27_strm1_cntl        = 'd0         ;
    std__pe7__lane27_strm1_data        = 'h1234_5678 ;
    std__pe7__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe7__lane28_strm0_cntl        = 'd0         ;
    std__pe7__lane28_strm0_data        = 'h1234_5678 ;
    std__pe7__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe7__lane28_strm1_cntl        = 'd0         ;
    std__pe7__lane28_strm1_data        = 'h1234_5678 ;
    std__pe7__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe7__lane29_strm0_cntl        = 'd0         ;
    std__pe7__lane29_strm0_data        = 'h1234_5678 ;
    std__pe7__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe7__lane29_strm1_cntl        = 'd0         ;
    std__pe7__lane29_strm1_data        = 'h1234_5678 ;
    std__pe7__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe7__lane30_strm0_cntl        = 'd0         ;
    std__pe7__lane30_strm0_data        = 'h1234_5678 ;
    std__pe7__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe7__lane30_strm1_cntl        = 'd0         ;
    std__pe7__lane30_strm1_data        = 'h1234_5678 ;
    std__pe7__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe7__lane31_strm0_cntl        = 'd0         ;
    std__pe7__lane31_strm0_data        = 'h1234_5678 ;
    std__pe7__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe7__lane31_strm1_cntl        = 'd0         ;
    std__pe7__lane31_strm1_data        = 'h1234_5678 ;
    std__pe7__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe8__lane0_strm0_cntl        = 'd0         ;
    std__pe8__lane0_strm0_data        = 'h1234_5678 ;
    std__pe8__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe8__lane0_strm1_cntl        = 'd0         ;
    std__pe8__lane0_strm1_data        = 'h1234_5678 ;
    std__pe8__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe8__lane1_strm0_cntl        = 'd0         ;
    std__pe8__lane1_strm0_data        = 'h1234_5678 ;
    std__pe8__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe8__lane1_strm1_cntl        = 'd0         ;
    std__pe8__lane1_strm1_data        = 'h1234_5678 ;
    std__pe8__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe8__lane2_strm0_cntl        = 'd0         ;
    std__pe8__lane2_strm0_data        = 'h1234_5678 ;
    std__pe8__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe8__lane2_strm1_cntl        = 'd0         ;
    std__pe8__lane2_strm1_data        = 'h1234_5678 ;
    std__pe8__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe8__lane3_strm0_cntl        = 'd0         ;
    std__pe8__lane3_strm0_data        = 'h1234_5678 ;
    std__pe8__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe8__lane3_strm1_cntl        = 'd0         ;
    std__pe8__lane3_strm1_data        = 'h1234_5678 ;
    std__pe8__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe8__lane4_strm0_cntl        = 'd0         ;
    std__pe8__lane4_strm0_data        = 'h1234_5678 ;
    std__pe8__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe8__lane4_strm1_cntl        = 'd0         ;
    std__pe8__lane4_strm1_data        = 'h1234_5678 ;
    std__pe8__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe8__lane5_strm0_cntl        = 'd0         ;
    std__pe8__lane5_strm0_data        = 'h1234_5678 ;
    std__pe8__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe8__lane5_strm1_cntl        = 'd0         ;
    std__pe8__lane5_strm1_data        = 'h1234_5678 ;
    std__pe8__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe8__lane6_strm0_cntl        = 'd0         ;
    std__pe8__lane6_strm0_data        = 'h1234_5678 ;
    std__pe8__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe8__lane6_strm1_cntl        = 'd0         ;
    std__pe8__lane6_strm1_data        = 'h1234_5678 ;
    std__pe8__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe8__lane7_strm0_cntl        = 'd0         ;
    std__pe8__lane7_strm0_data        = 'h1234_5678 ;
    std__pe8__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe8__lane7_strm1_cntl        = 'd0         ;
    std__pe8__lane7_strm1_data        = 'h1234_5678 ;
    std__pe8__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe8__lane8_strm0_cntl        = 'd0         ;
    std__pe8__lane8_strm0_data        = 'h1234_5678 ;
    std__pe8__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe8__lane8_strm1_cntl        = 'd0         ;
    std__pe8__lane8_strm1_data        = 'h1234_5678 ;
    std__pe8__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe8__lane9_strm0_cntl        = 'd0         ;
    std__pe8__lane9_strm0_data        = 'h1234_5678 ;
    std__pe8__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe8__lane9_strm1_cntl        = 'd0         ;
    std__pe8__lane9_strm1_data        = 'h1234_5678 ;
    std__pe8__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe8__lane10_strm0_cntl        = 'd0         ;
    std__pe8__lane10_strm0_data        = 'h1234_5678 ;
    std__pe8__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe8__lane10_strm1_cntl        = 'd0         ;
    std__pe8__lane10_strm1_data        = 'h1234_5678 ;
    std__pe8__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe8__lane11_strm0_cntl        = 'd0         ;
    std__pe8__lane11_strm0_data        = 'h1234_5678 ;
    std__pe8__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe8__lane11_strm1_cntl        = 'd0         ;
    std__pe8__lane11_strm1_data        = 'h1234_5678 ;
    std__pe8__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe8__lane12_strm0_cntl        = 'd0         ;
    std__pe8__lane12_strm0_data        = 'h1234_5678 ;
    std__pe8__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe8__lane12_strm1_cntl        = 'd0         ;
    std__pe8__lane12_strm1_data        = 'h1234_5678 ;
    std__pe8__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe8__lane13_strm0_cntl        = 'd0         ;
    std__pe8__lane13_strm0_data        = 'h1234_5678 ;
    std__pe8__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe8__lane13_strm1_cntl        = 'd0         ;
    std__pe8__lane13_strm1_data        = 'h1234_5678 ;
    std__pe8__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe8__lane14_strm0_cntl        = 'd0         ;
    std__pe8__lane14_strm0_data        = 'h1234_5678 ;
    std__pe8__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe8__lane14_strm1_cntl        = 'd0         ;
    std__pe8__lane14_strm1_data        = 'h1234_5678 ;
    std__pe8__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe8__lane15_strm0_cntl        = 'd0         ;
    std__pe8__lane15_strm0_data        = 'h1234_5678 ;
    std__pe8__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe8__lane15_strm1_cntl        = 'd0         ;
    std__pe8__lane15_strm1_data        = 'h1234_5678 ;
    std__pe8__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe8__lane16_strm0_cntl        = 'd0         ;
    std__pe8__lane16_strm0_data        = 'h1234_5678 ;
    std__pe8__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe8__lane16_strm1_cntl        = 'd0         ;
    std__pe8__lane16_strm1_data        = 'h1234_5678 ;
    std__pe8__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe8__lane17_strm0_cntl        = 'd0         ;
    std__pe8__lane17_strm0_data        = 'h1234_5678 ;
    std__pe8__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe8__lane17_strm1_cntl        = 'd0         ;
    std__pe8__lane17_strm1_data        = 'h1234_5678 ;
    std__pe8__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe8__lane18_strm0_cntl        = 'd0         ;
    std__pe8__lane18_strm0_data        = 'h1234_5678 ;
    std__pe8__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe8__lane18_strm1_cntl        = 'd0         ;
    std__pe8__lane18_strm1_data        = 'h1234_5678 ;
    std__pe8__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe8__lane19_strm0_cntl        = 'd0         ;
    std__pe8__lane19_strm0_data        = 'h1234_5678 ;
    std__pe8__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe8__lane19_strm1_cntl        = 'd0         ;
    std__pe8__lane19_strm1_data        = 'h1234_5678 ;
    std__pe8__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe8__lane20_strm0_cntl        = 'd0         ;
    std__pe8__lane20_strm0_data        = 'h1234_5678 ;
    std__pe8__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe8__lane20_strm1_cntl        = 'd0         ;
    std__pe8__lane20_strm1_data        = 'h1234_5678 ;
    std__pe8__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe8__lane21_strm0_cntl        = 'd0         ;
    std__pe8__lane21_strm0_data        = 'h1234_5678 ;
    std__pe8__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe8__lane21_strm1_cntl        = 'd0         ;
    std__pe8__lane21_strm1_data        = 'h1234_5678 ;
    std__pe8__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe8__lane22_strm0_cntl        = 'd0         ;
    std__pe8__lane22_strm0_data        = 'h1234_5678 ;
    std__pe8__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe8__lane22_strm1_cntl        = 'd0         ;
    std__pe8__lane22_strm1_data        = 'h1234_5678 ;
    std__pe8__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe8__lane23_strm0_cntl        = 'd0         ;
    std__pe8__lane23_strm0_data        = 'h1234_5678 ;
    std__pe8__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe8__lane23_strm1_cntl        = 'd0         ;
    std__pe8__lane23_strm1_data        = 'h1234_5678 ;
    std__pe8__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe8__lane24_strm0_cntl        = 'd0         ;
    std__pe8__lane24_strm0_data        = 'h1234_5678 ;
    std__pe8__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe8__lane24_strm1_cntl        = 'd0         ;
    std__pe8__lane24_strm1_data        = 'h1234_5678 ;
    std__pe8__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe8__lane25_strm0_cntl        = 'd0         ;
    std__pe8__lane25_strm0_data        = 'h1234_5678 ;
    std__pe8__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe8__lane25_strm1_cntl        = 'd0         ;
    std__pe8__lane25_strm1_data        = 'h1234_5678 ;
    std__pe8__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe8__lane26_strm0_cntl        = 'd0         ;
    std__pe8__lane26_strm0_data        = 'h1234_5678 ;
    std__pe8__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe8__lane26_strm1_cntl        = 'd0         ;
    std__pe8__lane26_strm1_data        = 'h1234_5678 ;
    std__pe8__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe8__lane27_strm0_cntl        = 'd0         ;
    std__pe8__lane27_strm0_data        = 'h1234_5678 ;
    std__pe8__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe8__lane27_strm1_cntl        = 'd0         ;
    std__pe8__lane27_strm1_data        = 'h1234_5678 ;
    std__pe8__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe8__lane28_strm0_cntl        = 'd0         ;
    std__pe8__lane28_strm0_data        = 'h1234_5678 ;
    std__pe8__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe8__lane28_strm1_cntl        = 'd0         ;
    std__pe8__lane28_strm1_data        = 'h1234_5678 ;
    std__pe8__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe8__lane29_strm0_cntl        = 'd0         ;
    std__pe8__lane29_strm0_data        = 'h1234_5678 ;
    std__pe8__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe8__lane29_strm1_cntl        = 'd0         ;
    std__pe8__lane29_strm1_data        = 'h1234_5678 ;
    std__pe8__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe8__lane30_strm0_cntl        = 'd0         ;
    std__pe8__lane30_strm0_data        = 'h1234_5678 ;
    std__pe8__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe8__lane30_strm1_cntl        = 'd0         ;
    std__pe8__lane30_strm1_data        = 'h1234_5678 ;
    std__pe8__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe8__lane31_strm0_cntl        = 'd0         ;
    std__pe8__lane31_strm0_data        = 'h1234_5678 ;
    std__pe8__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe8__lane31_strm1_cntl        = 'd0         ;
    std__pe8__lane31_strm1_data        = 'h1234_5678 ;
    std__pe8__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe9__lane0_strm0_cntl        = 'd0         ;
    std__pe9__lane0_strm0_data        = 'h1234_5678 ;
    std__pe9__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe9__lane0_strm1_cntl        = 'd0         ;
    std__pe9__lane0_strm1_data        = 'h1234_5678 ;
    std__pe9__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe9__lane1_strm0_cntl        = 'd0         ;
    std__pe9__lane1_strm0_data        = 'h1234_5678 ;
    std__pe9__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe9__lane1_strm1_cntl        = 'd0         ;
    std__pe9__lane1_strm1_data        = 'h1234_5678 ;
    std__pe9__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe9__lane2_strm0_cntl        = 'd0         ;
    std__pe9__lane2_strm0_data        = 'h1234_5678 ;
    std__pe9__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe9__lane2_strm1_cntl        = 'd0         ;
    std__pe9__lane2_strm1_data        = 'h1234_5678 ;
    std__pe9__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe9__lane3_strm0_cntl        = 'd0         ;
    std__pe9__lane3_strm0_data        = 'h1234_5678 ;
    std__pe9__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe9__lane3_strm1_cntl        = 'd0         ;
    std__pe9__lane3_strm1_data        = 'h1234_5678 ;
    std__pe9__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe9__lane4_strm0_cntl        = 'd0         ;
    std__pe9__lane4_strm0_data        = 'h1234_5678 ;
    std__pe9__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe9__lane4_strm1_cntl        = 'd0         ;
    std__pe9__lane4_strm1_data        = 'h1234_5678 ;
    std__pe9__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe9__lane5_strm0_cntl        = 'd0         ;
    std__pe9__lane5_strm0_data        = 'h1234_5678 ;
    std__pe9__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe9__lane5_strm1_cntl        = 'd0         ;
    std__pe9__lane5_strm1_data        = 'h1234_5678 ;
    std__pe9__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe9__lane6_strm0_cntl        = 'd0         ;
    std__pe9__lane6_strm0_data        = 'h1234_5678 ;
    std__pe9__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe9__lane6_strm1_cntl        = 'd0         ;
    std__pe9__lane6_strm1_data        = 'h1234_5678 ;
    std__pe9__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe9__lane7_strm0_cntl        = 'd0         ;
    std__pe9__lane7_strm0_data        = 'h1234_5678 ;
    std__pe9__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe9__lane7_strm1_cntl        = 'd0         ;
    std__pe9__lane7_strm1_data        = 'h1234_5678 ;
    std__pe9__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe9__lane8_strm0_cntl        = 'd0         ;
    std__pe9__lane8_strm0_data        = 'h1234_5678 ;
    std__pe9__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe9__lane8_strm1_cntl        = 'd0         ;
    std__pe9__lane8_strm1_data        = 'h1234_5678 ;
    std__pe9__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe9__lane9_strm0_cntl        = 'd0         ;
    std__pe9__lane9_strm0_data        = 'h1234_5678 ;
    std__pe9__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe9__lane9_strm1_cntl        = 'd0         ;
    std__pe9__lane9_strm1_data        = 'h1234_5678 ;
    std__pe9__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe9__lane10_strm0_cntl        = 'd0         ;
    std__pe9__lane10_strm0_data        = 'h1234_5678 ;
    std__pe9__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe9__lane10_strm1_cntl        = 'd0         ;
    std__pe9__lane10_strm1_data        = 'h1234_5678 ;
    std__pe9__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe9__lane11_strm0_cntl        = 'd0         ;
    std__pe9__lane11_strm0_data        = 'h1234_5678 ;
    std__pe9__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe9__lane11_strm1_cntl        = 'd0         ;
    std__pe9__lane11_strm1_data        = 'h1234_5678 ;
    std__pe9__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe9__lane12_strm0_cntl        = 'd0         ;
    std__pe9__lane12_strm0_data        = 'h1234_5678 ;
    std__pe9__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe9__lane12_strm1_cntl        = 'd0         ;
    std__pe9__lane12_strm1_data        = 'h1234_5678 ;
    std__pe9__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe9__lane13_strm0_cntl        = 'd0         ;
    std__pe9__lane13_strm0_data        = 'h1234_5678 ;
    std__pe9__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe9__lane13_strm1_cntl        = 'd0         ;
    std__pe9__lane13_strm1_data        = 'h1234_5678 ;
    std__pe9__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe9__lane14_strm0_cntl        = 'd0         ;
    std__pe9__lane14_strm0_data        = 'h1234_5678 ;
    std__pe9__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe9__lane14_strm1_cntl        = 'd0         ;
    std__pe9__lane14_strm1_data        = 'h1234_5678 ;
    std__pe9__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe9__lane15_strm0_cntl        = 'd0         ;
    std__pe9__lane15_strm0_data        = 'h1234_5678 ;
    std__pe9__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe9__lane15_strm1_cntl        = 'd0         ;
    std__pe9__lane15_strm1_data        = 'h1234_5678 ;
    std__pe9__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe9__lane16_strm0_cntl        = 'd0         ;
    std__pe9__lane16_strm0_data        = 'h1234_5678 ;
    std__pe9__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe9__lane16_strm1_cntl        = 'd0         ;
    std__pe9__lane16_strm1_data        = 'h1234_5678 ;
    std__pe9__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe9__lane17_strm0_cntl        = 'd0         ;
    std__pe9__lane17_strm0_data        = 'h1234_5678 ;
    std__pe9__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe9__lane17_strm1_cntl        = 'd0         ;
    std__pe9__lane17_strm1_data        = 'h1234_5678 ;
    std__pe9__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe9__lane18_strm0_cntl        = 'd0         ;
    std__pe9__lane18_strm0_data        = 'h1234_5678 ;
    std__pe9__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe9__lane18_strm1_cntl        = 'd0         ;
    std__pe9__lane18_strm1_data        = 'h1234_5678 ;
    std__pe9__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe9__lane19_strm0_cntl        = 'd0         ;
    std__pe9__lane19_strm0_data        = 'h1234_5678 ;
    std__pe9__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe9__lane19_strm1_cntl        = 'd0         ;
    std__pe9__lane19_strm1_data        = 'h1234_5678 ;
    std__pe9__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe9__lane20_strm0_cntl        = 'd0         ;
    std__pe9__lane20_strm0_data        = 'h1234_5678 ;
    std__pe9__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe9__lane20_strm1_cntl        = 'd0         ;
    std__pe9__lane20_strm1_data        = 'h1234_5678 ;
    std__pe9__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe9__lane21_strm0_cntl        = 'd0         ;
    std__pe9__lane21_strm0_data        = 'h1234_5678 ;
    std__pe9__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe9__lane21_strm1_cntl        = 'd0         ;
    std__pe9__lane21_strm1_data        = 'h1234_5678 ;
    std__pe9__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe9__lane22_strm0_cntl        = 'd0         ;
    std__pe9__lane22_strm0_data        = 'h1234_5678 ;
    std__pe9__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe9__lane22_strm1_cntl        = 'd0         ;
    std__pe9__lane22_strm1_data        = 'h1234_5678 ;
    std__pe9__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe9__lane23_strm0_cntl        = 'd0         ;
    std__pe9__lane23_strm0_data        = 'h1234_5678 ;
    std__pe9__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe9__lane23_strm1_cntl        = 'd0         ;
    std__pe9__lane23_strm1_data        = 'h1234_5678 ;
    std__pe9__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe9__lane24_strm0_cntl        = 'd0         ;
    std__pe9__lane24_strm0_data        = 'h1234_5678 ;
    std__pe9__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe9__lane24_strm1_cntl        = 'd0         ;
    std__pe9__lane24_strm1_data        = 'h1234_5678 ;
    std__pe9__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe9__lane25_strm0_cntl        = 'd0         ;
    std__pe9__lane25_strm0_data        = 'h1234_5678 ;
    std__pe9__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe9__lane25_strm1_cntl        = 'd0         ;
    std__pe9__lane25_strm1_data        = 'h1234_5678 ;
    std__pe9__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe9__lane26_strm0_cntl        = 'd0         ;
    std__pe9__lane26_strm0_data        = 'h1234_5678 ;
    std__pe9__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe9__lane26_strm1_cntl        = 'd0         ;
    std__pe9__lane26_strm1_data        = 'h1234_5678 ;
    std__pe9__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe9__lane27_strm0_cntl        = 'd0         ;
    std__pe9__lane27_strm0_data        = 'h1234_5678 ;
    std__pe9__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe9__lane27_strm1_cntl        = 'd0         ;
    std__pe9__lane27_strm1_data        = 'h1234_5678 ;
    std__pe9__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe9__lane28_strm0_cntl        = 'd0         ;
    std__pe9__lane28_strm0_data        = 'h1234_5678 ;
    std__pe9__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe9__lane28_strm1_cntl        = 'd0         ;
    std__pe9__lane28_strm1_data        = 'h1234_5678 ;
    std__pe9__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe9__lane29_strm0_cntl        = 'd0         ;
    std__pe9__lane29_strm0_data        = 'h1234_5678 ;
    std__pe9__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe9__lane29_strm1_cntl        = 'd0         ;
    std__pe9__lane29_strm1_data        = 'h1234_5678 ;
    std__pe9__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe9__lane30_strm0_cntl        = 'd0         ;
    std__pe9__lane30_strm0_data        = 'h1234_5678 ;
    std__pe9__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe9__lane30_strm1_cntl        = 'd0         ;
    std__pe9__lane30_strm1_data        = 'h1234_5678 ;
    std__pe9__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe9__lane31_strm0_cntl        = 'd0         ;
    std__pe9__lane31_strm0_data        = 'h1234_5678 ;
    std__pe9__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe9__lane31_strm1_cntl        = 'd0         ;
    std__pe9__lane31_strm1_data        = 'h1234_5678 ;
    std__pe9__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe10__lane0_strm0_cntl        = 'd0         ;
    std__pe10__lane0_strm0_data        = 'h1234_5678 ;
    std__pe10__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe10__lane0_strm1_cntl        = 'd0         ;
    std__pe10__lane0_strm1_data        = 'h1234_5678 ;
    std__pe10__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe10__lane1_strm0_cntl        = 'd0         ;
    std__pe10__lane1_strm0_data        = 'h1234_5678 ;
    std__pe10__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe10__lane1_strm1_cntl        = 'd0         ;
    std__pe10__lane1_strm1_data        = 'h1234_5678 ;
    std__pe10__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe10__lane2_strm0_cntl        = 'd0         ;
    std__pe10__lane2_strm0_data        = 'h1234_5678 ;
    std__pe10__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe10__lane2_strm1_cntl        = 'd0         ;
    std__pe10__lane2_strm1_data        = 'h1234_5678 ;
    std__pe10__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe10__lane3_strm0_cntl        = 'd0         ;
    std__pe10__lane3_strm0_data        = 'h1234_5678 ;
    std__pe10__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe10__lane3_strm1_cntl        = 'd0         ;
    std__pe10__lane3_strm1_data        = 'h1234_5678 ;
    std__pe10__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe10__lane4_strm0_cntl        = 'd0         ;
    std__pe10__lane4_strm0_data        = 'h1234_5678 ;
    std__pe10__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe10__lane4_strm1_cntl        = 'd0         ;
    std__pe10__lane4_strm1_data        = 'h1234_5678 ;
    std__pe10__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe10__lane5_strm0_cntl        = 'd0         ;
    std__pe10__lane5_strm0_data        = 'h1234_5678 ;
    std__pe10__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe10__lane5_strm1_cntl        = 'd0         ;
    std__pe10__lane5_strm1_data        = 'h1234_5678 ;
    std__pe10__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe10__lane6_strm0_cntl        = 'd0         ;
    std__pe10__lane6_strm0_data        = 'h1234_5678 ;
    std__pe10__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe10__lane6_strm1_cntl        = 'd0         ;
    std__pe10__lane6_strm1_data        = 'h1234_5678 ;
    std__pe10__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe10__lane7_strm0_cntl        = 'd0         ;
    std__pe10__lane7_strm0_data        = 'h1234_5678 ;
    std__pe10__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe10__lane7_strm1_cntl        = 'd0         ;
    std__pe10__lane7_strm1_data        = 'h1234_5678 ;
    std__pe10__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe10__lane8_strm0_cntl        = 'd0         ;
    std__pe10__lane8_strm0_data        = 'h1234_5678 ;
    std__pe10__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe10__lane8_strm1_cntl        = 'd0         ;
    std__pe10__lane8_strm1_data        = 'h1234_5678 ;
    std__pe10__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe10__lane9_strm0_cntl        = 'd0         ;
    std__pe10__lane9_strm0_data        = 'h1234_5678 ;
    std__pe10__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe10__lane9_strm1_cntl        = 'd0         ;
    std__pe10__lane9_strm1_data        = 'h1234_5678 ;
    std__pe10__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe10__lane10_strm0_cntl        = 'd0         ;
    std__pe10__lane10_strm0_data        = 'h1234_5678 ;
    std__pe10__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe10__lane10_strm1_cntl        = 'd0         ;
    std__pe10__lane10_strm1_data        = 'h1234_5678 ;
    std__pe10__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe10__lane11_strm0_cntl        = 'd0         ;
    std__pe10__lane11_strm0_data        = 'h1234_5678 ;
    std__pe10__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe10__lane11_strm1_cntl        = 'd0         ;
    std__pe10__lane11_strm1_data        = 'h1234_5678 ;
    std__pe10__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe10__lane12_strm0_cntl        = 'd0         ;
    std__pe10__lane12_strm0_data        = 'h1234_5678 ;
    std__pe10__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe10__lane12_strm1_cntl        = 'd0         ;
    std__pe10__lane12_strm1_data        = 'h1234_5678 ;
    std__pe10__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe10__lane13_strm0_cntl        = 'd0         ;
    std__pe10__lane13_strm0_data        = 'h1234_5678 ;
    std__pe10__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe10__lane13_strm1_cntl        = 'd0         ;
    std__pe10__lane13_strm1_data        = 'h1234_5678 ;
    std__pe10__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe10__lane14_strm0_cntl        = 'd0         ;
    std__pe10__lane14_strm0_data        = 'h1234_5678 ;
    std__pe10__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe10__lane14_strm1_cntl        = 'd0         ;
    std__pe10__lane14_strm1_data        = 'h1234_5678 ;
    std__pe10__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe10__lane15_strm0_cntl        = 'd0         ;
    std__pe10__lane15_strm0_data        = 'h1234_5678 ;
    std__pe10__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe10__lane15_strm1_cntl        = 'd0         ;
    std__pe10__lane15_strm1_data        = 'h1234_5678 ;
    std__pe10__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe10__lane16_strm0_cntl        = 'd0         ;
    std__pe10__lane16_strm0_data        = 'h1234_5678 ;
    std__pe10__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe10__lane16_strm1_cntl        = 'd0         ;
    std__pe10__lane16_strm1_data        = 'h1234_5678 ;
    std__pe10__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe10__lane17_strm0_cntl        = 'd0         ;
    std__pe10__lane17_strm0_data        = 'h1234_5678 ;
    std__pe10__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe10__lane17_strm1_cntl        = 'd0         ;
    std__pe10__lane17_strm1_data        = 'h1234_5678 ;
    std__pe10__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe10__lane18_strm0_cntl        = 'd0         ;
    std__pe10__lane18_strm0_data        = 'h1234_5678 ;
    std__pe10__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe10__lane18_strm1_cntl        = 'd0         ;
    std__pe10__lane18_strm1_data        = 'h1234_5678 ;
    std__pe10__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe10__lane19_strm0_cntl        = 'd0         ;
    std__pe10__lane19_strm0_data        = 'h1234_5678 ;
    std__pe10__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe10__lane19_strm1_cntl        = 'd0         ;
    std__pe10__lane19_strm1_data        = 'h1234_5678 ;
    std__pe10__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe10__lane20_strm0_cntl        = 'd0         ;
    std__pe10__lane20_strm0_data        = 'h1234_5678 ;
    std__pe10__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe10__lane20_strm1_cntl        = 'd0         ;
    std__pe10__lane20_strm1_data        = 'h1234_5678 ;
    std__pe10__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe10__lane21_strm0_cntl        = 'd0         ;
    std__pe10__lane21_strm0_data        = 'h1234_5678 ;
    std__pe10__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe10__lane21_strm1_cntl        = 'd0         ;
    std__pe10__lane21_strm1_data        = 'h1234_5678 ;
    std__pe10__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe10__lane22_strm0_cntl        = 'd0         ;
    std__pe10__lane22_strm0_data        = 'h1234_5678 ;
    std__pe10__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe10__lane22_strm1_cntl        = 'd0         ;
    std__pe10__lane22_strm1_data        = 'h1234_5678 ;
    std__pe10__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe10__lane23_strm0_cntl        = 'd0         ;
    std__pe10__lane23_strm0_data        = 'h1234_5678 ;
    std__pe10__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe10__lane23_strm1_cntl        = 'd0         ;
    std__pe10__lane23_strm1_data        = 'h1234_5678 ;
    std__pe10__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe10__lane24_strm0_cntl        = 'd0         ;
    std__pe10__lane24_strm0_data        = 'h1234_5678 ;
    std__pe10__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe10__lane24_strm1_cntl        = 'd0         ;
    std__pe10__lane24_strm1_data        = 'h1234_5678 ;
    std__pe10__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe10__lane25_strm0_cntl        = 'd0         ;
    std__pe10__lane25_strm0_data        = 'h1234_5678 ;
    std__pe10__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe10__lane25_strm1_cntl        = 'd0         ;
    std__pe10__lane25_strm1_data        = 'h1234_5678 ;
    std__pe10__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe10__lane26_strm0_cntl        = 'd0         ;
    std__pe10__lane26_strm0_data        = 'h1234_5678 ;
    std__pe10__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe10__lane26_strm1_cntl        = 'd0         ;
    std__pe10__lane26_strm1_data        = 'h1234_5678 ;
    std__pe10__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe10__lane27_strm0_cntl        = 'd0         ;
    std__pe10__lane27_strm0_data        = 'h1234_5678 ;
    std__pe10__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe10__lane27_strm1_cntl        = 'd0         ;
    std__pe10__lane27_strm1_data        = 'h1234_5678 ;
    std__pe10__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe10__lane28_strm0_cntl        = 'd0         ;
    std__pe10__lane28_strm0_data        = 'h1234_5678 ;
    std__pe10__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe10__lane28_strm1_cntl        = 'd0         ;
    std__pe10__lane28_strm1_data        = 'h1234_5678 ;
    std__pe10__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe10__lane29_strm0_cntl        = 'd0         ;
    std__pe10__lane29_strm0_data        = 'h1234_5678 ;
    std__pe10__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe10__lane29_strm1_cntl        = 'd0         ;
    std__pe10__lane29_strm1_data        = 'h1234_5678 ;
    std__pe10__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe10__lane30_strm0_cntl        = 'd0         ;
    std__pe10__lane30_strm0_data        = 'h1234_5678 ;
    std__pe10__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe10__lane30_strm1_cntl        = 'd0         ;
    std__pe10__lane30_strm1_data        = 'h1234_5678 ;
    std__pe10__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe10__lane31_strm0_cntl        = 'd0         ;
    std__pe10__lane31_strm0_data        = 'h1234_5678 ;
    std__pe10__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe10__lane31_strm1_cntl        = 'd0         ;
    std__pe10__lane31_strm1_data        = 'h1234_5678 ;
    std__pe10__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe11__lane0_strm0_cntl        = 'd0         ;
    std__pe11__lane0_strm0_data        = 'h1234_5678 ;
    std__pe11__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe11__lane0_strm1_cntl        = 'd0         ;
    std__pe11__lane0_strm1_data        = 'h1234_5678 ;
    std__pe11__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe11__lane1_strm0_cntl        = 'd0         ;
    std__pe11__lane1_strm0_data        = 'h1234_5678 ;
    std__pe11__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe11__lane1_strm1_cntl        = 'd0         ;
    std__pe11__lane1_strm1_data        = 'h1234_5678 ;
    std__pe11__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe11__lane2_strm0_cntl        = 'd0         ;
    std__pe11__lane2_strm0_data        = 'h1234_5678 ;
    std__pe11__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe11__lane2_strm1_cntl        = 'd0         ;
    std__pe11__lane2_strm1_data        = 'h1234_5678 ;
    std__pe11__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe11__lane3_strm0_cntl        = 'd0         ;
    std__pe11__lane3_strm0_data        = 'h1234_5678 ;
    std__pe11__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe11__lane3_strm1_cntl        = 'd0         ;
    std__pe11__lane3_strm1_data        = 'h1234_5678 ;
    std__pe11__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe11__lane4_strm0_cntl        = 'd0         ;
    std__pe11__lane4_strm0_data        = 'h1234_5678 ;
    std__pe11__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe11__lane4_strm1_cntl        = 'd0         ;
    std__pe11__lane4_strm1_data        = 'h1234_5678 ;
    std__pe11__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe11__lane5_strm0_cntl        = 'd0         ;
    std__pe11__lane5_strm0_data        = 'h1234_5678 ;
    std__pe11__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe11__lane5_strm1_cntl        = 'd0         ;
    std__pe11__lane5_strm1_data        = 'h1234_5678 ;
    std__pe11__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe11__lane6_strm0_cntl        = 'd0         ;
    std__pe11__lane6_strm0_data        = 'h1234_5678 ;
    std__pe11__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe11__lane6_strm1_cntl        = 'd0         ;
    std__pe11__lane6_strm1_data        = 'h1234_5678 ;
    std__pe11__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe11__lane7_strm0_cntl        = 'd0         ;
    std__pe11__lane7_strm0_data        = 'h1234_5678 ;
    std__pe11__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe11__lane7_strm1_cntl        = 'd0         ;
    std__pe11__lane7_strm1_data        = 'h1234_5678 ;
    std__pe11__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe11__lane8_strm0_cntl        = 'd0         ;
    std__pe11__lane8_strm0_data        = 'h1234_5678 ;
    std__pe11__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe11__lane8_strm1_cntl        = 'd0         ;
    std__pe11__lane8_strm1_data        = 'h1234_5678 ;
    std__pe11__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe11__lane9_strm0_cntl        = 'd0         ;
    std__pe11__lane9_strm0_data        = 'h1234_5678 ;
    std__pe11__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe11__lane9_strm1_cntl        = 'd0         ;
    std__pe11__lane9_strm1_data        = 'h1234_5678 ;
    std__pe11__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe11__lane10_strm0_cntl        = 'd0         ;
    std__pe11__lane10_strm0_data        = 'h1234_5678 ;
    std__pe11__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe11__lane10_strm1_cntl        = 'd0         ;
    std__pe11__lane10_strm1_data        = 'h1234_5678 ;
    std__pe11__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe11__lane11_strm0_cntl        = 'd0         ;
    std__pe11__lane11_strm0_data        = 'h1234_5678 ;
    std__pe11__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe11__lane11_strm1_cntl        = 'd0         ;
    std__pe11__lane11_strm1_data        = 'h1234_5678 ;
    std__pe11__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe11__lane12_strm0_cntl        = 'd0         ;
    std__pe11__lane12_strm0_data        = 'h1234_5678 ;
    std__pe11__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe11__lane12_strm1_cntl        = 'd0         ;
    std__pe11__lane12_strm1_data        = 'h1234_5678 ;
    std__pe11__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe11__lane13_strm0_cntl        = 'd0         ;
    std__pe11__lane13_strm0_data        = 'h1234_5678 ;
    std__pe11__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe11__lane13_strm1_cntl        = 'd0         ;
    std__pe11__lane13_strm1_data        = 'h1234_5678 ;
    std__pe11__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe11__lane14_strm0_cntl        = 'd0         ;
    std__pe11__lane14_strm0_data        = 'h1234_5678 ;
    std__pe11__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe11__lane14_strm1_cntl        = 'd0         ;
    std__pe11__lane14_strm1_data        = 'h1234_5678 ;
    std__pe11__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe11__lane15_strm0_cntl        = 'd0         ;
    std__pe11__lane15_strm0_data        = 'h1234_5678 ;
    std__pe11__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe11__lane15_strm1_cntl        = 'd0         ;
    std__pe11__lane15_strm1_data        = 'h1234_5678 ;
    std__pe11__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe11__lane16_strm0_cntl        = 'd0         ;
    std__pe11__lane16_strm0_data        = 'h1234_5678 ;
    std__pe11__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe11__lane16_strm1_cntl        = 'd0         ;
    std__pe11__lane16_strm1_data        = 'h1234_5678 ;
    std__pe11__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe11__lane17_strm0_cntl        = 'd0         ;
    std__pe11__lane17_strm0_data        = 'h1234_5678 ;
    std__pe11__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe11__lane17_strm1_cntl        = 'd0         ;
    std__pe11__lane17_strm1_data        = 'h1234_5678 ;
    std__pe11__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe11__lane18_strm0_cntl        = 'd0         ;
    std__pe11__lane18_strm0_data        = 'h1234_5678 ;
    std__pe11__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe11__lane18_strm1_cntl        = 'd0         ;
    std__pe11__lane18_strm1_data        = 'h1234_5678 ;
    std__pe11__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe11__lane19_strm0_cntl        = 'd0         ;
    std__pe11__lane19_strm0_data        = 'h1234_5678 ;
    std__pe11__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe11__lane19_strm1_cntl        = 'd0         ;
    std__pe11__lane19_strm1_data        = 'h1234_5678 ;
    std__pe11__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe11__lane20_strm0_cntl        = 'd0         ;
    std__pe11__lane20_strm0_data        = 'h1234_5678 ;
    std__pe11__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe11__lane20_strm1_cntl        = 'd0         ;
    std__pe11__lane20_strm1_data        = 'h1234_5678 ;
    std__pe11__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe11__lane21_strm0_cntl        = 'd0         ;
    std__pe11__lane21_strm0_data        = 'h1234_5678 ;
    std__pe11__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe11__lane21_strm1_cntl        = 'd0         ;
    std__pe11__lane21_strm1_data        = 'h1234_5678 ;
    std__pe11__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe11__lane22_strm0_cntl        = 'd0         ;
    std__pe11__lane22_strm0_data        = 'h1234_5678 ;
    std__pe11__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe11__lane22_strm1_cntl        = 'd0         ;
    std__pe11__lane22_strm1_data        = 'h1234_5678 ;
    std__pe11__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe11__lane23_strm0_cntl        = 'd0         ;
    std__pe11__lane23_strm0_data        = 'h1234_5678 ;
    std__pe11__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe11__lane23_strm1_cntl        = 'd0         ;
    std__pe11__lane23_strm1_data        = 'h1234_5678 ;
    std__pe11__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe11__lane24_strm0_cntl        = 'd0         ;
    std__pe11__lane24_strm0_data        = 'h1234_5678 ;
    std__pe11__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe11__lane24_strm1_cntl        = 'd0         ;
    std__pe11__lane24_strm1_data        = 'h1234_5678 ;
    std__pe11__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe11__lane25_strm0_cntl        = 'd0         ;
    std__pe11__lane25_strm0_data        = 'h1234_5678 ;
    std__pe11__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe11__lane25_strm1_cntl        = 'd0         ;
    std__pe11__lane25_strm1_data        = 'h1234_5678 ;
    std__pe11__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe11__lane26_strm0_cntl        = 'd0         ;
    std__pe11__lane26_strm0_data        = 'h1234_5678 ;
    std__pe11__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe11__lane26_strm1_cntl        = 'd0         ;
    std__pe11__lane26_strm1_data        = 'h1234_5678 ;
    std__pe11__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe11__lane27_strm0_cntl        = 'd0         ;
    std__pe11__lane27_strm0_data        = 'h1234_5678 ;
    std__pe11__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe11__lane27_strm1_cntl        = 'd0         ;
    std__pe11__lane27_strm1_data        = 'h1234_5678 ;
    std__pe11__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe11__lane28_strm0_cntl        = 'd0         ;
    std__pe11__lane28_strm0_data        = 'h1234_5678 ;
    std__pe11__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe11__lane28_strm1_cntl        = 'd0         ;
    std__pe11__lane28_strm1_data        = 'h1234_5678 ;
    std__pe11__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe11__lane29_strm0_cntl        = 'd0         ;
    std__pe11__lane29_strm0_data        = 'h1234_5678 ;
    std__pe11__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe11__lane29_strm1_cntl        = 'd0         ;
    std__pe11__lane29_strm1_data        = 'h1234_5678 ;
    std__pe11__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe11__lane30_strm0_cntl        = 'd0         ;
    std__pe11__lane30_strm0_data        = 'h1234_5678 ;
    std__pe11__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe11__lane30_strm1_cntl        = 'd0         ;
    std__pe11__lane30_strm1_data        = 'h1234_5678 ;
    std__pe11__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe11__lane31_strm0_cntl        = 'd0         ;
    std__pe11__lane31_strm0_data        = 'h1234_5678 ;
    std__pe11__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe11__lane31_strm1_cntl        = 'd0         ;
    std__pe11__lane31_strm1_data        = 'h1234_5678 ;
    std__pe11__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe12__lane0_strm0_cntl        = 'd0         ;
    std__pe12__lane0_strm0_data        = 'h1234_5678 ;
    std__pe12__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe12__lane0_strm1_cntl        = 'd0         ;
    std__pe12__lane0_strm1_data        = 'h1234_5678 ;
    std__pe12__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe12__lane1_strm0_cntl        = 'd0         ;
    std__pe12__lane1_strm0_data        = 'h1234_5678 ;
    std__pe12__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe12__lane1_strm1_cntl        = 'd0         ;
    std__pe12__lane1_strm1_data        = 'h1234_5678 ;
    std__pe12__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe12__lane2_strm0_cntl        = 'd0         ;
    std__pe12__lane2_strm0_data        = 'h1234_5678 ;
    std__pe12__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe12__lane2_strm1_cntl        = 'd0         ;
    std__pe12__lane2_strm1_data        = 'h1234_5678 ;
    std__pe12__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe12__lane3_strm0_cntl        = 'd0         ;
    std__pe12__lane3_strm0_data        = 'h1234_5678 ;
    std__pe12__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe12__lane3_strm1_cntl        = 'd0         ;
    std__pe12__lane3_strm1_data        = 'h1234_5678 ;
    std__pe12__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe12__lane4_strm0_cntl        = 'd0         ;
    std__pe12__lane4_strm0_data        = 'h1234_5678 ;
    std__pe12__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe12__lane4_strm1_cntl        = 'd0         ;
    std__pe12__lane4_strm1_data        = 'h1234_5678 ;
    std__pe12__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe12__lane5_strm0_cntl        = 'd0         ;
    std__pe12__lane5_strm0_data        = 'h1234_5678 ;
    std__pe12__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe12__lane5_strm1_cntl        = 'd0         ;
    std__pe12__lane5_strm1_data        = 'h1234_5678 ;
    std__pe12__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe12__lane6_strm0_cntl        = 'd0         ;
    std__pe12__lane6_strm0_data        = 'h1234_5678 ;
    std__pe12__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe12__lane6_strm1_cntl        = 'd0         ;
    std__pe12__lane6_strm1_data        = 'h1234_5678 ;
    std__pe12__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe12__lane7_strm0_cntl        = 'd0         ;
    std__pe12__lane7_strm0_data        = 'h1234_5678 ;
    std__pe12__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe12__lane7_strm1_cntl        = 'd0         ;
    std__pe12__lane7_strm1_data        = 'h1234_5678 ;
    std__pe12__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe12__lane8_strm0_cntl        = 'd0         ;
    std__pe12__lane8_strm0_data        = 'h1234_5678 ;
    std__pe12__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe12__lane8_strm1_cntl        = 'd0         ;
    std__pe12__lane8_strm1_data        = 'h1234_5678 ;
    std__pe12__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe12__lane9_strm0_cntl        = 'd0         ;
    std__pe12__lane9_strm0_data        = 'h1234_5678 ;
    std__pe12__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe12__lane9_strm1_cntl        = 'd0         ;
    std__pe12__lane9_strm1_data        = 'h1234_5678 ;
    std__pe12__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe12__lane10_strm0_cntl        = 'd0         ;
    std__pe12__lane10_strm0_data        = 'h1234_5678 ;
    std__pe12__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe12__lane10_strm1_cntl        = 'd0         ;
    std__pe12__lane10_strm1_data        = 'h1234_5678 ;
    std__pe12__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe12__lane11_strm0_cntl        = 'd0         ;
    std__pe12__lane11_strm0_data        = 'h1234_5678 ;
    std__pe12__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe12__lane11_strm1_cntl        = 'd0         ;
    std__pe12__lane11_strm1_data        = 'h1234_5678 ;
    std__pe12__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe12__lane12_strm0_cntl        = 'd0         ;
    std__pe12__lane12_strm0_data        = 'h1234_5678 ;
    std__pe12__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe12__lane12_strm1_cntl        = 'd0         ;
    std__pe12__lane12_strm1_data        = 'h1234_5678 ;
    std__pe12__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe12__lane13_strm0_cntl        = 'd0         ;
    std__pe12__lane13_strm0_data        = 'h1234_5678 ;
    std__pe12__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe12__lane13_strm1_cntl        = 'd0         ;
    std__pe12__lane13_strm1_data        = 'h1234_5678 ;
    std__pe12__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe12__lane14_strm0_cntl        = 'd0         ;
    std__pe12__lane14_strm0_data        = 'h1234_5678 ;
    std__pe12__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe12__lane14_strm1_cntl        = 'd0         ;
    std__pe12__lane14_strm1_data        = 'h1234_5678 ;
    std__pe12__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe12__lane15_strm0_cntl        = 'd0         ;
    std__pe12__lane15_strm0_data        = 'h1234_5678 ;
    std__pe12__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe12__lane15_strm1_cntl        = 'd0         ;
    std__pe12__lane15_strm1_data        = 'h1234_5678 ;
    std__pe12__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe12__lane16_strm0_cntl        = 'd0         ;
    std__pe12__lane16_strm0_data        = 'h1234_5678 ;
    std__pe12__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe12__lane16_strm1_cntl        = 'd0         ;
    std__pe12__lane16_strm1_data        = 'h1234_5678 ;
    std__pe12__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe12__lane17_strm0_cntl        = 'd0         ;
    std__pe12__lane17_strm0_data        = 'h1234_5678 ;
    std__pe12__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe12__lane17_strm1_cntl        = 'd0         ;
    std__pe12__lane17_strm1_data        = 'h1234_5678 ;
    std__pe12__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe12__lane18_strm0_cntl        = 'd0         ;
    std__pe12__lane18_strm0_data        = 'h1234_5678 ;
    std__pe12__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe12__lane18_strm1_cntl        = 'd0         ;
    std__pe12__lane18_strm1_data        = 'h1234_5678 ;
    std__pe12__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe12__lane19_strm0_cntl        = 'd0         ;
    std__pe12__lane19_strm0_data        = 'h1234_5678 ;
    std__pe12__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe12__lane19_strm1_cntl        = 'd0         ;
    std__pe12__lane19_strm1_data        = 'h1234_5678 ;
    std__pe12__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe12__lane20_strm0_cntl        = 'd0         ;
    std__pe12__lane20_strm0_data        = 'h1234_5678 ;
    std__pe12__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe12__lane20_strm1_cntl        = 'd0         ;
    std__pe12__lane20_strm1_data        = 'h1234_5678 ;
    std__pe12__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe12__lane21_strm0_cntl        = 'd0         ;
    std__pe12__lane21_strm0_data        = 'h1234_5678 ;
    std__pe12__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe12__lane21_strm1_cntl        = 'd0         ;
    std__pe12__lane21_strm1_data        = 'h1234_5678 ;
    std__pe12__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe12__lane22_strm0_cntl        = 'd0         ;
    std__pe12__lane22_strm0_data        = 'h1234_5678 ;
    std__pe12__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe12__lane22_strm1_cntl        = 'd0         ;
    std__pe12__lane22_strm1_data        = 'h1234_5678 ;
    std__pe12__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe12__lane23_strm0_cntl        = 'd0         ;
    std__pe12__lane23_strm0_data        = 'h1234_5678 ;
    std__pe12__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe12__lane23_strm1_cntl        = 'd0         ;
    std__pe12__lane23_strm1_data        = 'h1234_5678 ;
    std__pe12__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe12__lane24_strm0_cntl        = 'd0         ;
    std__pe12__lane24_strm0_data        = 'h1234_5678 ;
    std__pe12__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe12__lane24_strm1_cntl        = 'd0         ;
    std__pe12__lane24_strm1_data        = 'h1234_5678 ;
    std__pe12__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe12__lane25_strm0_cntl        = 'd0         ;
    std__pe12__lane25_strm0_data        = 'h1234_5678 ;
    std__pe12__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe12__lane25_strm1_cntl        = 'd0         ;
    std__pe12__lane25_strm1_data        = 'h1234_5678 ;
    std__pe12__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe12__lane26_strm0_cntl        = 'd0         ;
    std__pe12__lane26_strm0_data        = 'h1234_5678 ;
    std__pe12__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe12__lane26_strm1_cntl        = 'd0         ;
    std__pe12__lane26_strm1_data        = 'h1234_5678 ;
    std__pe12__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe12__lane27_strm0_cntl        = 'd0         ;
    std__pe12__lane27_strm0_data        = 'h1234_5678 ;
    std__pe12__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe12__lane27_strm1_cntl        = 'd0         ;
    std__pe12__lane27_strm1_data        = 'h1234_5678 ;
    std__pe12__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe12__lane28_strm0_cntl        = 'd0         ;
    std__pe12__lane28_strm0_data        = 'h1234_5678 ;
    std__pe12__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe12__lane28_strm1_cntl        = 'd0         ;
    std__pe12__lane28_strm1_data        = 'h1234_5678 ;
    std__pe12__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe12__lane29_strm0_cntl        = 'd0         ;
    std__pe12__lane29_strm0_data        = 'h1234_5678 ;
    std__pe12__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe12__lane29_strm1_cntl        = 'd0         ;
    std__pe12__lane29_strm1_data        = 'h1234_5678 ;
    std__pe12__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe12__lane30_strm0_cntl        = 'd0         ;
    std__pe12__lane30_strm0_data        = 'h1234_5678 ;
    std__pe12__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe12__lane30_strm1_cntl        = 'd0         ;
    std__pe12__lane30_strm1_data        = 'h1234_5678 ;
    std__pe12__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe12__lane31_strm0_cntl        = 'd0         ;
    std__pe12__lane31_strm0_data        = 'h1234_5678 ;
    std__pe12__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe12__lane31_strm1_cntl        = 'd0         ;
    std__pe12__lane31_strm1_data        = 'h1234_5678 ;
    std__pe12__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe13__lane0_strm0_cntl        = 'd0         ;
    std__pe13__lane0_strm0_data        = 'h1234_5678 ;
    std__pe13__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe13__lane0_strm1_cntl        = 'd0         ;
    std__pe13__lane0_strm1_data        = 'h1234_5678 ;
    std__pe13__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe13__lane1_strm0_cntl        = 'd0         ;
    std__pe13__lane1_strm0_data        = 'h1234_5678 ;
    std__pe13__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe13__lane1_strm1_cntl        = 'd0         ;
    std__pe13__lane1_strm1_data        = 'h1234_5678 ;
    std__pe13__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe13__lane2_strm0_cntl        = 'd0         ;
    std__pe13__lane2_strm0_data        = 'h1234_5678 ;
    std__pe13__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe13__lane2_strm1_cntl        = 'd0         ;
    std__pe13__lane2_strm1_data        = 'h1234_5678 ;
    std__pe13__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe13__lane3_strm0_cntl        = 'd0         ;
    std__pe13__lane3_strm0_data        = 'h1234_5678 ;
    std__pe13__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe13__lane3_strm1_cntl        = 'd0         ;
    std__pe13__lane3_strm1_data        = 'h1234_5678 ;
    std__pe13__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe13__lane4_strm0_cntl        = 'd0         ;
    std__pe13__lane4_strm0_data        = 'h1234_5678 ;
    std__pe13__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe13__lane4_strm1_cntl        = 'd0         ;
    std__pe13__lane4_strm1_data        = 'h1234_5678 ;
    std__pe13__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe13__lane5_strm0_cntl        = 'd0         ;
    std__pe13__lane5_strm0_data        = 'h1234_5678 ;
    std__pe13__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe13__lane5_strm1_cntl        = 'd0         ;
    std__pe13__lane5_strm1_data        = 'h1234_5678 ;
    std__pe13__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe13__lane6_strm0_cntl        = 'd0         ;
    std__pe13__lane6_strm0_data        = 'h1234_5678 ;
    std__pe13__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe13__lane6_strm1_cntl        = 'd0         ;
    std__pe13__lane6_strm1_data        = 'h1234_5678 ;
    std__pe13__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe13__lane7_strm0_cntl        = 'd0         ;
    std__pe13__lane7_strm0_data        = 'h1234_5678 ;
    std__pe13__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe13__lane7_strm1_cntl        = 'd0         ;
    std__pe13__lane7_strm1_data        = 'h1234_5678 ;
    std__pe13__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe13__lane8_strm0_cntl        = 'd0         ;
    std__pe13__lane8_strm0_data        = 'h1234_5678 ;
    std__pe13__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe13__lane8_strm1_cntl        = 'd0         ;
    std__pe13__lane8_strm1_data        = 'h1234_5678 ;
    std__pe13__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe13__lane9_strm0_cntl        = 'd0         ;
    std__pe13__lane9_strm0_data        = 'h1234_5678 ;
    std__pe13__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe13__lane9_strm1_cntl        = 'd0         ;
    std__pe13__lane9_strm1_data        = 'h1234_5678 ;
    std__pe13__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe13__lane10_strm0_cntl        = 'd0         ;
    std__pe13__lane10_strm0_data        = 'h1234_5678 ;
    std__pe13__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe13__lane10_strm1_cntl        = 'd0         ;
    std__pe13__lane10_strm1_data        = 'h1234_5678 ;
    std__pe13__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe13__lane11_strm0_cntl        = 'd0         ;
    std__pe13__lane11_strm0_data        = 'h1234_5678 ;
    std__pe13__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe13__lane11_strm1_cntl        = 'd0         ;
    std__pe13__lane11_strm1_data        = 'h1234_5678 ;
    std__pe13__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe13__lane12_strm0_cntl        = 'd0         ;
    std__pe13__lane12_strm0_data        = 'h1234_5678 ;
    std__pe13__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe13__lane12_strm1_cntl        = 'd0         ;
    std__pe13__lane12_strm1_data        = 'h1234_5678 ;
    std__pe13__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe13__lane13_strm0_cntl        = 'd0         ;
    std__pe13__lane13_strm0_data        = 'h1234_5678 ;
    std__pe13__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe13__lane13_strm1_cntl        = 'd0         ;
    std__pe13__lane13_strm1_data        = 'h1234_5678 ;
    std__pe13__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe13__lane14_strm0_cntl        = 'd0         ;
    std__pe13__lane14_strm0_data        = 'h1234_5678 ;
    std__pe13__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe13__lane14_strm1_cntl        = 'd0         ;
    std__pe13__lane14_strm1_data        = 'h1234_5678 ;
    std__pe13__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe13__lane15_strm0_cntl        = 'd0         ;
    std__pe13__lane15_strm0_data        = 'h1234_5678 ;
    std__pe13__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe13__lane15_strm1_cntl        = 'd0         ;
    std__pe13__lane15_strm1_data        = 'h1234_5678 ;
    std__pe13__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe13__lane16_strm0_cntl        = 'd0         ;
    std__pe13__lane16_strm0_data        = 'h1234_5678 ;
    std__pe13__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe13__lane16_strm1_cntl        = 'd0         ;
    std__pe13__lane16_strm1_data        = 'h1234_5678 ;
    std__pe13__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe13__lane17_strm0_cntl        = 'd0         ;
    std__pe13__lane17_strm0_data        = 'h1234_5678 ;
    std__pe13__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe13__lane17_strm1_cntl        = 'd0         ;
    std__pe13__lane17_strm1_data        = 'h1234_5678 ;
    std__pe13__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe13__lane18_strm0_cntl        = 'd0         ;
    std__pe13__lane18_strm0_data        = 'h1234_5678 ;
    std__pe13__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe13__lane18_strm1_cntl        = 'd0         ;
    std__pe13__lane18_strm1_data        = 'h1234_5678 ;
    std__pe13__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe13__lane19_strm0_cntl        = 'd0         ;
    std__pe13__lane19_strm0_data        = 'h1234_5678 ;
    std__pe13__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe13__lane19_strm1_cntl        = 'd0         ;
    std__pe13__lane19_strm1_data        = 'h1234_5678 ;
    std__pe13__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe13__lane20_strm0_cntl        = 'd0         ;
    std__pe13__lane20_strm0_data        = 'h1234_5678 ;
    std__pe13__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe13__lane20_strm1_cntl        = 'd0         ;
    std__pe13__lane20_strm1_data        = 'h1234_5678 ;
    std__pe13__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe13__lane21_strm0_cntl        = 'd0         ;
    std__pe13__lane21_strm0_data        = 'h1234_5678 ;
    std__pe13__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe13__lane21_strm1_cntl        = 'd0         ;
    std__pe13__lane21_strm1_data        = 'h1234_5678 ;
    std__pe13__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe13__lane22_strm0_cntl        = 'd0         ;
    std__pe13__lane22_strm0_data        = 'h1234_5678 ;
    std__pe13__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe13__lane22_strm1_cntl        = 'd0         ;
    std__pe13__lane22_strm1_data        = 'h1234_5678 ;
    std__pe13__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe13__lane23_strm0_cntl        = 'd0         ;
    std__pe13__lane23_strm0_data        = 'h1234_5678 ;
    std__pe13__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe13__lane23_strm1_cntl        = 'd0         ;
    std__pe13__lane23_strm1_data        = 'h1234_5678 ;
    std__pe13__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe13__lane24_strm0_cntl        = 'd0         ;
    std__pe13__lane24_strm0_data        = 'h1234_5678 ;
    std__pe13__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe13__lane24_strm1_cntl        = 'd0         ;
    std__pe13__lane24_strm1_data        = 'h1234_5678 ;
    std__pe13__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe13__lane25_strm0_cntl        = 'd0         ;
    std__pe13__lane25_strm0_data        = 'h1234_5678 ;
    std__pe13__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe13__lane25_strm1_cntl        = 'd0         ;
    std__pe13__lane25_strm1_data        = 'h1234_5678 ;
    std__pe13__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe13__lane26_strm0_cntl        = 'd0         ;
    std__pe13__lane26_strm0_data        = 'h1234_5678 ;
    std__pe13__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe13__lane26_strm1_cntl        = 'd0         ;
    std__pe13__lane26_strm1_data        = 'h1234_5678 ;
    std__pe13__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe13__lane27_strm0_cntl        = 'd0         ;
    std__pe13__lane27_strm0_data        = 'h1234_5678 ;
    std__pe13__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe13__lane27_strm1_cntl        = 'd0         ;
    std__pe13__lane27_strm1_data        = 'h1234_5678 ;
    std__pe13__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe13__lane28_strm0_cntl        = 'd0         ;
    std__pe13__lane28_strm0_data        = 'h1234_5678 ;
    std__pe13__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe13__lane28_strm1_cntl        = 'd0         ;
    std__pe13__lane28_strm1_data        = 'h1234_5678 ;
    std__pe13__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe13__lane29_strm0_cntl        = 'd0         ;
    std__pe13__lane29_strm0_data        = 'h1234_5678 ;
    std__pe13__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe13__lane29_strm1_cntl        = 'd0         ;
    std__pe13__lane29_strm1_data        = 'h1234_5678 ;
    std__pe13__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe13__lane30_strm0_cntl        = 'd0         ;
    std__pe13__lane30_strm0_data        = 'h1234_5678 ;
    std__pe13__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe13__lane30_strm1_cntl        = 'd0         ;
    std__pe13__lane30_strm1_data        = 'h1234_5678 ;
    std__pe13__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe13__lane31_strm0_cntl        = 'd0         ;
    std__pe13__lane31_strm0_data        = 'h1234_5678 ;
    std__pe13__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe13__lane31_strm1_cntl        = 'd0         ;
    std__pe13__lane31_strm1_data        = 'h1234_5678 ;
    std__pe13__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe14__lane0_strm0_cntl        = 'd0         ;
    std__pe14__lane0_strm0_data        = 'h1234_5678 ;
    std__pe14__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe14__lane0_strm1_cntl        = 'd0         ;
    std__pe14__lane0_strm1_data        = 'h1234_5678 ;
    std__pe14__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe14__lane1_strm0_cntl        = 'd0         ;
    std__pe14__lane1_strm0_data        = 'h1234_5678 ;
    std__pe14__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe14__lane1_strm1_cntl        = 'd0         ;
    std__pe14__lane1_strm1_data        = 'h1234_5678 ;
    std__pe14__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe14__lane2_strm0_cntl        = 'd0         ;
    std__pe14__lane2_strm0_data        = 'h1234_5678 ;
    std__pe14__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe14__lane2_strm1_cntl        = 'd0         ;
    std__pe14__lane2_strm1_data        = 'h1234_5678 ;
    std__pe14__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe14__lane3_strm0_cntl        = 'd0         ;
    std__pe14__lane3_strm0_data        = 'h1234_5678 ;
    std__pe14__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe14__lane3_strm1_cntl        = 'd0         ;
    std__pe14__lane3_strm1_data        = 'h1234_5678 ;
    std__pe14__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe14__lane4_strm0_cntl        = 'd0         ;
    std__pe14__lane4_strm0_data        = 'h1234_5678 ;
    std__pe14__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe14__lane4_strm1_cntl        = 'd0         ;
    std__pe14__lane4_strm1_data        = 'h1234_5678 ;
    std__pe14__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe14__lane5_strm0_cntl        = 'd0         ;
    std__pe14__lane5_strm0_data        = 'h1234_5678 ;
    std__pe14__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe14__lane5_strm1_cntl        = 'd0         ;
    std__pe14__lane5_strm1_data        = 'h1234_5678 ;
    std__pe14__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe14__lane6_strm0_cntl        = 'd0         ;
    std__pe14__lane6_strm0_data        = 'h1234_5678 ;
    std__pe14__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe14__lane6_strm1_cntl        = 'd0         ;
    std__pe14__lane6_strm1_data        = 'h1234_5678 ;
    std__pe14__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe14__lane7_strm0_cntl        = 'd0         ;
    std__pe14__lane7_strm0_data        = 'h1234_5678 ;
    std__pe14__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe14__lane7_strm1_cntl        = 'd0         ;
    std__pe14__lane7_strm1_data        = 'h1234_5678 ;
    std__pe14__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe14__lane8_strm0_cntl        = 'd0         ;
    std__pe14__lane8_strm0_data        = 'h1234_5678 ;
    std__pe14__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe14__lane8_strm1_cntl        = 'd0         ;
    std__pe14__lane8_strm1_data        = 'h1234_5678 ;
    std__pe14__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe14__lane9_strm0_cntl        = 'd0         ;
    std__pe14__lane9_strm0_data        = 'h1234_5678 ;
    std__pe14__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe14__lane9_strm1_cntl        = 'd0         ;
    std__pe14__lane9_strm1_data        = 'h1234_5678 ;
    std__pe14__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe14__lane10_strm0_cntl        = 'd0         ;
    std__pe14__lane10_strm0_data        = 'h1234_5678 ;
    std__pe14__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe14__lane10_strm1_cntl        = 'd0         ;
    std__pe14__lane10_strm1_data        = 'h1234_5678 ;
    std__pe14__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe14__lane11_strm0_cntl        = 'd0         ;
    std__pe14__lane11_strm0_data        = 'h1234_5678 ;
    std__pe14__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe14__lane11_strm1_cntl        = 'd0         ;
    std__pe14__lane11_strm1_data        = 'h1234_5678 ;
    std__pe14__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe14__lane12_strm0_cntl        = 'd0         ;
    std__pe14__lane12_strm0_data        = 'h1234_5678 ;
    std__pe14__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe14__lane12_strm1_cntl        = 'd0         ;
    std__pe14__lane12_strm1_data        = 'h1234_5678 ;
    std__pe14__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe14__lane13_strm0_cntl        = 'd0         ;
    std__pe14__lane13_strm0_data        = 'h1234_5678 ;
    std__pe14__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe14__lane13_strm1_cntl        = 'd0         ;
    std__pe14__lane13_strm1_data        = 'h1234_5678 ;
    std__pe14__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe14__lane14_strm0_cntl        = 'd0         ;
    std__pe14__lane14_strm0_data        = 'h1234_5678 ;
    std__pe14__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe14__lane14_strm1_cntl        = 'd0         ;
    std__pe14__lane14_strm1_data        = 'h1234_5678 ;
    std__pe14__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe14__lane15_strm0_cntl        = 'd0         ;
    std__pe14__lane15_strm0_data        = 'h1234_5678 ;
    std__pe14__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe14__lane15_strm1_cntl        = 'd0         ;
    std__pe14__lane15_strm1_data        = 'h1234_5678 ;
    std__pe14__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe14__lane16_strm0_cntl        = 'd0         ;
    std__pe14__lane16_strm0_data        = 'h1234_5678 ;
    std__pe14__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe14__lane16_strm1_cntl        = 'd0         ;
    std__pe14__lane16_strm1_data        = 'h1234_5678 ;
    std__pe14__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe14__lane17_strm0_cntl        = 'd0         ;
    std__pe14__lane17_strm0_data        = 'h1234_5678 ;
    std__pe14__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe14__lane17_strm1_cntl        = 'd0         ;
    std__pe14__lane17_strm1_data        = 'h1234_5678 ;
    std__pe14__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe14__lane18_strm0_cntl        = 'd0         ;
    std__pe14__lane18_strm0_data        = 'h1234_5678 ;
    std__pe14__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe14__lane18_strm1_cntl        = 'd0         ;
    std__pe14__lane18_strm1_data        = 'h1234_5678 ;
    std__pe14__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe14__lane19_strm0_cntl        = 'd0         ;
    std__pe14__lane19_strm0_data        = 'h1234_5678 ;
    std__pe14__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe14__lane19_strm1_cntl        = 'd0         ;
    std__pe14__lane19_strm1_data        = 'h1234_5678 ;
    std__pe14__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe14__lane20_strm0_cntl        = 'd0         ;
    std__pe14__lane20_strm0_data        = 'h1234_5678 ;
    std__pe14__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe14__lane20_strm1_cntl        = 'd0         ;
    std__pe14__lane20_strm1_data        = 'h1234_5678 ;
    std__pe14__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe14__lane21_strm0_cntl        = 'd0         ;
    std__pe14__lane21_strm0_data        = 'h1234_5678 ;
    std__pe14__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe14__lane21_strm1_cntl        = 'd0         ;
    std__pe14__lane21_strm1_data        = 'h1234_5678 ;
    std__pe14__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe14__lane22_strm0_cntl        = 'd0         ;
    std__pe14__lane22_strm0_data        = 'h1234_5678 ;
    std__pe14__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe14__lane22_strm1_cntl        = 'd0         ;
    std__pe14__lane22_strm1_data        = 'h1234_5678 ;
    std__pe14__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe14__lane23_strm0_cntl        = 'd0         ;
    std__pe14__lane23_strm0_data        = 'h1234_5678 ;
    std__pe14__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe14__lane23_strm1_cntl        = 'd0         ;
    std__pe14__lane23_strm1_data        = 'h1234_5678 ;
    std__pe14__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe14__lane24_strm0_cntl        = 'd0         ;
    std__pe14__lane24_strm0_data        = 'h1234_5678 ;
    std__pe14__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe14__lane24_strm1_cntl        = 'd0         ;
    std__pe14__lane24_strm1_data        = 'h1234_5678 ;
    std__pe14__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe14__lane25_strm0_cntl        = 'd0         ;
    std__pe14__lane25_strm0_data        = 'h1234_5678 ;
    std__pe14__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe14__lane25_strm1_cntl        = 'd0         ;
    std__pe14__lane25_strm1_data        = 'h1234_5678 ;
    std__pe14__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe14__lane26_strm0_cntl        = 'd0         ;
    std__pe14__lane26_strm0_data        = 'h1234_5678 ;
    std__pe14__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe14__lane26_strm1_cntl        = 'd0         ;
    std__pe14__lane26_strm1_data        = 'h1234_5678 ;
    std__pe14__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe14__lane27_strm0_cntl        = 'd0         ;
    std__pe14__lane27_strm0_data        = 'h1234_5678 ;
    std__pe14__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe14__lane27_strm1_cntl        = 'd0         ;
    std__pe14__lane27_strm1_data        = 'h1234_5678 ;
    std__pe14__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe14__lane28_strm0_cntl        = 'd0         ;
    std__pe14__lane28_strm0_data        = 'h1234_5678 ;
    std__pe14__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe14__lane28_strm1_cntl        = 'd0         ;
    std__pe14__lane28_strm1_data        = 'h1234_5678 ;
    std__pe14__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe14__lane29_strm0_cntl        = 'd0         ;
    std__pe14__lane29_strm0_data        = 'h1234_5678 ;
    std__pe14__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe14__lane29_strm1_cntl        = 'd0         ;
    std__pe14__lane29_strm1_data        = 'h1234_5678 ;
    std__pe14__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe14__lane30_strm0_cntl        = 'd0         ;
    std__pe14__lane30_strm0_data        = 'h1234_5678 ;
    std__pe14__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe14__lane30_strm1_cntl        = 'd0         ;
    std__pe14__lane30_strm1_data        = 'h1234_5678 ;
    std__pe14__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe14__lane31_strm0_cntl        = 'd0         ;
    std__pe14__lane31_strm0_data        = 'h1234_5678 ;
    std__pe14__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe14__lane31_strm1_cntl        = 'd0         ;
    std__pe14__lane31_strm1_data        = 'h1234_5678 ;
    std__pe14__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe15__lane0_strm0_cntl        = 'd0         ;
    std__pe15__lane0_strm0_data        = 'h1234_5678 ;
    std__pe15__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe15__lane0_strm1_cntl        = 'd0         ;
    std__pe15__lane0_strm1_data        = 'h1234_5678 ;
    std__pe15__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe15__lane1_strm0_cntl        = 'd0         ;
    std__pe15__lane1_strm0_data        = 'h1234_5678 ;
    std__pe15__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe15__lane1_strm1_cntl        = 'd0         ;
    std__pe15__lane1_strm1_data        = 'h1234_5678 ;
    std__pe15__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe15__lane2_strm0_cntl        = 'd0         ;
    std__pe15__lane2_strm0_data        = 'h1234_5678 ;
    std__pe15__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe15__lane2_strm1_cntl        = 'd0         ;
    std__pe15__lane2_strm1_data        = 'h1234_5678 ;
    std__pe15__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe15__lane3_strm0_cntl        = 'd0         ;
    std__pe15__lane3_strm0_data        = 'h1234_5678 ;
    std__pe15__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe15__lane3_strm1_cntl        = 'd0         ;
    std__pe15__lane3_strm1_data        = 'h1234_5678 ;
    std__pe15__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe15__lane4_strm0_cntl        = 'd0         ;
    std__pe15__lane4_strm0_data        = 'h1234_5678 ;
    std__pe15__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe15__lane4_strm1_cntl        = 'd0         ;
    std__pe15__lane4_strm1_data        = 'h1234_5678 ;
    std__pe15__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe15__lane5_strm0_cntl        = 'd0         ;
    std__pe15__lane5_strm0_data        = 'h1234_5678 ;
    std__pe15__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe15__lane5_strm1_cntl        = 'd0         ;
    std__pe15__lane5_strm1_data        = 'h1234_5678 ;
    std__pe15__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe15__lane6_strm0_cntl        = 'd0         ;
    std__pe15__lane6_strm0_data        = 'h1234_5678 ;
    std__pe15__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe15__lane6_strm1_cntl        = 'd0         ;
    std__pe15__lane6_strm1_data        = 'h1234_5678 ;
    std__pe15__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe15__lane7_strm0_cntl        = 'd0         ;
    std__pe15__lane7_strm0_data        = 'h1234_5678 ;
    std__pe15__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe15__lane7_strm1_cntl        = 'd0         ;
    std__pe15__lane7_strm1_data        = 'h1234_5678 ;
    std__pe15__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe15__lane8_strm0_cntl        = 'd0         ;
    std__pe15__lane8_strm0_data        = 'h1234_5678 ;
    std__pe15__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe15__lane8_strm1_cntl        = 'd0         ;
    std__pe15__lane8_strm1_data        = 'h1234_5678 ;
    std__pe15__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe15__lane9_strm0_cntl        = 'd0         ;
    std__pe15__lane9_strm0_data        = 'h1234_5678 ;
    std__pe15__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe15__lane9_strm1_cntl        = 'd0         ;
    std__pe15__lane9_strm1_data        = 'h1234_5678 ;
    std__pe15__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe15__lane10_strm0_cntl        = 'd0         ;
    std__pe15__lane10_strm0_data        = 'h1234_5678 ;
    std__pe15__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe15__lane10_strm1_cntl        = 'd0         ;
    std__pe15__lane10_strm1_data        = 'h1234_5678 ;
    std__pe15__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe15__lane11_strm0_cntl        = 'd0         ;
    std__pe15__lane11_strm0_data        = 'h1234_5678 ;
    std__pe15__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe15__lane11_strm1_cntl        = 'd0         ;
    std__pe15__lane11_strm1_data        = 'h1234_5678 ;
    std__pe15__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe15__lane12_strm0_cntl        = 'd0         ;
    std__pe15__lane12_strm0_data        = 'h1234_5678 ;
    std__pe15__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe15__lane12_strm1_cntl        = 'd0         ;
    std__pe15__lane12_strm1_data        = 'h1234_5678 ;
    std__pe15__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe15__lane13_strm0_cntl        = 'd0         ;
    std__pe15__lane13_strm0_data        = 'h1234_5678 ;
    std__pe15__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe15__lane13_strm1_cntl        = 'd0         ;
    std__pe15__lane13_strm1_data        = 'h1234_5678 ;
    std__pe15__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe15__lane14_strm0_cntl        = 'd0         ;
    std__pe15__lane14_strm0_data        = 'h1234_5678 ;
    std__pe15__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe15__lane14_strm1_cntl        = 'd0         ;
    std__pe15__lane14_strm1_data        = 'h1234_5678 ;
    std__pe15__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe15__lane15_strm0_cntl        = 'd0         ;
    std__pe15__lane15_strm0_data        = 'h1234_5678 ;
    std__pe15__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe15__lane15_strm1_cntl        = 'd0         ;
    std__pe15__lane15_strm1_data        = 'h1234_5678 ;
    std__pe15__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe15__lane16_strm0_cntl        = 'd0         ;
    std__pe15__lane16_strm0_data        = 'h1234_5678 ;
    std__pe15__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe15__lane16_strm1_cntl        = 'd0         ;
    std__pe15__lane16_strm1_data        = 'h1234_5678 ;
    std__pe15__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe15__lane17_strm0_cntl        = 'd0         ;
    std__pe15__lane17_strm0_data        = 'h1234_5678 ;
    std__pe15__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe15__lane17_strm1_cntl        = 'd0         ;
    std__pe15__lane17_strm1_data        = 'h1234_5678 ;
    std__pe15__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe15__lane18_strm0_cntl        = 'd0         ;
    std__pe15__lane18_strm0_data        = 'h1234_5678 ;
    std__pe15__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe15__lane18_strm1_cntl        = 'd0         ;
    std__pe15__lane18_strm1_data        = 'h1234_5678 ;
    std__pe15__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe15__lane19_strm0_cntl        = 'd0         ;
    std__pe15__lane19_strm0_data        = 'h1234_5678 ;
    std__pe15__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe15__lane19_strm1_cntl        = 'd0         ;
    std__pe15__lane19_strm1_data        = 'h1234_5678 ;
    std__pe15__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe15__lane20_strm0_cntl        = 'd0         ;
    std__pe15__lane20_strm0_data        = 'h1234_5678 ;
    std__pe15__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe15__lane20_strm1_cntl        = 'd0         ;
    std__pe15__lane20_strm1_data        = 'h1234_5678 ;
    std__pe15__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe15__lane21_strm0_cntl        = 'd0         ;
    std__pe15__lane21_strm0_data        = 'h1234_5678 ;
    std__pe15__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe15__lane21_strm1_cntl        = 'd0         ;
    std__pe15__lane21_strm1_data        = 'h1234_5678 ;
    std__pe15__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe15__lane22_strm0_cntl        = 'd0         ;
    std__pe15__lane22_strm0_data        = 'h1234_5678 ;
    std__pe15__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe15__lane22_strm1_cntl        = 'd0         ;
    std__pe15__lane22_strm1_data        = 'h1234_5678 ;
    std__pe15__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe15__lane23_strm0_cntl        = 'd0         ;
    std__pe15__lane23_strm0_data        = 'h1234_5678 ;
    std__pe15__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe15__lane23_strm1_cntl        = 'd0         ;
    std__pe15__lane23_strm1_data        = 'h1234_5678 ;
    std__pe15__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe15__lane24_strm0_cntl        = 'd0         ;
    std__pe15__lane24_strm0_data        = 'h1234_5678 ;
    std__pe15__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe15__lane24_strm1_cntl        = 'd0         ;
    std__pe15__lane24_strm1_data        = 'h1234_5678 ;
    std__pe15__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe15__lane25_strm0_cntl        = 'd0         ;
    std__pe15__lane25_strm0_data        = 'h1234_5678 ;
    std__pe15__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe15__lane25_strm1_cntl        = 'd0         ;
    std__pe15__lane25_strm1_data        = 'h1234_5678 ;
    std__pe15__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe15__lane26_strm0_cntl        = 'd0         ;
    std__pe15__lane26_strm0_data        = 'h1234_5678 ;
    std__pe15__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe15__lane26_strm1_cntl        = 'd0         ;
    std__pe15__lane26_strm1_data        = 'h1234_5678 ;
    std__pe15__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe15__lane27_strm0_cntl        = 'd0         ;
    std__pe15__lane27_strm0_data        = 'h1234_5678 ;
    std__pe15__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe15__lane27_strm1_cntl        = 'd0         ;
    std__pe15__lane27_strm1_data        = 'h1234_5678 ;
    std__pe15__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe15__lane28_strm0_cntl        = 'd0         ;
    std__pe15__lane28_strm0_data        = 'h1234_5678 ;
    std__pe15__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe15__lane28_strm1_cntl        = 'd0         ;
    std__pe15__lane28_strm1_data        = 'h1234_5678 ;
    std__pe15__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe15__lane29_strm0_cntl        = 'd0         ;
    std__pe15__lane29_strm0_data        = 'h1234_5678 ;
    std__pe15__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe15__lane29_strm1_cntl        = 'd0         ;
    std__pe15__lane29_strm1_data        = 'h1234_5678 ;
    std__pe15__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe15__lane30_strm0_cntl        = 'd0         ;
    std__pe15__lane30_strm0_data        = 'h1234_5678 ;
    std__pe15__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe15__lane30_strm1_cntl        = 'd0         ;
    std__pe15__lane30_strm1_data        = 'h1234_5678 ;
    std__pe15__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe15__lane31_strm0_cntl        = 'd0         ;
    std__pe15__lane31_strm0_data        = 'h1234_5678 ;
    std__pe15__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe15__lane31_strm1_cntl        = 'd0         ;
    std__pe15__lane31_strm1_data        = 'h1234_5678 ;
    std__pe15__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe16__lane0_strm0_cntl        = 'd0         ;
    std__pe16__lane0_strm0_data        = 'h1234_5678 ;
    std__pe16__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe16__lane0_strm1_cntl        = 'd0         ;
    std__pe16__lane0_strm1_data        = 'h1234_5678 ;
    std__pe16__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe16__lane1_strm0_cntl        = 'd0         ;
    std__pe16__lane1_strm0_data        = 'h1234_5678 ;
    std__pe16__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe16__lane1_strm1_cntl        = 'd0         ;
    std__pe16__lane1_strm1_data        = 'h1234_5678 ;
    std__pe16__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe16__lane2_strm0_cntl        = 'd0         ;
    std__pe16__lane2_strm0_data        = 'h1234_5678 ;
    std__pe16__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe16__lane2_strm1_cntl        = 'd0         ;
    std__pe16__lane2_strm1_data        = 'h1234_5678 ;
    std__pe16__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe16__lane3_strm0_cntl        = 'd0         ;
    std__pe16__lane3_strm0_data        = 'h1234_5678 ;
    std__pe16__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe16__lane3_strm1_cntl        = 'd0         ;
    std__pe16__lane3_strm1_data        = 'h1234_5678 ;
    std__pe16__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe16__lane4_strm0_cntl        = 'd0         ;
    std__pe16__lane4_strm0_data        = 'h1234_5678 ;
    std__pe16__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe16__lane4_strm1_cntl        = 'd0         ;
    std__pe16__lane4_strm1_data        = 'h1234_5678 ;
    std__pe16__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe16__lane5_strm0_cntl        = 'd0         ;
    std__pe16__lane5_strm0_data        = 'h1234_5678 ;
    std__pe16__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe16__lane5_strm1_cntl        = 'd0         ;
    std__pe16__lane5_strm1_data        = 'h1234_5678 ;
    std__pe16__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe16__lane6_strm0_cntl        = 'd0         ;
    std__pe16__lane6_strm0_data        = 'h1234_5678 ;
    std__pe16__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe16__lane6_strm1_cntl        = 'd0         ;
    std__pe16__lane6_strm1_data        = 'h1234_5678 ;
    std__pe16__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe16__lane7_strm0_cntl        = 'd0         ;
    std__pe16__lane7_strm0_data        = 'h1234_5678 ;
    std__pe16__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe16__lane7_strm1_cntl        = 'd0         ;
    std__pe16__lane7_strm1_data        = 'h1234_5678 ;
    std__pe16__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe16__lane8_strm0_cntl        = 'd0         ;
    std__pe16__lane8_strm0_data        = 'h1234_5678 ;
    std__pe16__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe16__lane8_strm1_cntl        = 'd0         ;
    std__pe16__lane8_strm1_data        = 'h1234_5678 ;
    std__pe16__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe16__lane9_strm0_cntl        = 'd0         ;
    std__pe16__lane9_strm0_data        = 'h1234_5678 ;
    std__pe16__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe16__lane9_strm1_cntl        = 'd0         ;
    std__pe16__lane9_strm1_data        = 'h1234_5678 ;
    std__pe16__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe16__lane10_strm0_cntl        = 'd0         ;
    std__pe16__lane10_strm0_data        = 'h1234_5678 ;
    std__pe16__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe16__lane10_strm1_cntl        = 'd0         ;
    std__pe16__lane10_strm1_data        = 'h1234_5678 ;
    std__pe16__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe16__lane11_strm0_cntl        = 'd0         ;
    std__pe16__lane11_strm0_data        = 'h1234_5678 ;
    std__pe16__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe16__lane11_strm1_cntl        = 'd0         ;
    std__pe16__lane11_strm1_data        = 'h1234_5678 ;
    std__pe16__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe16__lane12_strm0_cntl        = 'd0         ;
    std__pe16__lane12_strm0_data        = 'h1234_5678 ;
    std__pe16__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe16__lane12_strm1_cntl        = 'd0         ;
    std__pe16__lane12_strm1_data        = 'h1234_5678 ;
    std__pe16__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe16__lane13_strm0_cntl        = 'd0         ;
    std__pe16__lane13_strm0_data        = 'h1234_5678 ;
    std__pe16__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe16__lane13_strm1_cntl        = 'd0         ;
    std__pe16__lane13_strm1_data        = 'h1234_5678 ;
    std__pe16__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe16__lane14_strm0_cntl        = 'd0         ;
    std__pe16__lane14_strm0_data        = 'h1234_5678 ;
    std__pe16__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe16__lane14_strm1_cntl        = 'd0         ;
    std__pe16__lane14_strm1_data        = 'h1234_5678 ;
    std__pe16__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe16__lane15_strm0_cntl        = 'd0         ;
    std__pe16__lane15_strm0_data        = 'h1234_5678 ;
    std__pe16__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe16__lane15_strm1_cntl        = 'd0         ;
    std__pe16__lane15_strm1_data        = 'h1234_5678 ;
    std__pe16__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe16__lane16_strm0_cntl        = 'd0         ;
    std__pe16__lane16_strm0_data        = 'h1234_5678 ;
    std__pe16__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe16__lane16_strm1_cntl        = 'd0         ;
    std__pe16__lane16_strm1_data        = 'h1234_5678 ;
    std__pe16__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe16__lane17_strm0_cntl        = 'd0         ;
    std__pe16__lane17_strm0_data        = 'h1234_5678 ;
    std__pe16__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe16__lane17_strm1_cntl        = 'd0         ;
    std__pe16__lane17_strm1_data        = 'h1234_5678 ;
    std__pe16__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe16__lane18_strm0_cntl        = 'd0         ;
    std__pe16__lane18_strm0_data        = 'h1234_5678 ;
    std__pe16__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe16__lane18_strm1_cntl        = 'd0         ;
    std__pe16__lane18_strm1_data        = 'h1234_5678 ;
    std__pe16__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe16__lane19_strm0_cntl        = 'd0         ;
    std__pe16__lane19_strm0_data        = 'h1234_5678 ;
    std__pe16__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe16__lane19_strm1_cntl        = 'd0         ;
    std__pe16__lane19_strm1_data        = 'h1234_5678 ;
    std__pe16__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe16__lane20_strm0_cntl        = 'd0         ;
    std__pe16__lane20_strm0_data        = 'h1234_5678 ;
    std__pe16__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe16__lane20_strm1_cntl        = 'd0         ;
    std__pe16__lane20_strm1_data        = 'h1234_5678 ;
    std__pe16__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe16__lane21_strm0_cntl        = 'd0         ;
    std__pe16__lane21_strm0_data        = 'h1234_5678 ;
    std__pe16__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe16__lane21_strm1_cntl        = 'd0         ;
    std__pe16__lane21_strm1_data        = 'h1234_5678 ;
    std__pe16__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe16__lane22_strm0_cntl        = 'd0         ;
    std__pe16__lane22_strm0_data        = 'h1234_5678 ;
    std__pe16__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe16__lane22_strm1_cntl        = 'd0         ;
    std__pe16__lane22_strm1_data        = 'h1234_5678 ;
    std__pe16__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe16__lane23_strm0_cntl        = 'd0         ;
    std__pe16__lane23_strm0_data        = 'h1234_5678 ;
    std__pe16__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe16__lane23_strm1_cntl        = 'd0         ;
    std__pe16__lane23_strm1_data        = 'h1234_5678 ;
    std__pe16__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe16__lane24_strm0_cntl        = 'd0         ;
    std__pe16__lane24_strm0_data        = 'h1234_5678 ;
    std__pe16__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe16__lane24_strm1_cntl        = 'd0         ;
    std__pe16__lane24_strm1_data        = 'h1234_5678 ;
    std__pe16__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe16__lane25_strm0_cntl        = 'd0         ;
    std__pe16__lane25_strm0_data        = 'h1234_5678 ;
    std__pe16__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe16__lane25_strm1_cntl        = 'd0         ;
    std__pe16__lane25_strm1_data        = 'h1234_5678 ;
    std__pe16__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe16__lane26_strm0_cntl        = 'd0         ;
    std__pe16__lane26_strm0_data        = 'h1234_5678 ;
    std__pe16__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe16__lane26_strm1_cntl        = 'd0         ;
    std__pe16__lane26_strm1_data        = 'h1234_5678 ;
    std__pe16__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe16__lane27_strm0_cntl        = 'd0         ;
    std__pe16__lane27_strm0_data        = 'h1234_5678 ;
    std__pe16__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe16__lane27_strm1_cntl        = 'd0         ;
    std__pe16__lane27_strm1_data        = 'h1234_5678 ;
    std__pe16__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe16__lane28_strm0_cntl        = 'd0         ;
    std__pe16__lane28_strm0_data        = 'h1234_5678 ;
    std__pe16__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe16__lane28_strm1_cntl        = 'd0         ;
    std__pe16__lane28_strm1_data        = 'h1234_5678 ;
    std__pe16__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe16__lane29_strm0_cntl        = 'd0         ;
    std__pe16__lane29_strm0_data        = 'h1234_5678 ;
    std__pe16__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe16__lane29_strm1_cntl        = 'd0         ;
    std__pe16__lane29_strm1_data        = 'h1234_5678 ;
    std__pe16__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe16__lane30_strm0_cntl        = 'd0         ;
    std__pe16__lane30_strm0_data        = 'h1234_5678 ;
    std__pe16__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe16__lane30_strm1_cntl        = 'd0         ;
    std__pe16__lane30_strm1_data        = 'h1234_5678 ;
    std__pe16__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe16__lane31_strm0_cntl        = 'd0         ;
    std__pe16__lane31_strm0_data        = 'h1234_5678 ;
    std__pe16__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe16__lane31_strm1_cntl        = 'd0         ;
    std__pe16__lane31_strm1_data        = 'h1234_5678 ;
    std__pe16__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe17__lane0_strm0_cntl        = 'd0         ;
    std__pe17__lane0_strm0_data        = 'h1234_5678 ;
    std__pe17__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe17__lane0_strm1_cntl        = 'd0         ;
    std__pe17__lane0_strm1_data        = 'h1234_5678 ;
    std__pe17__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe17__lane1_strm0_cntl        = 'd0         ;
    std__pe17__lane1_strm0_data        = 'h1234_5678 ;
    std__pe17__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe17__lane1_strm1_cntl        = 'd0         ;
    std__pe17__lane1_strm1_data        = 'h1234_5678 ;
    std__pe17__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe17__lane2_strm0_cntl        = 'd0         ;
    std__pe17__lane2_strm0_data        = 'h1234_5678 ;
    std__pe17__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe17__lane2_strm1_cntl        = 'd0         ;
    std__pe17__lane2_strm1_data        = 'h1234_5678 ;
    std__pe17__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe17__lane3_strm0_cntl        = 'd0         ;
    std__pe17__lane3_strm0_data        = 'h1234_5678 ;
    std__pe17__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe17__lane3_strm1_cntl        = 'd0         ;
    std__pe17__lane3_strm1_data        = 'h1234_5678 ;
    std__pe17__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe17__lane4_strm0_cntl        = 'd0         ;
    std__pe17__lane4_strm0_data        = 'h1234_5678 ;
    std__pe17__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe17__lane4_strm1_cntl        = 'd0         ;
    std__pe17__lane4_strm1_data        = 'h1234_5678 ;
    std__pe17__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe17__lane5_strm0_cntl        = 'd0         ;
    std__pe17__lane5_strm0_data        = 'h1234_5678 ;
    std__pe17__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe17__lane5_strm1_cntl        = 'd0         ;
    std__pe17__lane5_strm1_data        = 'h1234_5678 ;
    std__pe17__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe17__lane6_strm0_cntl        = 'd0         ;
    std__pe17__lane6_strm0_data        = 'h1234_5678 ;
    std__pe17__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe17__lane6_strm1_cntl        = 'd0         ;
    std__pe17__lane6_strm1_data        = 'h1234_5678 ;
    std__pe17__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe17__lane7_strm0_cntl        = 'd0         ;
    std__pe17__lane7_strm0_data        = 'h1234_5678 ;
    std__pe17__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe17__lane7_strm1_cntl        = 'd0         ;
    std__pe17__lane7_strm1_data        = 'h1234_5678 ;
    std__pe17__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe17__lane8_strm0_cntl        = 'd0         ;
    std__pe17__lane8_strm0_data        = 'h1234_5678 ;
    std__pe17__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe17__lane8_strm1_cntl        = 'd0         ;
    std__pe17__lane8_strm1_data        = 'h1234_5678 ;
    std__pe17__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe17__lane9_strm0_cntl        = 'd0         ;
    std__pe17__lane9_strm0_data        = 'h1234_5678 ;
    std__pe17__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe17__lane9_strm1_cntl        = 'd0         ;
    std__pe17__lane9_strm1_data        = 'h1234_5678 ;
    std__pe17__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe17__lane10_strm0_cntl        = 'd0         ;
    std__pe17__lane10_strm0_data        = 'h1234_5678 ;
    std__pe17__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe17__lane10_strm1_cntl        = 'd0         ;
    std__pe17__lane10_strm1_data        = 'h1234_5678 ;
    std__pe17__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe17__lane11_strm0_cntl        = 'd0         ;
    std__pe17__lane11_strm0_data        = 'h1234_5678 ;
    std__pe17__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe17__lane11_strm1_cntl        = 'd0         ;
    std__pe17__lane11_strm1_data        = 'h1234_5678 ;
    std__pe17__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe17__lane12_strm0_cntl        = 'd0         ;
    std__pe17__lane12_strm0_data        = 'h1234_5678 ;
    std__pe17__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe17__lane12_strm1_cntl        = 'd0         ;
    std__pe17__lane12_strm1_data        = 'h1234_5678 ;
    std__pe17__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe17__lane13_strm0_cntl        = 'd0         ;
    std__pe17__lane13_strm0_data        = 'h1234_5678 ;
    std__pe17__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe17__lane13_strm1_cntl        = 'd0         ;
    std__pe17__lane13_strm1_data        = 'h1234_5678 ;
    std__pe17__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe17__lane14_strm0_cntl        = 'd0         ;
    std__pe17__lane14_strm0_data        = 'h1234_5678 ;
    std__pe17__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe17__lane14_strm1_cntl        = 'd0         ;
    std__pe17__lane14_strm1_data        = 'h1234_5678 ;
    std__pe17__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe17__lane15_strm0_cntl        = 'd0         ;
    std__pe17__lane15_strm0_data        = 'h1234_5678 ;
    std__pe17__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe17__lane15_strm1_cntl        = 'd0         ;
    std__pe17__lane15_strm1_data        = 'h1234_5678 ;
    std__pe17__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe17__lane16_strm0_cntl        = 'd0         ;
    std__pe17__lane16_strm0_data        = 'h1234_5678 ;
    std__pe17__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe17__lane16_strm1_cntl        = 'd0         ;
    std__pe17__lane16_strm1_data        = 'h1234_5678 ;
    std__pe17__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe17__lane17_strm0_cntl        = 'd0         ;
    std__pe17__lane17_strm0_data        = 'h1234_5678 ;
    std__pe17__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe17__lane17_strm1_cntl        = 'd0         ;
    std__pe17__lane17_strm1_data        = 'h1234_5678 ;
    std__pe17__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe17__lane18_strm0_cntl        = 'd0         ;
    std__pe17__lane18_strm0_data        = 'h1234_5678 ;
    std__pe17__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe17__lane18_strm1_cntl        = 'd0         ;
    std__pe17__lane18_strm1_data        = 'h1234_5678 ;
    std__pe17__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe17__lane19_strm0_cntl        = 'd0         ;
    std__pe17__lane19_strm0_data        = 'h1234_5678 ;
    std__pe17__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe17__lane19_strm1_cntl        = 'd0         ;
    std__pe17__lane19_strm1_data        = 'h1234_5678 ;
    std__pe17__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe17__lane20_strm0_cntl        = 'd0         ;
    std__pe17__lane20_strm0_data        = 'h1234_5678 ;
    std__pe17__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe17__lane20_strm1_cntl        = 'd0         ;
    std__pe17__lane20_strm1_data        = 'h1234_5678 ;
    std__pe17__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe17__lane21_strm0_cntl        = 'd0         ;
    std__pe17__lane21_strm0_data        = 'h1234_5678 ;
    std__pe17__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe17__lane21_strm1_cntl        = 'd0         ;
    std__pe17__lane21_strm1_data        = 'h1234_5678 ;
    std__pe17__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe17__lane22_strm0_cntl        = 'd0         ;
    std__pe17__lane22_strm0_data        = 'h1234_5678 ;
    std__pe17__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe17__lane22_strm1_cntl        = 'd0         ;
    std__pe17__lane22_strm1_data        = 'h1234_5678 ;
    std__pe17__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe17__lane23_strm0_cntl        = 'd0         ;
    std__pe17__lane23_strm0_data        = 'h1234_5678 ;
    std__pe17__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe17__lane23_strm1_cntl        = 'd0         ;
    std__pe17__lane23_strm1_data        = 'h1234_5678 ;
    std__pe17__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe17__lane24_strm0_cntl        = 'd0         ;
    std__pe17__lane24_strm0_data        = 'h1234_5678 ;
    std__pe17__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe17__lane24_strm1_cntl        = 'd0         ;
    std__pe17__lane24_strm1_data        = 'h1234_5678 ;
    std__pe17__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe17__lane25_strm0_cntl        = 'd0         ;
    std__pe17__lane25_strm0_data        = 'h1234_5678 ;
    std__pe17__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe17__lane25_strm1_cntl        = 'd0         ;
    std__pe17__lane25_strm1_data        = 'h1234_5678 ;
    std__pe17__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe17__lane26_strm0_cntl        = 'd0         ;
    std__pe17__lane26_strm0_data        = 'h1234_5678 ;
    std__pe17__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe17__lane26_strm1_cntl        = 'd0         ;
    std__pe17__lane26_strm1_data        = 'h1234_5678 ;
    std__pe17__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe17__lane27_strm0_cntl        = 'd0         ;
    std__pe17__lane27_strm0_data        = 'h1234_5678 ;
    std__pe17__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe17__lane27_strm1_cntl        = 'd0         ;
    std__pe17__lane27_strm1_data        = 'h1234_5678 ;
    std__pe17__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe17__lane28_strm0_cntl        = 'd0         ;
    std__pe17__lane28_strm0_data        = 'h1234_5678 ;
    std__pe17__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe17__lane28_strm1_cntl        = 'd0         ;
    std__pe17__lane28_strm1_data        = 'h1234_5678 ;
    std__pe17__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe17__lane29_strm0_cntl        = 'd0         ;
    std__pe17__lane29_strm0_data        = 'h1234_5678 ;
    std__pe17__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe17__lane29_strm1_cntl        = 'd0         ;
    std__pe17__lane29_strm1_data        = 'h1234_5678 ;
    std__pe17__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe17__lane30_strm0_cntl        = 'd0         ;
    std__pe17__lane30_strm0_data        = 'h1234_5678 ;
    std__pe17__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe17__lane30_strm1_cntl        = 'd0         ;
    std__pe17__lane30_strm1_data        = 'h1234_5678 ;
    std__pe17__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe17__lane31_strm0_cntl        = 'd0         ;
    std__pe17__lane31_strm0_data        = 'h1234_5678 ;
    std__pe17__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe17__lane31_strm1_cntl        = 'd0         ;
    std__pe17__lane31_strm1_data        = 'h1234_5678 ;
    std__pe17__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe18__lane0_strm0_cntl        = 'd0         ;
    std__pe18__lane0_strm0_data        = 'h1234_5678 ;
    std__pe18__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe18__lane0_strm1_cntl        = 'd0         ;
    std__pe18__lane0_strm1_data        = 'h1234_5678 ;
    std__pe18__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe18__lane1_strm0_cntl        = 'd0         ;
    std__pe18__lane1_strm0_data        = 'h1234_5678 ;
    std__pe18__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe18__lane1_strm1_cntl        = 'd0         ;
    std__pe18__lane1_strm1_data        = 'h1234_5678 ;
    std__pe18__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe18__lane2_strm0_cntl        = 'd0         ;
    std__pe18__lane2_strm0_data        = 'h1234_5678 ;
    std__pe18__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe18__lane2_strm1_cntl        = 'd0         ;
    std__pe18__lane2_strm1_data        = 'h1234_5678 ;
    std__pe18__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe18__lane3_strm0_cntl        = 'd0         ;
    std__pe18__lane3_strm0_data        = 'h1234_5678 ;
    std__pe18__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe18__lane3_strm1_cntl        = 'd0         ;
    std__pe18__lane3_strm1_data        = 'h1234_5678 ;
    std__pe18__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe18__lane4_strm0_cntl        = 'd0         ;
    std__pe18__lane4_strm0_data        = 'h1234_5678 ;
    std__pe18__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe18__lane4_strm1_cntl        = 'd0         ;
    std__pe18__lane4_strm1_data        = 'h1234_5678 ;
    std__pe18__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe18__lane5_strm0_cntl        = 'd0         ;
    std__pe18__lane5_strm0_data        = 'h1234_5678 ;
    std__pe18__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe18__lane5_strm1_cntl        = 'd0         ;
    std__pe18__lane5_strm1_data        = 'h1234_5678 ;
    std__pe18__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe18__lane6_strm0_cntl        = 'd0         ;
    std__pe18__lane6_strm0_data        = 'h1234_5678 ;
    std__pe18__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe18__lane6_strm1_cntl        = 'd0         ;
    std__pe18__lane6_strm1_data        = 'h1234_5678 ;
    std__pe18__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe18__lane7_strm0_cntl        = 'd0         ;
    std__pe18__lane7_strm0_data        = 'h1234_5678 ;
    std__pe18__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe18__lane7_strm1_cntl        = 'd0         ;
    std__pe18__lane7_strm1_data        = 'h1234_5678 ;
    std__pe18__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe18__lane8_strm0_cntl        = 'd0         ;
    std__pe18__lane8_strm0_data        = 'h1234_5678 ;
    std__pe18__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe18__lane8_strm1_cntl        = 'd0         ;
    std__pe18__lane8_strm1_data        = 'h1234_5678 ;
    std__pe18__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe18__lane9_strm0_cntl        = 'd0         ;
    std__pe18__lane9_strm0_data        = 'h1234_5678 ;
    std__pe18__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe18__lane9_strm1_cntl        = 'd0         ;
    std__pe18__lane9_strm1_data        = 'h1234_5678 ;
    std__pe18__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe18__lane10_strm0_cntl        = 'd0         ;
    std__pe18__lane10_strm0_data        = 'h1234_5678 ;
    std__pe18__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe18__lane10_strm1_cntl        = 'd0         ;
    std__pe18__lane10_strm1_data        = 'h1234_5678 ;
    std__pe18__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe18__lane11_strm0_cntl        = 'd0         ;
    std__pe18__lane11_strm0_data        = 'h1234_5678 ;
    std__pe18__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe18__lane11_strm1_cntl        = 'd0         ;
    std__pe18__lane11_strm1_data        = 'h1234_5678 ;
    std__pe18__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe18__lane12_strm0_cntl        = 'd0         ;
    std__pe18__lane12_strm0_data        = 'h1234_5678 ;
    std__pe18__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe18__lane12_strm1_cntl        = 'd0         ;
    std__pe18__lane12_strm1_data        = 'h1234_5678 ;
    std__pe18__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe18__lane13_strm0_cntl        = 'd0         ;
    std__pe18__lane13_strm0_data        = 'h1234_5678 ;
    std__pe18__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe18__lane13_strm1_cntl        = 'd0         ;
    std__pe18__lane13_strm1_data        = 'h1234_5678 ;
    std__pe18__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe18__lane14_strm0_cntl        = 'd0         ;
    std__pe18__lane14_strm0_data        = 'h1234_5678 ;
    std__pe18__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe18__lane14_strm1_cntl        = 'd0         ;
    std__pe18__lane14_strm1_data        = 'h1234_5678 ;
    std__pe18__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe18__lane15_strm0_cntl        = 'd0         ;
    std__pe18__lane15_strm0_data        = 'h1234_5678 ;
    std__pe18__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe18__lane15_strm1_cntl        = 'd0         ;
    std__pe18__lane15_strm1_data        = 'h1234_5678 ;
    std__pe18__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe18__lane16_strm0_cntl        = 'd0         ;
    std__pe18__lane16_strm0_data        = 'h1234_5678 ;
    std__pe18__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe18__lane16_strm1_cntl        = 'd0         ;
    std__pe18__lane16_strm1_data        = 'h1234_5678 ;
    std__pe18__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe18__lane17_strm0_cntl        = 'd0         ;
    std__pe18__lane17_strm0_data        = 'h1234_5678 ;
    std__pe18__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe18__lane17_strm1_cntl        = 'd0         ;
    std__pe18__lane17_strm1_data        = 'h1234_5678 ;
    std__pe18__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe18__lane18_strm0_cntl        = 'd0         ;
    std__pe18__lane18_strm0_data        = 'h1234_5678 ;
    std__pe18__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe18__lane18_strm1_cntl        = 'd0         ;
    std__pe18__lane18_strm1_data        = 'h1234_5678 ;
    std__pe18__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe18__lane19_strm0_cntl        = 'd0         ;
    std__pe18__lane19_strm0_data        = 'h1234_5678 ;
    std__pe18__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe18__lane19_strm1_cntl        = 'd0         ;
    std__pe18__lane19_strm1_data        = 'h1234_5678 ;
    std__pe18__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe18__lane20_strm0_cntl        = 'd0         ;
    std__pe18__lane20_strm0_data        = 'h1234_5678 ;
    std__pe18__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe18__lane20_strm1_cntl        = 'd0         ;
    std__pe18__lane20_strm1_data        = 'h1234_5678 ;
    std__pe18__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe18__lane21_strm0_cntl        = 'd0         ;
    std__pe18__lane21_strm0_data        = 'h1234_5678 ;
    std__pe18__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe18__lane21_strm1_cntl        = 'd0         ;
    std__pe18__lane21_strm1_data        = 'h1234_5678 ;
    std__pe18__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe18__lane22_strm0_cntl        = 'd0         ;
    std__pe18__lane22_strm0_data        = 'h1234_5678 ;
    std__pe18__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe18__lane22_strm1_cntl        = 'd0         ;
    std__pe18__lane22_strm1_data        = 'h1234_5678 ;
    std__pe18__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe18__lane23_strm0_cntl        = 'd0         ;
    std__pe18__lane23_strm0_data        = 'h1234_5678 ;
    std__pe18__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe18__lane23_strm1_cntl        = 'd0         ;
    std__pe18__lane23_strm1_data        = 'h1234_5678 ;
    std__pe18__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe18__lane24_strm0_cntl        = 'd0         ;
    std__pe18__lane24_strm0_data        = 'h1234_5678 ;
    std__pe18__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe18__lane24_strm1_cntl        = 'd0         ;
    std__pe18__lane24_strm1_data        = 'h1234_5678 ;
    std__pe18__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe18__lane25_strm0_cntl        = 'd0         ;
    std__pe18__lane25_strm0_data        = 'h1234_5678 ;
    std__pe18__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe18__lane25_strm1_cntl        = 'd0         ;
    std__pe18__lane25_strm1_data        = 'h1234_5678 ;
    std__pe18__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe18__lane26_strm0_cntl        = 'd0         ;
    std__pe18__lane26_strm0_data        = 'h1234_5678 ;
    std__pe18__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe18__lane26_strm1_cntl        = 'd0         ;
    std__pe18__lane26_strm1_data        = 'h1234_5678 ;
    std__pe18__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe18__lane27_strm0_cntl        = 'd0         ;
    std__pe18__lane27_strm0_data        = 'h1234_5678 ;
    std__pe18__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe18__lane27_strm1_cntl        = 'd0         ;
    std__pe18__lane27_strm1_data        = 'h1234_5678 ;
    std__pe18__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe18__lane28_strm0_cntl        = 'd0         ;
    std__pe18__lane28_strm0_data        = 'h1234_5678 ;
    std__pe18__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe18__lane28_strm1_cntl        = 'd0         ;
    std__pe18__lane28_strm1_data        = 'h1234_5678 ;
    std__pe18__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe18__lane29_strm0_cntl        = 'd0         ;
    std__pe18__lane29_strm0_data        = 'h1234_5678 ;
    std__pe18__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe18__lane29_strm1_cntl        = 'd0         ;
    std__pe18__lane29_strm1_data        = 'h1234_5678 ;
    std__pe18__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe18__lane30_strm0_cntl        = 'd0         ;
    std__pe18__lane30_strm0_data        = 'h1234_5678 ;
    std__pe18__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe18__lane30_strm1_cntl        = 'd0         ;
    std__pe18__lane30_strm1_data        = 'h1234_5678 ;
    std__pe18__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe18__lane31_strm0_cntl        = 'd0         ;
    std__pe18__lane31_strm0_data        = 'h1234_5678 ;
    std__pe18__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe18__lane31_strm1_cntl        = 'd0         ;
    std__pe18__lane31_strm1_data        = 'h1234_5678 ;
    std__pe18__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe19__lane0_strm0_cntl        = 'd0         ;
    std__pe19__lane0_strm0_data        = 'h1234_5678 ;
    std__pe19__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe19__lane0_strm1_cntl        = 'd0         ;
    std__pe19__lane0_strm1_data        = 'h1234_5678 ;
    std__pe19__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe19__lane1_strm0_cntl        = 'd0         ;
    std__pe19__lane1_strm0_data        = 'h1234_5678 ;
    std__pe19__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe19__lane1_strm1_cntl        = 'd0         ;
    std__pe19__lane1_strm1_data        = 'h1234_5678 ;
    std__pe19__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe19__lane2_strm0_cntl        = 'd0         ;
    std__pe19__lane2_strm0_data        = 'h1234_5678 ;
    std__pe19__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe19__lane2_strm1_cntl        = 'd0         ;
    std__pe19__lane2_strm1_data        = 'h1234_5678 ;
    std__pe19__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe19__lane3_strm0_cntl        = 'd0         ;
    std__pe19__lane3_strm0_data        = 'h1234_5678 ;
    std__pe19__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe19__lane3_strm1_cntl        = 'd0         ;
    std__pe19__lane3_strm1_data        = 'h1234_5678 ;
    std__pe19__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe19__lane4_strm0_cntl        = 'd0         ;
    std__pe19__lane4_strm0_data        = 'h1234_5678 ;
    std__pe19__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe19__lane4_strm1_cntl        = 'd0         ;
    std__pe19__lane4_strm1_data        = 'h1234_5678 ;
    std__pe19__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe19__lane5_strm0_cntl        = 'd0         ;
    std__pe19__lane5_strm0_data        = 'h1234_5678 ;
    std__pe19__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe19__lane5_strm1_cntl        = 'd0         ;
    std__pe19__lane5_strm1_data        = 'h1234_5678 ;
    std__pe19__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe19__lane6_strm0_cntl        = 'd0         ;
    std__pe19__lane6_strm0_data        = 'h1234_5678 ;
    std__pe19__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe19__lane6_strm1_cntl        = 'd0         ;
    std__pe19__lane6_strm1_data        = 'h1234_5678 ;
    std__pe19__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe19__lane7_strm0_cntl        = 'd0         ;
    std__pe19__lane7_strm0_data        = 'h1234_5678 ;
    std__pe19__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe19__lane7_strm1_cntl        = 'd0         ;
    std__pe19__lane7_strm1_data        = 'h1234_5678 ;
    std__pe19__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe19__lane8_strm0_cntl        = 'd0         ;
    std__pe19__lane8_strm0_data        = 'h1234_5678 ;
    std__pe19__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe19__lane8_strm1_cntl        = 'd0         ;
    std__pe19__lane8_strm1_data        = 'h1234_5678 ;
    std__pe19__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe19__lane9_strm0_cntl        = 'd0         ;
    std__pe19__lane9_strm0_data        = 'h1234_5678 ;
    std__pe19__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe19__lane9_strm1_cntl        = 'd0         ;
    std__pe19__lane9_strm1_data        = 'h1234_5678 ;
    std__pe19__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe19__lane10_strm0_cntl        = 'd0         ;
    std__pe19__lane10_strm0_data        = 'h1234_5678 ;
    std__pe19__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe19__lane10_strm1_cntl        = 'd0         ;
    std__pe19__lane10_strm1_data        = 'h1234_5678 ;
    std__pe19__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe19__lane11_strm0_cntl        = 'd0         ;
    std__pe19__lane11_strm0_data        = 'h1234_5678 ;
    std__pe19__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe19__lane11_strm1_cntl        = 'd0         ;
    std__pe19__lane11_strm1_data        = 'h1234_5678 ;
    std__pe19__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe19__lane12_strm0_cntl        = 'd0         ;
    std__pe19__lane12_strm0_data        = 'h1234_5678 ;
    std__pe19__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe19__lane12_strm1_cntl        = 'd0         ;
    std__pe19__lane12_strm1_data        = 'h1234_5678 ;
    std__pe19__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe19__lane13_strm0_cntl        = 'd0         ;
    std__pe19__lane13_strm0_data        = 'h1234_5678 ;
    std__pe19__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe19__lane13_strm1_cntl        = 'd0         ;
    std__pe19__lane13_strm1_data        = 'h1234_5678 ;
    std__pe19__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe19__lane14_strm0_cntl        = 'd0         ;
    std__pe19__lane14_strm0_data        = 'h1234_5678 ;
    std__pe19__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe19__lane14_strm1_cntl        = 'd0         ;
    std__pe19__lane14_strm1_data        = 'h1234_5678 ;
    std__pe19__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe19__lane15_strm0_cntl        = 'd0         ;
    std__pe19__lane15_strm0_data        = 'h1234_5678 ;
    std__pe19__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe19__lane15_strm1_cntl        = 'd0         ;
    std__pe19__lane15_strm1_data        = 'h1234_5678 ;
    std__pe19__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe19__lane16_strm0_cntl        = 'd0         ;
    std__pe19__lane16_strm0_data        = 'h1234_5678 ;
    std__pe19__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe19__lane16_strm1_cntl        = 'd0         ;
    std__pe19__lane16_strm1_data        = 'h1234_5678 ;
    std__pe19__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe19__lane17_strm0_cntl        = 'd0         ;
    std__pe19__lane17_strm0_data        = 'h1234_5678 ;
    std__pe19__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe19__lane17_strm1_cntl        = 'd0         ;
    std__pe19__lane17_strm1_data        = 'h1234_5678 ;
    std__pe19__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe19__lane18_strm0_cntl        = 'd0         ;
    std__pe19__lane18_strm0_data        = 'h1234_5678 ;
    std__pe19__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe19__lane18_strm1_cntl        = 'd0         ;
    std__pe19__lane18_strm1_data        = 'h1234_5678 ;
    std__pe19__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe19__lane19_strm0_cntl        = 'd0         ;
    std__pe19__lane19_strm0_data        = 'h1234_5678 ;
    std__pe19__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe19__lane19_strm1_cntl        = 'd0         ;
    std__pe19__lane19_strm1_data        = 'h1234_5678 ;
    std__pe19__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe19__lane20_strm0_cntl        = 'd0         ;
    std__pe19__lane20_strm0_data        = 'h1234_5678 ;
    std__pe19__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe19__lane20_strm1_cntl        = 'd0         ;
    std__pe19__lane20_strm1_data        = 'h1234_5678 ;
    std__pe19__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe19__lane21_strm0_cntl        = 'd0         ;
    std__pe19__lane21_strm0_data        = 'h1234_5678 ;
    std__pe19__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe19__lane21_strm1_cntl        = 'd0         ;
    std__pe19__lane21_strm1_data        = 'h1234_5678 ;
    std__pe19__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe19__lane22_strm0_cntl        = 'd0         ;
    std__pe19__lane22_strm0_data        = 'h1234_5678 ;
    std__pe19__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe19__lane22_strm1_cntl        = 'd0         ;
    std__pe19__lane22_strm1_data        = 'h1234_5678 ;
    std__pe19__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe19__lane23_strm0_cntl        = 'd0         ;
    std__pe19__lane23_strm0_data        = 'h1234_5678 ;
    std__pe19__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe19__lane23_strm1_cntl        = 'd0         ;
    std__pe19__lane23_strm1_data        = 'h1234_5678 ;
    std__pe19__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe19__lane24_strm0_cntl        = 'd0         ;
    std__pe19__lane24_strm0_data        = 'h1234_5678 ;
    std__pe19__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe19__lane24_strm1_cntl        = 'd0         ;
    std__pe19__lane24_strm1_data        = 'h1234_5678 ;
    std__pe19__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe19__lane25_strm0_cntl        = 'd0         ;
    std__pe19__lane25_strm0_data        = 'h1234_5678 ;
    std__pe19__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe19__lane25_strm1_cntl        = 'd0         ;
    std__pe19__lane25_strm1_data        = 'h1234_5678 ;
    std__pe19__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe19__lane26_strm0_cntl        = 'd0         ;
    std__pe19__lane26_strm0_data        = 'h1234_5678 ;
    std__pe19__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe19__lane26_strm1_cntl        = 'd0         ;
    std__pe19__lane26_strm1_data        = 'h1234_5678 ;
    std__pe19__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe19__lane27_strm0_cntl        = 'd0         ;
    std__pe19__lane27_strm0_data        = 'h1234_5678 ;
    std__pe19__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe19__lane27_strm1_cntl        = 'd0         ;
    std__pe19__lane27_strm1_data        = 'h1234_5678 ;
    std__pe19__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe19__lane28_strm0_cntl        = 'd0         ;
    std__pe19__lane28_strm0_data        = 'h1234_5678 ;
    std__pe19__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe19__lane28_strm1_cntl        = 'd0         ;
    std__pe19__lane28_strm1_data        = 'h1234_5678 ;
    std__pe19__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe19__lane29_strm0_cntl        = 'd0         ;
    std__pe19__lane29_strm0_data        = 'h1234_5678 ;
    std__pe19__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe19__lane29_strm1_cntl        = 'd0         ;
    std__pe19__lane29_strm1_data        = 'h1234_5678 ;
    std__pe19__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe19__lane30_strm0_cntl        = 'd0         ;
    std__pe19__lane30_strm0_data        = 'h1234_5678 ;
    std__pe19__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe19__lane30_strm1_cntl        = 'd0         ;
    std__pe19__lane30_strm1_data        = 'h1234_5678 ;
    std__pe19__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe19__lane31_strm0_cntl        = 'd0         ;
    std__pe19__lane31_strm0_data        = 'h1234_5678 ;
    std__pe19__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe19__lane31_strm1_cntl        = 'd0         ;
    std__pe19__lane31_strm1_data        = 'h1234_5678 ;
    std__pe19__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe20__lane0_strm0_cntl        = 'd0         ;
    std__pe20__lane0_strm0_data        = 'h1234_5678 ;
    std__pe20__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe20__lane0_strm1_cntl        = 'd0         ;
    std__pe20__lane0_strm1_data        = 'h1234_5678 ;
    std__pe20__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe20__lane1_strm0_cntl        = 'd0         ;
    std__pe20__lane1_strm0_data        = 'h1234_5678 ;
    std__pe20__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe20__lane1_strm1_cntl        = 'd0         ;
    std__pe20__lane1_strm1_data        = 'h1234_5678 ;
    std__pe20__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe20__lane2_strm0_cntl        = 'd0         ;
    std__pe20__lane2_strm0_data        = 'h1234_5678 ;
    std__pe20__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe20__lane2_strm1_cntl        = 'd0         ;
    std__pe20__lane2_strm1_data        = 'h1234_5678 ;
    std__pe20__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe20__lane3_strm0_cntl        = 'd0         ;
    std__pe20__lane3_strm0_data        = 'h1234_5678 ;
    std__pe20__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe20__lane3_strm1_cntl        = 'd0         ;
    std__pe20__lane3_strm1_data        = 'h1234_5678 ;
    std__pe20__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe20__lane4_strm0_cntl        = 'd0         ;
    std__pe20__lane4_strm0_data        = 'h1234_5678 ;
    std__pe20__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe20__lane4_strm1_cntl        = 'd0         ;
    std__pe20__lane4_strm1_data        = 'h1234_5678 ;
    std__pe20__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe20__lane5_strm0_cntl        = 'd0         ;
    std__pe20__lane5_strm0_data        = 'h1234_5678 ;
    std__pe20__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe20__lane5_strm1_cntl        = 'd0         ;
    std__pe20__lane5_strm1_data        = 'h1234_5678 ;
    std__pe20__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe20__lane6_strm0_cntl        = 'd0         ;
    std__pe20__lane6_strm0_data        = 'h1234_5678 ;
    std__pe20__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe20__lane6_strm1_cntl        = 'd0         ;
    std__pe20__lane6_strm1_data        = 'h1234_5678 ;
    std__pe20__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe20__lane7_strm0_cntl        = 'd0         ;
    std__pe20__lane7_strm0_data        = 'h1234_5678 ;
    std__pe20__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe20__lane7_strm1_cntl        = 'd0         ;
    std__pe20__lane7_strm1_data        = 'h1234_5678 ;
    std__pe20__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe20__lane8_strm0_cntl        = 'd0         ;
    std__pe20__lane8_strm0_data        = 'h1234_5678 ;
    std__pe20__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe20__lane8_strm1_cntl        = 'd0         ;
    std__pe20__lane8_strm1_data        = 'h1234_5678 ;
    std__pe20__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe20__lane9_strm0_cntl        = 'd0         ;
    std__pe20__lane9_strm0_data        = 'h1234_5678 ;
    std__pe20__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe20__lane9_strm1_cntl        = 'd0         ;
    std__pe20__lane9_strm1_data        = 'h1234_5678 ;
    std__pe20__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe20__lane10_strm0_cntl        = 'd0         ;
    std__pe20__lane10_strm0_data        = 'h1234_5678 ;
    std__pe20__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe20__lane10_strm1_cntl        = 'd0         ;
    std__pe20__lane10_strm1_data        = 'h1234_5678 ;
    std__pe20__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe20__lane11_strm0_cntl        = 'd0         ;
    std__pe20__lane11_strm0_data        = 'h1234_5678 ;
    std__pe20__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe20__lane11_strm1_cntl        = 'd0         ;
    std__pe20__lane11_strm1_data        = 'h1234_5678 ;
    std__pe20__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe20__lane12_strm0_cntl        = 'd0         ;
    std__pe20__lane12_strm0_data        = 'h1234_5678 ;
    std__pe20__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe20__lane12_strm1_cntl        = 'd0         ;
    std__pe20__lane12_strm1_data        = 'h1234_5678 ;
    std__pe20__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe20__lane13_strm0_cntl        = 'd0         ;
    std__pe20__lane13_strm0_data        = 'h1234_5678 ;
    std__pe20__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe20__lane13_strm1_cntl        = 'd0         ;
    std__pe20__lane13_strm1_data        = 'h1234_5678 ;
    std__pe20__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe20__lane14_strm0_cntl        = 'd0         ;
    std__pe20__lane14_strm0_data        = 'h1234_5678 ;
    std__pe20__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe20__lane14_strm1_cntl        = 'd0         ;
    std__pe20__lane14_strm1_data        = 'h1234_5678 ;
    std__pe20__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe20__lane15_strm0_cntl        = 'd0         ;
    std__pe20__lane15_strm0_data        = 'h1234_5678 ;
    std__pe20__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe20__lane15_strm1_cntl        = 'd0         ;
    std__pe20__lane15_strm1_data        = 'h1234_5678 ;
    std__pe20__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe20__lane16_strm0_cntl        = 'd0         ;
    std__pe20__lane16_strm0_data        = 'h1234_5678 ;
    std__pe20__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe20__lane16_strm1_cntl        = 'd0         ;
    std__pe20__lane16_strm1_data        = 'h1234_5678 ;
    std__pe20__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe20__lane17_strm0_cntl        = 'd0         ;
    std__pe20__lane17_strm0_data        = 'h1234_5678 ;
    std__pe20__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe20__lane17_strm1_cntl        = 'd0         ;
    std__pe20__lane17_strm1_data        = 'h1234_5678 ;
    std__pe20__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe20__lane18_strm0_cntl        = 'd0         ;
    std__pe20__lane18_strm0_data        = 'h1234_5678 ;
    std__pe20__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe20__lane18_strm1_cntl        = 'd0         ;
    std__pe20__lane18_strm1_data        = 'h1234_5678 ;
    std__pe20__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe20__lane19_strm0_cntl        = 'd0         ;
    std__pe20__lane19_strm0_data        = 'h1234_5678 ;
    std__pe20__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe20__lane19_strm1_cntl        = 'd0         ;
    std__pe20__lane19_strm1_data        = 'h1234_5678 ;
    std__pe20__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe20__lane20_strm0_cntl        = 'd0         ;
    std__pe20__lane20_strm0_data        = 'h1234_5678 ;
    std__pe20__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe20__lane20_strm1_cntl        = 'd0         ;
    std__pe20__lane20_strm1_data        = 'h1234_5678 ;
    std__pe20__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe20__lane21_strm0_cntl        = 'd0         ;
    std__pe20__lane21_strm0_data        = 'h1234_5678 ;
    std__pe20__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe20__lane21_strm1_cntl        = 'd0         ;
    std__pe20__lane21_strm1_data        = 'h1234_5678 ;
    std__pe20__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe20__lane22_strm0_cntl        = 'd0         ;
    std__pe20__lane22_strm0_data        = 'h1234_5678 ;
    std__pe20__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe20__lane22_strm1_cntl        = 'd0         ;
    std__pe20__lane22_strm1_data        = 'h1234_5678 ;
    std__pe20__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe20__lane23_strm0_cntl        = 'd0         ;
    std__pe20__lane23_strm0_data        = 'h1234_5678 ;
    std__pe20__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe20__lane23_strm1_cntl        = 'd0         ;
    std__pe20__lane23_strm1_data        = 'h1234_5678 ;
    std__pe20__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe20__lane24_strm0_cntl        = 'd0         ;
    std__pe20__lane24_strm0_data        = 'h1234_5678 ;
    std__pe20__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe20__lane24_strm1_cntl        = 'd0         ;
    std__pe20__lane24_strm1_data        = 'h1234_5678 ;
    std__pe20__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe20__lane25_strm0_cntl        = 'd0         ;
    std__pe20__lane25_strm0_data        = 'h1234_5678 ;
    std__pe20__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe20__lane25_strm1_cntl        = 'd0         ;
    std__pe20__lane25_strm1_data        = 'h1234_5678 ;
    std__pe20__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe20__lane26_strm0_cntl        = 'd0         ;
    std__pe20__lane26_strm0_data        = 'h1234_5678 ;
    std__pe20__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe20__lane26_strm1_cntl        = 'd0         ;
    std__pe20__lane26_strm1_data        = 'h1234_5678 ;
    std__pe20__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe20__lane27_strm0_cntl        = 'd0         ;
    std__pe20__lane27_strm0_data        = 'h1234_5678 ;
    std__pe20__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe20__lane27_strm1_cntl        = 'd0         ;
    std__pe20__lane27_strm1_data        = 'h1234_5678 ;
    std__pe20__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe20__lane28_strm0_cntl        = 'd0         ;
    std__pe20__lane28_strm0_data        = 'h1234_5678 ;
    std__pe20__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe20__lane28_strm1_cntl        = 'd0         ;
    std__pe20__lane28_strm1_data        = 'h1234_5678 ;
    std__pe20__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe20__lane29_strm0_cntl        = 'd0         ;
    std__pe20__lane29_strm0_data        = 'h1234_5678 ;
    std__pe20__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe20__lane29_strm1_cntl        = 'd0         ;
    std__pe20__lane29_strm1_data        = 'h1234_5678 ;
    std__pe20__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe20__lane30_strm0_cntl        = 'd0         ;
    std__pe20__lane30_strm0_data        = 'h1234_5678 ;
    std__pe20__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe20__lane30_strm1_cntl        = 'd0         ;
    std__pe20__lane30_strm1_data        = 'h1234_5678 ;
    std__pe20__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe20__lane31_strm0_cntl        = 'd0         ;
    std__pe20__lane31_strm0_data        = 'h1234_5678 ;
    std__pe20__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe20__lane31_strm1_cntl        = 'd0         ;
    std__pe20__lane31_strm1_data        = 'h1234_5678 ;
    std__pe20__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe21__lane0_strm0_cntl        = 'd0         ;
    std__pe21__lane0_strm0_data        = 'h1234_5678 ;
    std__pe21__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe21__lane0_strm1_cntl        = 'd0         ;
    std__pe21__lane0_strm1_data        = 'h1234_5678 ;
    std__pe21__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe21__lane1_strm0_cntl        = 'd0         ;
    std__pe21__lane1_strm0_data        = 'h1234_5678 ;
    std__pe21__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe21__lane1_strm1_cntl        = 'd0         ;
    std__pe21__lane1_strm1_data        = 'h1234_5678 ;
    std__pe21__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe21__lane2_strm0_cntl        = 'd0         ;
    std__pe21__lane2_strm0_data        = 'h1234_5678 ;
    std__pe21__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe21__lane2_strm1_cntl        = 'd0         ;
    std__pe21__lane2_strm1_data        = 'h1234_5678 ;
    std__pe21__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe21__lane3_strm0_cntl        = 'd0         ;
    std__pe21__lane3_strm0_data        = 'h1234_5678 ;
    std__pe21__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe21__lane3_strm1_cntl        = 'd0         ;
    std__pe21__lane3_strm1_data        = 'h1234_5678 ;
    std__pe21__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe21__lane4_strm0_cntl        = 'd0         ;
    std__pe21__lane4_strm0_data        = 'h1234_5678 ;
    std__pe21__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe21__lane4_strm1_cntl        = 'd0         ;
    std__pe21__lane4_strm1_data        = 'h1234_5678 ;
    std__pe21__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe21__lane5_strm0_cntl        = 'd0         ;
    std__pe21__lane5_strm0_data        = 'h1234_5678 ;
    std__pe21__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe21__lane5_strm1_cntl        = 'd0         ;
    std__pe21__lane5_strm1_data        = 'h1234_5678 ;
    std__pe21__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe21__lane6_strm0_cntl        = 'd0         ;
    std__pe21__lane6_strm0_data        = 'h1234_5678 ;
    std__pe21__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe21__lane6_strm1_cntl        = 'd0         ;
    std__pe21__lane6_strm1_data        = 'h1234_5678 ;
    std__pe21__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe21__lane7_strm0_cntl        = 'd0         ;
    std__pe21__lane7_strm0_data        = 'h1234_5678 ;
    std__pe21__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe21__lane7_strm1_cntl        = 'd0         ;
    std__pe21__lane7_strm1_data        = 'h1234_5678 ;
    std__pe21__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe21__lane8_strm0_cntl        = 'd0         ;
    std__pe21__lane8_strm0_data        = 'h1234_5678 ;
    std__pe21__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe21__lane8_strm1_cntl        = 'd0         ;
    std__pe21__lane8_strm1_data        = 'h1234_5678 ;
    std__pe21__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe21__lane9_strm0_cntl        = 'd0         ;
    std__pe21__lane9_strm0_data        = 'h1234_5678 ;
    std__pe21__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe21__lane9_strm1_cntl        = 'd0         ;
    std__pe21__lane9_strm1_data        = 'h1234_5678 ;
    std__pe21__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe21__lane10_strm0_cntl        = 'd0         ;
    std__pe21__lane10_strm0_data        = 'h1234_5678 ;
    std__pe21__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe21__lane10_strm1_cntl        = 'd0         ;
    std__pe21__lane10_strm1_data        = 'h1234_5678 ;
    std__pe21__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe21__lane11_strm0_cntl        = 'd0         ;
    std__pe21__lane11_strm0_data        = 'h1234_5678 ;
    std__pe21__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe21__lane11_strm1_cntl        = 'd0         ;
    std__pe21__lane11_strm1_data        = 'h1234_5678 ;
    std__pe21__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe21__lane12_strm0_cntl        = 'd0         ;
    std__pe21__lane12_strm0_data        = 'h1234_5678 ;
    std__pe21__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe21__lane12_strm1_cntl        = 'd0         ;
    std__pe21__lane12_strm1_data        = 'h1234_5678 ;
    std__pe21__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe21__lane13_strm0_cntl        = 'd0         ;
    std__pe21__lane13_strm0_data        = 'h1234_5678 ;
    std__pe21__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe21__lane13_strm1_cntl        = 'd0         ;
    std__pe21__lane13_strm1_data        = 'h1234_5678 ;
    std__pe21__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe21__lane14_strm0_cntl        = 'd0         ;
    std__pe21__lane14_strm0_data        = 'h1234_5678 ;
    std__pe21__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe21__lane14_strm1_cntl        = 'd0         ;
    std__pe21__lane14_strm1_data        = 'h1234_5678 ;
    std__pe21__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe21__lane15_strm0_cntl        = 'd0         ;
    std__pe21__lane15_strm0_data        = 'h1234_5678 ;
    std__pe21__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe21__lane15_strm1_cntl        = 'd0         ;
    std__pe21__lane15_strm1_data        = 'h1234_5678 ;
    std__pe21__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe21__lane16_strm0_cntl        = 'd0         ;
    std__pe21__lane16_strm0_data        = 'h1234_5678 ;
    std__pe21__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe21__lane16_strm1_cntl        = 'd0         ;
    std__pe21__lane16_strm1_data        = 'h1234_5678 ;
    std__pe21__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe21__lane17_strm0_cntl        = 'd0         ;
    std__pe21__lane17_strm0_data        = 'h1234_5678 ;
    std__pe21__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe21__lane17_strm1_cntl        = 'd0         ;
    std__pe21__lane17_strm1_data        = 'h1234_5678 ;
    std__pe21__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe21__lane18_strm0_cntl        = 'd0         ;
    std__pe21__lane18_strm0_data        = 'h1234_5678 ;
    std__pe21__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe21__lane18_strm1_cntl        = 'd0         ;
    std__pe21__lane18_strm1_data        = 'h1234_5678 ;
    std__pe21__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe21__lane19_strm0_cntl        = 'd0         ;
    std__pe21__lane19_strm0_data        = 'h1234_5678 ;
    std__pe21__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe21__lane19_strm1_cntl        = 'd0         ;
    std__pe21__lane19_strm1_data        = 'h1234_5678 ;
    std__pe21__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe21__lane20_strm0_cntl        = 'd0         ;
    std__pe21__lane20_strm0_data        = 'h1234_5678 ;
    std__pe21__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe21__lane20_strm1_cntl        = 'd0         ;
    std__pe21__lane20_strm1_data        = 'h1234_5678 ;
    std__pe21__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe21__lane21_strm0_cntl        = 'd0         ;
    std__pe21__lane21_strm0_data        = 'h1234_5678 ;
    std__pe21__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe21__lane21_strm1_cntl        = 'd0         ;
    std__pe21__lane21_strm1_data        = 'h1234_5678 ;
    std__pe21__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe21__lane22_strm0_cntl        = 'd0         ;
    std__pe21__lane22_strm0_data        = 'h1234_5678 ;
    std__pe21__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe21__lane22_strm1_cntl        = 'd0         ;
    std__pe21__lane22_strm1_data        = 'h1234_5678 ;
    std__pe21__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe21__lane23_strm0_cntl        = 'd0         ;
    std__pe21__lane23_strm0_data        = 'h1234_5678 ;
    std__pe21__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe21__lane23_strm1_cntl        = 'd0         ;
    std__pe21__lane23_strm1_data        = 'h1234_5678 ;
    std__pe21__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe21__lane24_strm0_cntl        = 'd0         ;
    std__pe21__lane24_strm0_data        = 'h1234_5678 ;
    std__pe21__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe21__lane24_strm1_cntl        = 'd0         ;
    std__pe21__lane24_strm1_data        = 'h1234_5678 ;
    std__pe21__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe21__lane25_strm0_cntl        = 'd0         ;
    std__pe21__lane25_strm0_data        = 'h1234_5678 ;
    std__pe21__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe21__lane25_strm1_cntl        = 'd0         ;
    std__pe21__lane25_strm1_data        = 'h1234_5678 ;
    std__pe21__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe21__lane26_strm0_cntl        = 'd0         ;
    std__pe21__lane26_strm0_data        = 'h1234_5678 ;
    std__pe21__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe21__lane26_strm1_cntl        = 'd0         ;
    std__pe21__lane26_strm1_data        = 'h1234_5678 ;
    std__pe21__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe21__lane27_strm0_cntl        = 'd0         ;
    std__pe21__lane27_strm0_data        = 'h1234_5678 ;
    std__pe21__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe21__lane27_strm1_cntl        = 'd0         ;
    std__pe21__lane27_strm1_data        = 'h1234_5678 ;
    std__pe21__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe21__lane28_strm0_cntl        = 'd0         ;
    std__pe21__lane28_strm0_data        = 'h1234_5678 ;
    std__pe21__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe21__lane28_strm1_cntl        = 'd0         ;
    std__pe21__lane28_strm1_data        = 'h1234_5678 ;
    std__pe21__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe21__lane29_strm0_cntl        = 'd0         ;
    std__pe21__lane29_strm0_data        = 'h1234_5678 ;
    std__pe21__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe21__lane29_strm1_cntl        = 'd0         ;
    std__pe21__lane29_strm1_data        = 'h1234_5678 ;
    std__pe21__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe21__lane30_strm0_cntl        = 'd0         ;
    std__pe21__lane30_strm0_data        = 'h1234_5678 ;
    std__pe21__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe21__lane30_strm1_cntl        = 'd0         ;
    std__pe21__lane30_strm1_data        = 'h1234_5678 ;
    std__pe21__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe21__lane31_strm0_cntl        = 'd0         ;
    std__pe21__lane31_strm0_data        = 'h1234_5678 ;
    std__pe21__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe21__lane31_strm1_cntl        = 'd0         ;
    std__pe21__lane31_strm1_data        = 'h1234_5678 ;
    std__pe21__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe22__lane0_strm0_cntl        = 'd0         ;
    std__pe22__lane0_strm0_data        = 'h1234_5678 ;
    std__pe22__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe22__lane0_strm1_cntl        = 'd0         ;
    std__pe22__lane0_strm1_data        = 'h1234_5678 ;
    std__pe22__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe22__lane1_strm0_cntl        = 'd0         ;
    std__pe22__lane1_strm0_data        = 'h1234_5678 ;
    std__pe22__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe22__lane1_strm1_cntl        = 'd0         ;
    std__pe22__lane1_strm1_data        = 'h1234_5678 ;
    std__pe22__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe22__lane2_strm0_cntl        = 'd0         ;
    std__pe22__lane2_strm0_data        = 'h1234_5678 ;
    std__pe22__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe22__lane2_strm1_cntl        = 'd0         ;
    std__pe22__lane2_strm1_data        = 'h1234_5678 ;
    std__pe22__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe22__lane3_strm0_cntl        = 'd0         ;
    std__pe22__lane3_strm0_data        = 'h1234_5678 ;
    std__pe22__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe22__lane3_strm1_cntl        = 'd0         ;
    std__pe22__lane3_strm1_data        = 'h1234_5678 ;
    std__pe22__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe22__lane4_strm0_cntl        = 'd0         ;
    std__pe22__lane4_strm0_data        = 'h1234_5678 ;
    std__pe22__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe22__lane4_strm1_cntl        = 'd0         ;
    std__pe22__lane4_strm1_data        = 'h1234_5678 ;
    std__pe22__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe22__lane5_strm0_cntl        = 'd0         ;
    std__pe22__lane5_strm0_data        = 'h1234_5678 ;
    std__pe22__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe22__lane5_strm1_cntl        = 'd0         ;
    std__pe22__lane5_strm1_data        = 'h1234_5678 ;
    std__pe22__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe22__lane6_strm0_cntl        = 'd0         ;
    std__pe22__lane6_strm0_data        = 'h1234_5678 ;
    std__pe22__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe22__lane6_strm1_cntl        = 'd0         ;
    std__pe22__lane6_strm1_data        = 'h1234_5678 ;
    std__pe22__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe22__lane7_strm0_cntl        = 'd0         ;
    std__pe22__lane7_strm0_data        = 'h1234_5678 ;
    std__pe22__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe22__lane7_strm1_cntl        = 'd0         ;
    std__pe22__lane7_strm1_data        = 'h1234_5678 ;
    std__pe22__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe22__lane8_strm0_cntl        = 'd0         ;
    std__pe22__lane8_strm0_data        = 'h1234_5678 ;
    std__pe22__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe22__lane8_strm1_cntl        = 'd0         ;
    std__pe22__lane8_strm1_data        = 'h1234_5678 ;
    std__pe22__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe22__lane9_strm0_cntl        = 'd0         ;
    std__pe22__lane9_strm0_data        = 'h1234_5678 ;
    std__pe22__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe22__lane9_strm1_cntl        = 'd0         ;
    std__pe22__lane9_strm1_data        = 'h1234_5678 ;
    std__pe22__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe22__lane10_strm0_cntl        = 'd0         ;
    std__pe22__lane10_strm0_data        = 'h1234_5678 ;
    std__pe22__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe22__lane10_strm1_cntl        = 'd0         ;
    std__pe22__lane10_strm1_data        = 'h1234_5678 ;
    std__pe22__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe22__lane11_strm0_cntl        = 'd0         ;
    std__pe22__lane11_strm0_data        = 'h1234_5678 ;
    std__pe22__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe22__lane11_strm1_cntl        = 'd0         ;
    std__pe22__lane11_strm1_data        = 'h1234_5678 ;
    std__pe22__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe22__lane12_strm0_cntl        = 'd0         ;
    std__pe22__lane12_strm0_data        = 'h1234_5678 ;
    std__pe22__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe22__lane12_strm1_cntl        = 'd0         ;
    std__pe22__lane12_strm1_data        = 'h1234_5678 ;
    std__pe22__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe22__lane13_strm0_cntl        = 'd0         ;
    std__pe22__lane13_strm0_data        = 'h1234_5678 ;
    std__pe22__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe22__lane13_strm1_cntl        = 'd0         ;
    std__pe22__lane13_strm1_data        = 'h1234_5678 ;
    std__pe22__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe22__lane14_strm0_cntl        = 'd0         ;
    std__pe22__lane14_strm0_data        = 'h1234_5678 ;
    std__pe22__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe22__lane14_strm1_cntl        = 'd0         ;
    std__pe22__lane14_strm1_data        = 'h1234_5678 ;
    std__pe22__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe22__lane15_strm0_cntl        = 'd0         ;
    std__pe22__lane15_strm0_data        = 'h1234_5678 ;
    std__pe22__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe22__lane15_strm1_cntl        = 'd0         ;
    std__pe22__lane15_strm1_data        = 'h1234_5678 ;
    std__pe22__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe22__lane16_strm0_cntl        = 'd0         ;
    std__pe22__lane16_strm0_data        = 'h1234_5678 ;
    std__pe22__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe22__lane16_strm1_cntl        = 'd0         ;
    std__pe22__lane16_strm1_data        = 'h1234_5678 ;
    std__pe22__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe22__lane17_strm0_cntl        = 'd0         ;
    std__pe22__lane17_strm0_data        = 'h1234_5678 ;
    std__pe22__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe22__lane17_strm1_cntl        = 'd0         ;
    std__pe22__lane17_strm1_data        = 'h1234_5678 ;
    std__pe22__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe22__lane18_strm0_cntl        = 'd0         ;
    std__pe22__lane18_strm0_data        = 'h1234_5678 ;
    std__pe22__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe22__lane18_strm1_cntl        = 'd0         ;
    std__pe22__lane18_strm1_data        = 'h1234_5678 ;
    std__pe22__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe22__lane19_strm0_cntl        = 'd0         ;
    std__pe22__lane19_strm0_data        = 'h1234_5678 ;
    std__pe22__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe22__lane19_strm1_cntl        = 'd0         ;
    std__pe22__lane19_strm1_data        = 'h1234_5678 ;
    std__pe22__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe22__lane20_strm0_cntl        = 'd0         ;
    std__pe22__lane20_strm0_data        = 'h1234_5678 ;
    std__pe22__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe22__lane20_strm1_cntl        = 'd0         ;
    std__pe22__lane20_strm1_data        = 'h1234_5678 ;
    std__pe22__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe22__lane21_strm0_cntl        = 'd0         ;
    std__pe22__lane21_strm0_data        = 'h1234_5678 ;
    std__pe22__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe22__lane21_strm1_cntl        = 'd0         ;
    std__pe22__lane21_strm1_data        = 'h1234_5678 ;
    std__pe22__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe22__lane22_strm0_cntl        = 'd0         ;
    std__pe22__lane22_strm0_data        = 'h1234_5678 ;
    std__pe22__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe22__lane22_strm1_cntl        = 'd0         ;
    std__pe22__lane22_strm1_data        = 'h1234_5678 ;
    std__pe22__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe22__lane23_strm0_cntl        = 'd0         ;
    std__pe22__lane23_strm0_data        = 'h1234_5678 ;
    std__pe22__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe22__lane23_strm1_cntl        = 'd0         ;
    std__pe22__lane23_strm1_data        = 'h1234_5678 ;
    std__pe22__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe22__lane24_strm0_cntl        = 'd0         ;
    std__pe22__lane24_strm0_data        = 'h1234_5678 ;
    std__pe22__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe22__lane24_strm1_cntl        = 'd0         ;
    std__pe22__lane24_strm1_data        = 'h1234_5678 ;
    std__pe22__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe22__lane25_strm0_cntl        = 'd0         ;
    std__pe22__lane25_strm0_data        = 'h1234_5678 ;
    std__pe22__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe22__lane25_strm1_cntl        = 'd0         ;
    std__pe22__lane25_strm1_data        = 'h1234_5678 ;
    std__pe22__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe22__lane26_strm0_cntl        = 'd0         ;
    std__pe22__lane26_strm0_data        = 'h1234_5678 ;
    std__pe22__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe22__lane26_strm1_cntl        = 'd0         ;
    std__pe22__lane26_strm1_data        = 'h1234_5678 ;
    std__pe22__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe22__lane27_strm0_cntl        = 'd0         ;
    std__pe22__lane27_strm0_data        = 'h1234_5678 ;
    std__pe22__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe22__lane27_strm1_cntl        = 'd0         ;
    std__pe22__lane27_strm1_data        = 'h1234_5678 ;
    std__pe22__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe22__lane28_strm0_cntl        = 'd0         ;
    std__pe22__lane28_strm0_data        = 'h1234_5678 ;
    std__pe22__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe22__lane28_strm1_cntl        = 'd0         ;
    std__pe22__lane28_strm1_data        = 'h1234_5678 ;
    std__pe22__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe22__lane29_strm0_cntl        = 'd0         ;
    std__pe22__lane29_strm0_data        = 'h1234_5678 ;
    std__pe22__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe22__lane29_strm1_cntl        = 'd0         ;
    std__pe22__lane29_strm1_data        = 'h1234_5678 ;
    std__pe22__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe22__lane30_strm0_cntl        = 'd0         ;
    std__pe22__lane30_strm0_data        = 'h1234_5678 ;
    std__pe22__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe22__lane30_strm1_cntl        = 'd0         ;
    std__pe22__lane30_strm1_data        = 'h1234_5678 ;
    std__pe22__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe22__lane31_strm0_cntl        = 'd0         ;
    std__pe22__lane31_strm0_data        = 'h1234_5678 ;
    std__pe22__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe22__lane31_strm1_cntl        = 'd0         ;
    std__pe22__lane31_strm1_data        = 'h1234_5678 ;
    std__pe22__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe23__lane0_strm0_cntl        = 'd0         ;
    std__pe23__lane0_strm0_data        = 'h1234_5678 ;
    std__pe23__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe23__lane0_strm1_cntl        = 'd0         ;
    std__pe23__lane0_strm1_data        = 'h1234_5678 ;
    std__pe23__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe23__lane1_strm0_cntl        = 'd0         ;
    std__pe23__lane1_strm0_data        = 'h1234_5678 ;
    std__pe23__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe23__lane1_strm1_cntl        = 'd0         ;
    std__pe23__lane1_strm1_data        = 'h1234_5678 ;
    std__pe23__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe23__lane2_strm0_cntl        = 'd0         ;
    std__pe23__lane2_strm0_data        = 'h1234_5678 ;
    std__pe23__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe23__lane2_strm1_cntl        = 'd0         ;
    std__pe23__lane2_strm1_data        = 'h1234_5678 ;
    std__pe23__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe23__lane3_strm0_cntl        = 'd0         ;
    std__pe23__lane3_strm0_data        = 'h1234_5678 ;
    std__pe23__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe23__lane3_strm1_cntl        = 'd0         ;
    std__pe23__lane3_strm1_data        = 'h1234_5678 ;
    std__pe23__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe23__lane4_strm0_cntl        = 'd0         ;
    std__pe23__lane4_strm0_data        = 'h1234_5678 ;
    std__pe23__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe23__lane4_strm1_cntl        = 'd0         ;
    std__pe23__lane4_strm1_data        = 'h1234_5678 ;
    std__pe23__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe23__lane5_strm0_cntl        = 'd0         ;
    std__pe23__lane5_strm0_data        = 'h1234_5678 ;
    std__pe23__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe23__lane5_strm1_cntl        = 'd0         ;
    std__pe23__lane5_strm1_data        = 'h1234_5678 ;
    std__pe23__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe23__lane6_strm0_cntl        = 'd0         ;
    std__pe23__lane6_strm0_data        = 'h1234_5678 ;
    std__pe23__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe23__lane6_strm1_cntl        = 'd0         ;
    std__pe23__lane6_strm1_data        = 'h1234_5678 ;
    std__pe23__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe23__lane7_strm0_cntl        = 'd0         ;
    std__pe23__lane7_strm0_data        = 'h1234_5678 ;
    std__pe23__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe23__lane7_strm1_cntl        = 'd0         ;
    std__pe23__lane7_strm1_data        = 'h1234_5678 ;
    std__pe23__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe23__lane8_strm0_cntl        = 'd0         ;
    std__pe23__lane8_strm0_data        = 'h1234_5678 ;
    std__pe23__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe23__lane8_strm1_cntl        = 'd0         ;
    std__pe23__lane8_strm1_data        = 'h1234_5678 ;
    std__pe23__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe23__lane9_strm0_cntl        = 'd0         ;
    std__pe23__lane9_strm0_data        = 'h1234_5678 ;
    std__pe23__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe23__lane9_strm1_cntl        = 'd0         ;
    std__pe23__lane9_strm1_data        = 'h1234_5678 ;
    std__pe23__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe23__lane10_strm0_cntl        = 'd0         ;
    std__pe23__lane10_strm0_data        = 'h1234_5678 ;
    std__pe23__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe23__lane10_strm1_cntl        = 'd0         ;
    std__pe23__lane10_strm1_data        = 'h1234_5678 ;
    std__pe23__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe23__lane11_strm0_cntl        = 'd0         ;
    std__pe23__lane11_strm0_data        = 'h1234_5678 ;
    std__pe23__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe23__lane11_strm1_cntl        = 'd0         ;
    std__pe23__lane11_strm1_data        = 'h1234_5678 ;
    std__pe23__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe23__lane12_strm0_cntl        = 'd0         ;
    std__pe23__lane12_strm0_data        = 'h1234_5678 ;
    std__pe23__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe23__lane12_strm1_cntl        = 'd0         ;
    std__pe23__lane12_strm1_data        = 'h1234_5678 ;
    std__pe23__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe23__lane13_strm0_cntl        = 'd0         ;
    std__pe23__lane13_strm0_data        = 'h1234_5678 ;
    std__pe23__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe23__lane13_strm1_cntl        = 'd0         ;
    std__pe23__lane13_strm1_data        = 'h1234_5678 ;
    std__pe23__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe23__lane14_strm0_cntl        = 'd0         ;
    std__pe23__lane14_strm0_data        = 'h1234_5678 ;
    std__pe23__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe23__lane14_strm1_cntl        = 'd0         ;
    std__pe23__lane14_strm1_data        = 'h1234_5678 ;
    std__pe23__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe23__lane15_strm0_cntl        = 'd0         ;
    std__pe23__lane15_strm0_data        = 'h1234_5678 ;
    std__pe23__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe23__lane15_strm1_cntl        = 'd0         ;
    std__pe23__lane15_strm1_data        = 'h1234_5678 ;
    std__pe23__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe23__lane16_strm0_cntl        = 'd0         ;
    std__pe23__lane16_strm0_data        = 'h1234_5678 ;
    std__pe23__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe23__lane16_strm1_cntl        = 'd0         ;
    std__pe23__lane16_strm1_data        = 'h1234_5678 ;
    std__pe23__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe23__lane17_strm0_cntl        = 'd0         ;
    std__pe23__lane17_strm0_data        = 'h1234_5678 ;
    std__pe23__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe23__lane17_strm1_cntl        = 'd0         ;
    std__pe23__lane17_strm1_data        = 'h1234_5678 ;
    std__pe23__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe23__lane18_strm0_cntl        = 'd0         ;
    std__pe23__lane18_strm0_data        = 'h1234_5678 ;
    std__pe23__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe23__lane18_strm1_cntl        = 'd0         ;
    std__pe23__lane18_strm1_data        = 'h1234_5678 ;
    std__pe23__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe23__lane19_strm0_cntl        = 'd0         ;
    std__pe23__lane19_strm0_data        = 'h1234_5678 ;
    std__pe23__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe23__lane19_strm1_cntl        = 'd0         ;
    std__pe23__lane19_strm1_data        = 'h1234_5678 ;
    std__pe23__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe23__lane20_strm0_cntl        = 'd0         ;
    std__pe23__lane20_strm0_data        = 'h1234_5678 ;
    std__pe23__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe23__lane20_strm1_cntl        = 'd0         ;
    std__pe23__lane20_strm1_data        = 'h1234_5678 ;
    std__pe23__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe23__lane21_strm0_cntl        = 'd0         ;
    std__pe23__lane21_strm0_data        = 'h1234_5678 ;
    std__pe23__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe23__lane21_strm1_cntl        = 'd0         ;
    std__pe23__lane21_strm1_data        = 'h1234_5678 ;
    std__pe23__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe23__lane22_strm0_cntl        = 'd0         ;
    std__pe23__lane22_strm0_data        = 'h1234_5678 ;
    std__pe23__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe23__lane22_strm1_cntl        = 'd0         ;
    std__pe23__lane22_strm1_data        = 'h1234_5678 ;
    std__pe23__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe23__lane23_strm0_cntl        = 'd0         ;
    std__pe23__lane23_strm0_data        = 'h1234_5678 ;
    std__pe23__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe23__lane23_strm1_cntl        = 'd0         ;
    std__pe23__lane23_strm1_data        = 'h1234_5678 ;
    std__pe23__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe23__lane24_strm0_cntl        = 'd0         ;
    std__pe23__lane24_strm0_data        = 'h1234_5678 ;
    std__pe23__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe23__lane24_strm1_cntl        = 'd0         ;
    std__pe23__lane24_strm1_data        = 'h1234_5678 ;
    std__pe23__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe23__lane25_strm0_cntl        = 'd0         ;
    std__pe23__lane25_strm0_data        = 'h1234_5678 ;
    std__pe23__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe23__lane25_strm1_cntl        = 'd0         ;
    std__pe23__lane25_strm1_data        = 'h1234_5678 ;
    std__pe23__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe23__lane26_strm0_cntl        = 'd0         ;
    std__pe23__lane26_strm0_data        = 'h1234_5678 ;
    std__pe23__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe23__lane26_strm1_cntl        = 'd0         ;
    std__pe23__lane26_strm1_data        = 'h1234_5678 ;
    std__pe23__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe23__lane27_strm0_cntl        = 'd0         ;
    std__pe23__lane27_strm0_data        = 'h1234_5678 ;
    std__pe23__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe23__lane27_strm1_cntl        = 'd0         ;
    std__pe23__lane27_strm1_data        = 'h1234_5678 ;
    std__pe23__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe23__lane28_strm0_cntl        = 'd0         ;
    std__pe23__lane28_strm0_data        = 'h1234_5678 ;
    std__pe23__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe23__lane28_strm1_cntl        = 'd0         ;
    std__pe23__lane28_strm1_data        = 'h1234_5678 ;
    std__pe23__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe23__lane29_strm0_cntl        = 'd0         ;
    std__pe23__lane29_strm0_data        = 'h1234_5678 ;
    std__pe23__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe23__lane29_strm1_cntl        = 'd0         ;
    std__pe23__lane29_strm1_data        = 'h1234_5678 ;
    std__pe23__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe23__lane30_strm0_cntl        = 'd0         ;
    std__pe23__lane30_strm0_data        = 'h1234_5678 ;
    std__pe23__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe23__lane30_strm1_cntl        = 'd0         ;
    std__pe23__lane30_strm1_data        = 'h1234_5678 ;
    std__pe23__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe23__lane31_strm0_cntl        = 'd0         ;
    std__pe23__lane31_strm0_data        = 'h1234_5678 ;
    std__pe23__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe23__lane31_strm1_cntl        = 'd0         ;
    std__pe23__lane31_strm1_data        = 'h1234_5678 ;
    std__pe23__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe24__lane0_strm0_cntl        = 'd0         ;
    std__pe24__lane0_strm0_data        = 'h1234_5678 ;
    std__pe24__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe24__lane0_strm1_cntl        = 'd0         ;
    std__pe24__lane0_strm1_data        = 'h1234_5678 ;
    std__pe24__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe24__lane1_strm0_cntl        = 'd0         ;
    std__pe24__lane1_strm0_data        = 'h1234_5678 ;
    std__pe24__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe24__lane1_strm1_cntl        = 'd0         ;
    std__pe24__lane1_strm1_data        = 'h1234_5678 ;
    std__pe24__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe24__lane2_strm0_cntl        = 'd0         ;
    std__pe24__lane2_strm0_data        = 'h1234_5678 ;
    std__pe24__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe24__lane2_strm1_cntl        = 'd0         ;
    std__pe24__lane2_strm1_data        = 'h1234_5678 ;
    std__pe24__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe24__lane3_strm0_cntl        = 'd0         ;
    std__pe24__lane3_strm0_data        = 'h1234_5678 ;
    std__pe24__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe24__lane3_strm1_cntl        = 'd0         ;
    std__pe24__lane3_strm1_data        = 'h1234_5678 ;
    std__pe24__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe24__lane4_strm0_cntl        = 'd0         ;
    std__pe24__lane4_strm0_data        = 'h1234_5678 ;
    std__pe24__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe24__lane4_strm1_cntl        = 'd0         ;
    std__pe24__lane4_strm1_data        = 'h1234_5678 ;
    std__pe24__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe24__lane5_strm0_cntl        = 'd0         ;
    std__pe24__lane5_strm0_data        = 'h1234_5678 ;
    std__pe24__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe24__lane5_strm1_cntl        = 'd0         ;
    std__pe24__lane5_strm1_data        = 'h1234_5678 ;
    std__pe24__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe24__lane6_strm0_cntl        = 'd0         ;
    std__pe24__lane6_strm0_data        = 'h1234_5678 ;
    std__pe24__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe24__lane6_strm1_cntl        = 'd0         ;
    std__pe24__lane6_strm1_data        = 'h1234_5678 ;
    std__pe24__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe24__lane7_strm0_cntl        = 'd0         ;
    std__pe24__lane7_strm0_data        = 'h1234_5678 ;
    std__pe24__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe24__lane7_strm1_cntl        = 'd0         ;
    std__pe24__lane7_strm1_data        = 'h1234_5678 ;
    std__pe24__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe24__lane8_strm0_cntl        = 'd0         ;
    std__pe24__lane8_strm0_data        = 'h1234_5678 ;
    std__pe24__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe24__lane8_strm1_cntl        = 'd0         ;
    std__pe24__lane8_strm1_data        = 'h1234_5678 ;
    std__pe24__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe24__lane9_strm0_cntl        = 'd0         ;
    std__pe24__lane9_strm0_data        = 'h1234_5678 ;
    std__pe24__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe24__lane9_strm1_cntl        = 'd0         ;
    std__pe24__lane9_strm1_data        = 'h1234_5678 ;
    std__pe24__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe24__lane10_strm0_cntl        = 'd0         ;
    std__pe24__lane10_strm0_data        = 'h1234_5678 ;
    std__pe24__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe24__lane10_strm1_cntl        = 'd0         ;
    std__pe24__lane10_strm1_data        = 'h1234_5678 ;
    std__pe24__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe24__lane11_strm0_cntl        = 'd0         ;
    std__pe24__lane11_strm0_data        = 'h1234_5678 ;
    std__pe24__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe24__lane11_strm1_cntl        = 'd0         ;
    std__pe24__lane11_strm1_data        = 'h1234_5678 ;
    std__pe24__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe24__lane12_strm0_cntl        = 'd0         ;
    std__pe24__lane12_strm0_data        = 'h1234_5678 ;
    std__pe24__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe24__lane12_strm1_cntl        = 'd0         ;
    std__pe24__lane12_strm1_data        = 'h1234_5678 ;
    std__pe24__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe24__lane13_strm0_cntl        = 'd0         ;
    std__pe24__lane13_strm0_data        = 'h1234_5678 ;
    std__pe24__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe24__lane13_strm1_cntl        = 'd0         ;
    std__pe24__lane13_strm1_data        = 'h1234_5678 ;
    std__pe24__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe24__lane14_strm0_cntl        = 'd0         ;
    std__pe24__lane14_strm0_data        = 'h1234_5678 ;
    std__pe24__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe24__lane14_strm1_cntl        = 'd0         ;
    std__pe24__lane14_strm1_data        = 'h1234_5678 ;
    std__pe24__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe24__lane15_strm0_cntl        = 'd0         ;
    std__pe24__lane15_strm0_data        = 'h1234_5678 ;
    std__pe24__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe24__lane15_strm1_cntl        = 'd0         ;
    std__pe24__lane15_strm1_data        = 'h1234_5678 ;
    std__pe24__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe24__lane16_strm0_cntl        = 'd0         ;
    std__pe24__lane16_strm0_data        = 'h1234_5678 ;
    std__pe24__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe24__lane16_strm1_cntl        = 'd0         ;
    std__pe24__lane16_strm1_data        = 'h1234_5678 ;
    std__pe24__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe24__lane17_strm0_cntl        = 'd0         ;
    std__pe24__lane17_strm0_data        = 'h1234_5678 ;
    std__pe24__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe24__lane17_strm1_cntl        = 'd0         ;
    std__pe24__lane17_strm1_data        = 'h1234_5678 ;
    std__pe24__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe24__lane18_strm0_cntl        = 'd0         ;
    std__pe24__lane18_strm0_data        = 'h1234_5678 ;
    std__pe24__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe24__lane18_strm1_cntl        = 'd0         ;
    std__pe24__lane18_strm1_data        = 'h1234_5678 ;
    std__pe24__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe24__lane19_strm0_cntl        = 'd0         ;
    std__pe24__lane19_strm0_data        = 'h1234_5678 ;
    std__pe24__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe24__lane19_strm1_cntl        = 'd0         ;
    std__pe24__lane19_strm1_data        = 'h1234_5678 ;
    std__pe24__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe24__lane20_strm0_cntl        = 'd0         ;
    std__pe24__lane20_strm0_data        = 'h1234_5678 ;
    std__pe24__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe24__lane20_strm1_cntl        = 'd0         ;
    std__pe24__lane20_strm1_data        = 'h1234_5678 ;
    std__pe24__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe24__lane21_strm0_cntl        = 'd0         ;
    std__pe24__lane21_strm0_data        = 'h1234_5678 ;
    std__pe24__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe24__lane21_strm1_cntl        = 'd0         ;
    std__pe24__lane21_strm1_data        = 'h1234_5678 ;
    std__pe24__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe24__lane22_strm0_cntl        = 'd0         ;
    std__pe24__lane22_strm0_data        = 'h1234_5678 ;
    std__pe24__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe24__lane22_strm1_cntl        = 'd0         ;
    std__pe24__lane22_strm1_data        = 'h1234_5678 ;
    std__pe24__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe24__lane23_strm0_cntl        = 'd0         ;
    std__pe24__lane23_strm0_data        = 'h1234_5678 ;
    std__pe24__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe24__lane23_strm1_cntl        = 'd0         ;
    std__pe24__lane23_strm1_data        = 'h1234_5678 ;
    std__pe24__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe24__lane24_strm0_cntl        = 'd0         ;
    std__pe24__lane24_strm0_data        = 'h1234_5678 ;
    std__pe24__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe24__lane24_strm1_cntl        = 'd0         ;
    std__pe24__lane24_strm1_data        = 'h1234_5678 ;
    std__pe24__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe24__lane25_strm0_cntl        = 'd0         ;
    std__pe24__lane25_strm0_data        = 'h1234_5678 ;
    std__pe24__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe24__lane25_strm1_cntl        = 'd0         ;
    std__pe24__lane25_strm1_data        = 'h1234_5678 ;
    std__pe24__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe24__lane26_strm0_cntl        = 'd0         ;
    std__pe24__lane26_strm0_data        = 'h1234_5678 ;
    std__pe24__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe24__lane26_strm1_cntl        = 'd0         ;
    std__pe24__lane26_strm1_data        = 'h1234_5678 ;
    std__pe24__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe24__lane27_strm0_cntl        = 'd0         ;
    std__pe24__lane27_strm0_data        = 'h1234_5678 ;
    std__pe24__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe24__lane27_strm1_cntl        = 'd0         ;
    std__pe24__lane27_strm1_data        = 'h1234_5678 ;
    std__pe24__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe24__lane28_strm0_cntl        = 'd0         ;
    std__pe24__lane28_strm0_data        = 'h1234_5678 ;
    std__pe24__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe24__lane28_strm1_cntl        = 'd0         ;
    std__pe24__lane28_strm1_data        = 'h1234_5678 ;
    std__pe24__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe24__lane29_strm0_cntl        = 'd0         ;
    std__pe24__lane29_strm0_data        = 'h1234_5678 ;
    std__pe24__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe24__lane29_strm1_cntl        = 'd0         ;
    std__pe24__lane29_strm1_data        = 'h1234_5678 ;
    std__pe24__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe24__lane30_strm0_cntl        = 'd0         ;
    std__pe24__lane30_strm0_data        = 'h1234_5678 ;
    std__pe24__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe24__lane30_strm1_cntl        = 'd0         ;
    std__pe24__lane30_strm1_data        = 'h1234_5678 ;
    std__pe24__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe24__lane31_strm0_cntl        = 'd0         ;
    std__pe24__lane31_strm0_data        = 'h1234_5678 ;
    std__pe24__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe24__lane31_strm1_cntl        = 'd0         ;
    std__pe24__lane31_strm1_data        = 'h1234_5678 ;
    std__pe24__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe25__lane0_strm0_cntl        = 'd0         ;
    std__pe25__lane0_strm0_data        = 'h1234_5678 ;
    std__pe25__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe25__lane0_strm1_cntl        = 'd0         ;
    std__pe25__lane0_strm1_data        = 'h1234_5678 ;
    std__pe25__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe25__lane1_strm0_cntl        = 'd0         ;
    std__pe25__lane1_strm0_data        = 'h1234_5678 ;
    std__pe25__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe25__lane1_strm1_cntl        = 'd0         ;
    std__pe25__lane1_strm1_data        = 'h1234_5678 ;
    std__pe25__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe25__lane2_strm0_cntl        = 'd0         ;
    std__pe25__lane2_strm0_data        = 'h1234_5678 ;
    std__pe25__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe25__lane2_strm1_cntl        = 'd0         ;
    std__pe25__lane2_strm1_data        = 'h1234_5678 ;
    std__pe25__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe25__lane3_strm0_cntl        = 'd0         ;
    std__pe25__lane3_strm0_data        = 'h1234_5678 ;
    std__pe25__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe25__lane3_strm1_cntl        = 'd0         ;
    std__pe25__lane3_strm1_data        = 'h1234_5678 ;
    std__pe25__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe25__lane4_strm0_cntl        = 'd0         ;
    std__pe25__lane4_strm0_data        = 'h1234_5678 ;
    std__pe25__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe25__lane4_strm1_cntl        = 'd0         ;
    std__pe25__lane4_strm1_data        = 'h1234_5678 ;
    std__pe25__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe25__lane5_strm0_cntl        = 'd0         ;
    std__pe25__lane5_strm0_data        = 'h1234_5678 ;
    std__pe25__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe25__lane5_strm1_cntl        = 'd0         ;
    std__pe25__lane5_strm1_data        = 'h1234_5678 ;
    std__pe25__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe25__lane6_strm0_cntl        = 'd0         ;
    std__pe25__lane6_strm0_data        = 'h1234_5678 ;
    std__pe25__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe25__lane6_strm1_cntl        = 'd0         ;
    std__pe25__lane6_strm1_data        = 'h1234_5678 ;
    std__pe25__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe25__lane7_strm0_cntl        = 'd0         ;
    std__pe25__lane7_strm0_data        = 'h1234_5678 ;
    std__pe25__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe25__lane7_strm1_cntl        = 'd0         ;
    std__pe25__lane7_strm1_data        = 'h1234_5678 ;
    std__pe25__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe25__lane8_strm0_cntl        = 'd0         ;
    std__pe25__lane8_strm0_data        = 'h1234_5678 ;
    std__pe25__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe25__lane8_strm1_cntl        = 'd0         ;
    std__pe25__lane8_strm1_data        = 'h1234_5678 ;
    std__pe25__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe25__lane9_strm0_cntl        = 'd0         ;
    std__pe25__lane9_strm0_data        = 'h1234_5678 ;
    std__pe25__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe25__lane9_strm1_cntl        = 'd0         ;
    std__pe25__lane9_strm1_data        = 'h1234_5678 ;
    std__pe25__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe25__lane10_strm0_cntl        = 'd0         ;
    std__pe25__lane10_strm0_data        = 'h1234_5678 ;
    std__pe25__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe25__lane10_strm1_cntl        = 'd0         ;
    std__pe25__lane10_strm1_data        = 'h1234_5678 ;
    std__pe25__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe25__lane11_strm0_cntl        = 'd0         ;
    std__pe25__lane11_strm0_data        = 'h1234_5678 ;
    std__pe25__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe25__lane11_strm1_cntl        = 'd0         ;
    std__pe25__lane11_strm1_data        = 'h1234_5678 ;
    std__pe25__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe25__lane12_strm0_cntl        = 'd0         ;
    std__pe25__lane12_strm0_data        = 'h1234_5678 ;
    std__pe25__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe25__lane12_strm1_cntl        = 'd0         ;
    std__pe25__lane12_strm1_data        = 'h1234_5678 ;
    std__pe25__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe25__lane13_strm0_cntl        = 'd0         ;
    std__pe25__lane13_strm0_data        = 'h1234_5678 ;
    std__pe25__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe25__lane13_strm1_cntl        = 'd0         ;
    std__pe25__lane13_strm1_data        = 'h1234_5678 ;
    std__pe25__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe25__lane14_strm0_cntl        = 'd0         ;
    std__pe25__lane14_strm0_data        = 'h1234_5678 ;
    std__pe25__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe25__lane14_strm1_cntl        = 'd0         ;
    std__pe25__lane14_strm1_data        = 'h1234_5678 ;
    std__pe25__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe25__lane15_strm0_cntl        = 'd0         ;
    std__pe25__lane15_strm0_data        = 'h1234_5678 ;
    std__pe25__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe25__lane15_strm1_cntl        = 'd0         ;
    std__pe25__lane15_strm1_data        = 'h1234_5678 ;
    std__pe25__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe25__lane16_strm0_cntl        = 'd0         ;
    std__pe25__lane16_strm0_data        = 'h1234_5678 ;
    std__pe25__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe25__lane16_strm1_cntl        = 'd0         ;
    std__pe25__lane16_strm1_data        = 'h1234_5678 ;
    std__pe25__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe25__lane17_strm0_cntl        = 'd0         ;
    std__pe25__lane17_strm0_data        = 'h1234_5678 ;
    std__pe25__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe25__lane17_strm1_cntl        = 'd0         ;
    std__pe25__lane17_strm1_data        = 'h1234_5678 ;
    std__pe25__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe25__lane18_strm0_cntl        = 'd0         ;
    std__pe25__lane18_strm0_data        = 'h1234_5678 ;
    std__pe25__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe25__lane18_strm1_cntl        = 'd0         ;
    std__pe25__lane18_strm1_data        = 'h1234_5678 ;
    std__pe25__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe25__lane19_strm0_cntl        = 'd0         ;
    std__pe25__lane19_strm0_data        = 'h1234_5678 ;
    std__pe25__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe25__lane19_strm1_cntl        = 'd0         ;
    std__pe25__lane19_strm1_data        = 'h1234_5678 ;
    std__pe25__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe25__lane20_strm0_cntl        = 'd0         ;
    std__pe25__lane20_strm0_data        = 'h1234_5678 ;
    std__pe25__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe25__lane20_strm1_cntl        = 'd0         ;
    std__pe25__lane20_strm1_data        = 'h1234_5678 ;
    std__pe25__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe25__lane21_strm0_cntl        = 'd0         ;
    std__pe25__lane21_strm0_data        = 'h1234_5678 ;
    std__pe25__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe25__lane21_strm1_cntl        = 'd0         ;
    std__pe25__lane21_strm1_data        = 'h1234_5678 ;
    std__pe25__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe25__lane22_strm0_cntl        = 'd0         ;
    std__pe25__lane22_strm0_data        = 'h1234_5678 ;
    std__pe25__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe25__lane22_strm1_cntl        = 'd0         ;
    std__pe25__lane22_strm1_data        = 'h1234_5678 ;
    std__pe25__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe25__lane23_strm0_cntl        = 'd0         ;
    std__pe25__lane23_strm0_data        = 'h1234_5678 ;
    std__pe25__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe25__lane23_strm1_cntl        = 'd0         ;
    std__pe25__lane23_strm1_data        = 'h1234_5678 ;
    std__pe25__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe25__lane24_strm0_cntl        = 'd0         ;
    std__pe25__lane24_strm0_data        = 'h1234_5678 ;
    std__pe25__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe25__lane24_strm1_cntl        = 'd0         ;
    std__pe25__lane24_strm1_data        = 'h1234_5678 ;
    std__pe25__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe25__lane25_strm0_cntl        = 'd0         ;
    std__pe25__lane25_strm0_data        = 'h1234_5678 ;
    std__pe25__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe25__lane25_strm1_cntl        = 'd0         ;
    std__pe25__lane25_strm1_data        = 'h1234_5678 ;
    std__pe25__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe25__lane26_strm0_cntl        = 'd0         ;
    std__pe25__lane26_strm0_data        = 'h1234_5678 ;
    std__pe25__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe25__lane26_strm1_cntl        = 'd0         ;
    std__pe25__lane26_strm1_data        = 'h1234_5678 ;
    std__pe25__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe25__lane27_strm0_cntl        = 'd0         ;
    std__pe25__lane27_strm0_data        = 'h1234_5678 ;
    std__pe25__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe25__lane27_strm1_cntl        = 'd0         ;
    std__pe25__lane27_strm1_data        = 'h1234_5678 ;
    std__pe25__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe25__lane28_strm0_cntl        = 'd0         ;
    std__pe25__lane28_strm0_data        = 'h1234_5678 ;
    std__pe25__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe25__lane28_strm1_cntl        = 'd0         ;
    std__pe25__lane28_strm1_data        = 'h1234_5678 ;
    std__pe25__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe25__lane29_strm0_cntl        = 'd0         ;
    std__pe25__lane29_strm0_data        = 'h1234_5678 ;
    std__pe25__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe25__lane29_strm1_cntl        = 'd0         ;
    std__pe25__lane29_strm1_data        = 'h1234_5678 ;
    std__pe25__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe25__lane30_strm0_cntl        = 'd0         ;
    std__pe25__lane30_strm0_data        = 'h1234_5678 ;
    std__pe25__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe25__lane30_strm1_cntl        = 'd0         ;
    std__pe25__lane30_strm1_data        = 'h1234_5678 ;
    std__pe25__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe25__lane31_strm0_cntl        = 'd0         ;
    std__pe25__lane31_strm0_data        = 'h1234_5678 ;
    std__pe25__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe25__lane31_strm1_cntl        = 'd0         ;
    std__pe25__lane31_strm1_data        = 'h1234_5678 ;
    std__pe25__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe26__lane0_strm0_cntl        = 'd0         ;
    std__pe26__lane0_strm0_data        = 'h1234_5678 ;
    std__pe26__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe26__lane0_strm1_cntl        = 'd0         ;
    std__pe26__lane0_strm1_data        = 'h1234_5678 ;
    std__pe26__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe26__lane1_strm0_cntl        = 'd0         ;
    std__pe26__lane1_strm0_data        = 'h1234_5678 ;
    std__pe26__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe26__lane1_strm1_cntl        = 'd0         ;
    std__pe26__lane1_strm1_data        = 'h1234_5678 ;
    std__pe26__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe26__lane2_strm0_cntl        = 'd0         ;
    std__pe26__lane2_strm0_data        = 'h1234_5678 ;
    std__pe26__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe26__lane2_strm1_cntl        = 'd0         ;
    std__pe26__lane2_strm1_data        = 'h1234_5678 ;
    std__pe26__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe26__lane3_strm0_cntl        = 'd0         ;
    std__pe26__lane3_strm0_data        = 'h1234_5678 ;
    std__pe26__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe26__lane3_strm1_cntl        = 'd0         ;
    std__pe26__lane3_strm1_data        = 'h1234_5678 ;
    std__pe26__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe26__lane4_strm0_cntl        = 'd0         ;
    std__pe26__lane4_strm0_data        = 'h1234_5678 ;
    std__pe26__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe26__lane4_strm1_cntl        = 'd0         ;
    std__pe26__lane4_strm1_data        = 'h1234_5678 ;
    std__pe26__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe26__lane5_strm0_cntl        = 'd0         ;
    std__pe26__lane5_strm0_data        = 'h1234_5678 ;
    std__pe26__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe26__lane5_strm1_cntl        = 'd0         ;
    std__pe26__lane5_strm1_data        = 'h1234_5678 ;
    std__pe26__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe26__lane6_strm0_cntl        = 'd0         ;
    std__pe26__lane6_strm0_data        = 'h1234_5678 ;
    std__pe26__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe26__lane6_strm1_cntl        = 'd0         ;
    std__pe26__lane6_strm1_data        = 'h1234_5678 ;
    std__pe26__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe26__lane7_strm0_cntl        = 'd0         ;
    std__pe26__lane7_strm0_data        = 'h1234_5678 ;
    std__pe26__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe26__lane7_strm1_cntl        = 'd0         ;
    std__pe26__lane7_strm1_data        = 'h1234_5678 ;
    std__pe26__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe26__lane8_strm0_cntl        = 'd0         ;
    std__pe26__lane8_strm0_data        = 'h1234_5678 ;
    std__pe26__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe26__lane8_strm1_cntl        = 'd0         ;
    std__pe26__lane8_strm1_data        = 'h1234_5678 ;
    std__pe26__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe26__lane9_strm0_cntl        = 'd0         ;
    std__pe26__lane9_strm0_data        = 'h1234_5678 ;
    std__pe26__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe26__lane9_strm1_cntl        = 'd0         ;
    std__pe26__lane9_strm1_data        = 'h1234_5678 ;
    std__pe26__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe26__lane10_strm0_cntl        = 'd0         ;
    std__pe26__lane10_strm0_data        = 'h1234_5678 ;
    std__pe26__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe26__lane10_strm1_cntl        = 'd0         ;
    std__pe26__lane10_strm1_data        = 'h1234_5678 ;
    std__pe26__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe26__lane11_strm0_cntl        = 'd0         ;
    std__pe26__lane11_strm0_data        = 'h1234_5678 ;
    std__pe26__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe26__lane11_strm1_cntl        = 'd0         ;
    std__pe26__lane11_strm1_data        = 'h1234_5678 ;
    std__pe26__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe26__lane12_strm0_cntl        = 'd0         ;
    std__pe26__lane12_strm0_data        = 'h1234_5678 ;
    std__pe26__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe26__lane12_strm1_cntl        = 'd0         ;
    std__pe26__lane12_strm1_data        = 'h1234_5678 ;
    std__pe26__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe26__lane13_strm0_cntl        = 'd0         ;
    std__pe26__lane13_strm0_data        = 'h1234_5678 ;
    std__pe26__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe26__lane13_strm1_cntl        = 'd0         ;
    std__pe26__lane13_strm1_data        = 'h1234_5678 ;
    std__pe26__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe26__lane14_strm0_cntl        = 'd0         ;
    std__pe26__lane14_strm0_data        = 'h1234_5678 ;
    std__pe26__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe26__lane14_strm1_cntl        = 'd0         ;
    std__pe26__lane14_strm1_data        = 'h1234_5678 ;
    std__pe26__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe26__lane15_strm0_cntl        = 'd0         ;
    std__pe26__lane15_strm0_data        = 'h1234_5678 ;
    std__pe26__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe26__lane15_strm1_cntl        = 'd0         ;
    std__pe26__lane15_strm1_data        = 'h1234_5678 ;
    std__pe26__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe26__lane16_strm0_cntl        = 'd0         ;
    std__pe26__lane16_strm0_data        = 'h1234_5678 ;
    std__pe26__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe26__lane16_strm1_cntl        = 'd0         ;
    std__pe26__lane16_strm1_data        = 'h1234_5678 ;
    std__pe26__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe26__lane17_strm0_cntl        = 'd0         ;
    std__pe26__lane17_strm0_data        = 'h1234_5678 ;
    std__pe26__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe26__lane17_strm1_cntl        = 'd0         ;
    std__pe26__lane17_strm1_data        = 'h1234_5678 ;
    std__pe26__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe26__lane18_strm0_cntl        = 'd0         ;
    std__pe26__lane18_strm0_data        = 'h1234_5678 ;
    std__pe26__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe26__lane18_strm1_cntl        = 'd0         ;
    std__pe26__lane18_strm1_data        = 'h1234_5678 ;
    std__pe26__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe26__lane19_strm0_cntl        = 'd0         ;
    std__pe26__lane19_strm0_data        = 'h1234_5678 ;
    std__pe26__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe26__lane19_strm1_cntl        = 'd0         ;
    std__pe26__lane19_strm1_data        = 'h1234_5678 ;
    std__pe26__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe26__lane20_strm0_cntl        = 'd0         ;
    std__pe26__lane20_strm0_data        = 'h1234_5678 ;
    std__pe26__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe26__lane20_strm1_cntl        = 'd0         ;
    std__pe26__lane20_strm1_data        = 'h1234_5678 ;
    std__pe26__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe26__lane21_strm0_cntl        = 'd0         ;
    std__pe26__lane21_strm0_data        = 'h1234_5678 ;
    std__pe26__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe26__lane21_strm1_cntl        = 'd0         ;
    std__pe26__lane21_strm1_data        = 'h1234_5678 ;
    std__pe26__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe26__lane22_strm0_cntl        = 'd0         ;
    std__pe26__lane22_strm0_data        = 'h1234_5678 ;
    std__pe26__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe26__lane22_strm1_cntl        = 'd0         ;
    std__pe26__lane22_strm1_data        = 'h1234_5678 ;
    std__pe26__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe26__lane23_strm0_cntl        = 'd0         ;
    std__pe26__lane23_strm0_data        = 'h1234_5678 ;
    std__pe26__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe26__lane23_strm1_cntl        = 'd0         ;
    std__pe26__lane23_strm1_data        = 'h1234_5678 ;
    std__pe26__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe26__lane24_strm0_cntl        = 'd0         ;
    std__pe26__lane24_strm0_data        = 'h1234_5678 ;
    std__pe26__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe26__lane24_strm1_cntl        = 'd0         ;
    std__pe26__lane24_strm1_data        = 'h1234_5678 ;
    std__pe26__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe26__lane25_strm0_cntl        = 'd0         ;
    std__pe26__lane25_strm0_data        = 'h1234_5678 ;
    std__pe26__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe26__lane25_strm1_cntl        = 'd0         ;
    std__pe26__lane25_strm1_data        = 'h1234_5678 ;
    std__pe26__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe26__lane26_strm0_cntl        = 'd0         ;
    std__pe26__lane26_strm0_data        = 'h1234_5678 ;
    std__pe26__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe26__lane26_strm1_cntl        = 'd0         ;
    std__pe26__lane26_strm1_data        = 'h1234_5678 ;
    std__pe26__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe26__lane27_strm0_cntl        = 'd0         ;
    std__pe26__lane27_strm0_data        = 'h1234_5678 ;
    std__pe26__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe26__lane27_strm1_cntl        = 'd0         ;
    std__pe26__lane27_strm1_data        = 'h1234_5678 ;
    std__pe26__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe26__lane28_strm0_cntl        = 'd0         ;
    std__pe26__lane28_strm0_data        = 'h1234_5678 ;
    std__pe26__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe26__lane28_strm1_cntl        = 'd0         ;
    std__pe26__lane28_strm1_data        = 'h1234_5678 ;
    std__pe26__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe26__lane29_strm0_cntl        = 'd0         ;
    std__pe26__lane29_strm0_data        = 'h1234_5678 ;
    std__pe26__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe26__lane29_strm1_cntl        = 'd0         ;
    std__pe26__lane29_strm1_data        = 'h1234_5678 ;
    std__pe26__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe26__lane30_strm0_cntl        = 'd0         ;
    std__pe26__lane30_strm0_data        = 'h1234_5678 ;
    std__pe26__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe26__lane30_strm1_cntl        = 'd0         ;
    std__pe26__lane30_strm1_data        = 'h1234_5678 ;
    std__pe26__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe26__lane31_strm0_cntl        = 'd0         ;
    std__pe26__lane31_strm0_data        = 'h1234_5678 ;
    std__pe26__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe26__lane31_strm1_cntl        = 'd0         ;
    std__pe26__lane31_strm1_data        = 'h1234_5678 ;
    std__pe26__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe27__lane0_strm0_cntl        = 'd0         ;
    std__pe27__lane0_strm0_data        = 'h1234_5678 ;
    std__pe27__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe27__lane0_strm1_cntl        = 'd0         ;
    std__pe27__lane0_strm1_data        = 'h1234_5678 ;
    std__pe27__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe27__lane1_strm0_cntl        = 'd0         ;
    std__pe27__lane1_strm0_data        = 'h1234_5678 ;
    std__pe27__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe27__lane1_strm1_cntl        = 'd0         ;
    std__pe27__lane1_strm1_data        = 'h1234_5678 ;
    std__pe27__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe27__lane2_strm0_cntl        = 'd0         ;
    std__pe27__lane2_strm0_data        = 'h1234_5678 ;
    std__pe27__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe27__lane2_strm1_cntl        = 'd0         ;
    std__pe27__lane2_strm1_data        = 'h1234_5678 ;
    std__pe27__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe27__lane3_strm0_cntl        = 'd0         ;
    std__pe27__lane3_strm0_data        = 'h1234_5678 ;
    std__pe27__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe27__lane3_strm1_cntl        = 'd0         ;
    std__pe27__lane3_strm1_data        = 'h1234_5678 ;
    std__pe27__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe27__lane4_strm0_cntl        = 'd0         ;
    std__pe27__lane4_strm0_data        = 'h1234_5678 ;
    std__pe27__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe27__lane4_strm1_cntl        = 'd0         ;
    std__pe27__lane4_strm1_data        = 'h1234_5678 ;
    std__pe27__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe27__lane5_strm0_cntl        = 'd0         ;
    std__pe27__lane5_strm0_data        = 'h1234_5678 ;
    std__pe27__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe27__lane5_strm1_cntl        = 'd0         ;
    std__pe27__lane5_strm1_data        = 'h1234_5678 ;
    std__pe27__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe27__lane6_strm0_cntl        = 'd0         ;
    std__pe27__lane6_strm0_data        = 'h1234_5678 ;
    std__pe27__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe27__lane6_strm1_cntl        = 'd0         ;
    std__pe27__lane6_strm1_data        = 'h1234_5678 ;
    std__pe27__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe27__lane7_strm0_cntl        = 'd0         ;
    std__pe27__lane7_strm0_data        = 'h1234_5678 ;
    std__pe27__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe27__lane7_strm1_cntl        = 'd0         ;
    std__pe27__lane7_strm1_data        = 'h1234_5678 ;
    std__pe27__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe27__lane8_strm0_cntl        = 'd0         ;
    std__pe27__lane8_strm0_data        = 'h1234_5678 ;
    std__pe27__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe27__lane8_strm1_cntl        = 'd0         ;
    std__pe27__lane8_strm1_data        = 'h1234_5678 ;
    std__pe27__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe27__lane9_strm0_cntl        = 'd0         ;
    std__pe27__lane9_strm0_data        = 'h1234_5678 ;
    std__pe27__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe27__lane9_strm1_cntl        = 'd0         ;
    std__pe27__lane9_strm1_data        = 'h1234_5678 ;
    std__pe27__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe27__lane10_strm0_cntl        = 'd0         ;
    std__pe27__lane10_strm0_data        = 'h1234_5678 ;
    std__pe27__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe27__lane10_strm1_cntl        = 'd0         ;
    std__pe27__lane10_strm1_data        = 'h1234_5678 ;
    std__pe27__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe27__lane11_strm0_cntl        = 'd0         ;
    std__pe27__lane11_strm0_data        = 'h1234_5678 ;
    std__pe27__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe27__lane11_strm1_cntl        = 'd0         ;
    std__pe27__lane11_strm1_data        = 'h1234_5678 ;
    std__pe27__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe27__lane12_strm0_cntl        = 'd0         ;
    std__pe27__lane12_strm0_data        = 'h1234_5678 ;
    std__pe27__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe27__lane12_strm1_cntl        = 'd0         ;
    std__pe27__lane12_strm1_data        = 'h1234_5678 ;
    std__pe27__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe27__lane13_strm0_cntl        = 'd0         ;
    std__pe27__lane13_strm0_data        = 'h1234_5678 ;
    std__pe27__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe27__lane13_strm1_cntl        = 'd0         ;
    std__pe27__lane13_strm1_data        = 'h1234_5678 ;
    std__pe27__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe27__lane14_strm0_cntl        = 'd0         ;
    std__pe27__lane14_strm0_data        = 'h1234_5678 ;
    std__pe27__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe27__lane14_strm1_cntl        = 'd0         ;
    std__pe27__lane14_strm1_data        = 'h1234_5678 ;
    std__pe27__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe27__lane15_strm0_cntl        = 'd0         ;
    std__pe27__lane15_strm0_data        = 'h1234_5678 ;
    std__pe27__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe27__lane15_strm1_cntl        = 'd0         ;
    std__pe27__lane15_strm1_data        = 'h1234_5678 ;
    std__pe27__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe27__lane16_strm0_cntl        = 'd0         ;
    std__pe27__lane16_strm0_data        = 'h1234_5678 ;
    std__pe27__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe27__lane16_strm1_cntl        = 'd0         ;
    std__pe27__lane16_strm1_data        = 'h1234_5678 ;
    std__pe27__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe27__lane17_strm0_cntl        = 'd0         ;
    std__pe27__lane17_strm0_data        = 'h1234_5678 ;
    std__pe27__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe27__lane17_strm1_cntl        = 'd0         ;
    std__pe27__lane17_strm1_data        = 'h1234_5678 ;
    std__pe27__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe27__lane18_strm0_cntl        = 'd0         ;
    std__pe27__lane18_strm0_data        = 'h1234_5678 ;
    std__pe27__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe27__lane18_strm1_cntl        = 'd0         ;
    std__pe27__lane18_strm1_data        = 'h1234_5678 ;
    std__pe27__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe27__lane19_strm0_cntl        = 'd0         ;
    std__pe27__lane19_strm0_data        = 'h1234_5678 ;
    std__pe27__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe27__lane19_strm1_cntl        = 'd0         ;
    std__pe27__lane19_strm1_data        = 'h1234_5678 ;
    std__pe27__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe27__lane20_strm0_cntl        = 'd0         ;
    std__pe27__lane20_strm0_data        = 'h1234_5678 ;
    std__pe27__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe27__lane20_strm1_cntl        = 'd0         ;
    std__pe27__lane20_strm1_data        = 'h1234_5678 ;
    std__pe27__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe27__lane21_strm0_cntl        = 'd0         ;
    std__pe27__lane21_strm0_data        = 'h1234_5678 ;
    std__pe27__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe27__lane21_strm1_cntl        = 'd0         ;
    std__pe27__lane21_strm1_data        = 'h1234_5678 ;
    std__pe27__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe27__lane22_strm0_cntl        = 'd0         ;
    std__pe27__lane22_strm0_data        = 'h1234_5678 ;
    std__pe27__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe27__lane22_strm1_cntl        = 'd0         ;
    std__pe27__lane22_strm1_data        = 'h1234_5678 ;
    std__pe27__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe27__lane23_strm0_cntl        = 'd0         ;
    std__pe27__lane23_strm0_data        = 'h1234_5678 ;
    std__pe27__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe27__lane23_strm1_cntl        = 'd0         ;
    std__pe27__lane23_strm1_data        = 'h1234_5678 ;
    std__pe27__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe27__lane24_strm0_cntl        = 'd0         ;
    std__pe27__lane24_strm0_data        = 'h1234_5678 ;
    std__pe27__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe27__lane24_strm1_cntl        = 'd0         ;
    std__pe27__lane24_strm1_data        = 'h1234_5678 ;
    std__pe27__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe27__lane25_strm0_cntl        = 'd0         ;
    std__pe27__lane25_strm0_data        = 'h1234_5678 ;
    std__pe27__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe27__lane25_strm1_cntl        = 'd0         ;
    std__pe27__lane25_strm1_data        = 'h1234_5678 ;
    std__pe27__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe27__lane26_strm0_cntl        = 'd0         ;
    std__pe27__lane26_strm0_data        = 'h1234_5678 ;
    std__pe27__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe27__lane26_strm1_cntl        = 'd0         ;
    std__pe27__lane26_strm1_data        = 'h1234_5678 ;
    std__pe27__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe27__lane27_strm0_cntl        = 'd0         ;
    std__pe27__lane27_strm0_data        = 'h1234_5678 ;
    std__pe27__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe27__lane27_strm1_cntl        = 'd0         ;
    std__pe27__lane27_strm1_data        = 'h1234_5678 ;
    std__pe27__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe27__lane28_strm0_cntl        = 'd0         ;
    std__pe27__lane28_strm0_data        = 'h1234_5678 ;
    std__pe27__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe27__lane28_strm1_cntl        = 'd0         ;
    std__pe27__lane28_strm1_data        = 'h1234_5678 ;
    std__pe27__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe27__lane29_strm0_cntl        = 'd0         ;
    std__pe27__lane29_strm0_data        = 'h1234_5678 ;
    std__pe27__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe27__lane29_strm1_cntl        = 'd0         ;
    std__pe27__lane29_strm1_data        = 'h1234_5678 ;
    std__pe27__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe27__lane30_strm0_cntl        = 'd0         ;
    std__pe27__lane30_strm0_data        = 'h1234_5678 ;
    std__pe27__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe27__lane30_strm1_cntl        = 'd0         ;
    std__pe27__lane30_strm1_data        = 'h1234_5678 ;
    std__pe27__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe27__lane31_strm0_cntl        = 'd0         ;
    std__pe27__lane31_strm0_data        = 'h1234_5678 ;
    std__pe27__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe27__lane31_strm1_cntl        = 'd0         ;
    std__pe27__lane31_strm1_data        = 'h1234_5678 ;
    std__pe27__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe28__lane0_strm0_cntl        = 'd0         ;
    std__pe28__lane0_strm0_data        = 'h1234_5678 ;
    std__pe28__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe28__lane0_strm1_cntl        = 'd0         ;
    std__pe28__lane0_strm1_data        = 'h1234_5678 ;
    std__pe28__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe28__lane1_strm0_cntl        = 'd0         ;
    std__pe28__lane1_strm0_data        = 'h1234_5678 ;
    std__pe28__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe28__lane1_strm1_cntl        = 'd0         ;
    std__pe28__lane1_strm1_data        = 'h1234_5678 ;
    std__pe28__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe28__lane2_strm0_cntl        = 'd0         ;
    std__pe28__lane2_strm0_data        = 'h1234_5678 ;
    std__pe28__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe28__lane2_strm1_cntl        = 'd0         ;
    std__pe28__lane2_strm1_data        = 'h1234_5678 ;
    std__pe28__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe28__lane3_strm0_cntl        = 'd0         ;
    std__pe28__lane3_strm0_data        = 'h1234_5678 ;
    std__pe28__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe28__lane3_strm1_cntl        = 'd0         ;
    std__pe28__lane3_strm1_data        = 'h1234_5678 ;
    std__pe28__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe28__lane4_strm0_cntl        = 'd0         ;
    std__pe28__lane4_strm0_data        = 'h1234_5678 ;
    std__pe28__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe28__lane4_strm1_cntl        = 'd0         ;
    std__pe28__lane4_strm1_data        = 'h1234_5678 ;
    std__pe28__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe28__lane5_strm0_cntl        = 'd0         ;
    std__pe28__lane5_strm0_data        = 'h1234_5678 ;
    std__pe28__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe28__lane5_strm1_cntl        = 'd0         ;
    std__pe28__lane5_strm1_data        = 'h1234_5678 ;
    std__pe28__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe28__lane6_strm0_cntl        = 'd0         ;
    std__pe28__lane6_strm0_data        = 'h1234_5678 ;
    std__pe28__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe28__lane6_strm1_cntl        = 'd0         ;
    std__pe28__lane6_strm1_data        = 'h1234_5678 ;
    std__pe28__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe28__lane7_strm0_cntl        = 'd0         ;
    std__pe28__lane7_strm0_data        = 'h1234_5678 ;
    std__pe28__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe28__lane7_strm1_cntl        = 'd0         ;
    std__pe28__lane7_strm1_data        = 'h1234_5678 ;
    std__pe28__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe28__lane8_strm0_cntl        = 'd0         ;
    std__pe28__lane8_strm0_data        = 'h1234_5678 ;
    std__pe28__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe28__lane8_strm1_cntl        = 'd0         ;
    std__pe28__lane8_strm1_data        = 'h1234_5678 ;
    std__pe28__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe28__lane9_strm0_cntl        = 'd0         ;
    std__pe28__lane9_strm0_data        = 'h1234_5678 ;
    std__pe28__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe28__lane9_strm1_cntl        = 'd0         ;
    std__pe28__lane9_strm1_data        = 'h1234_5678 ;
    std__pe28__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe28__lane10_strm0_cntl        = 'd0         ;
    std__pe28__lane10_strm0_data        = 'h1234_5678 ;
    std__pe28__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe28__lane10_strm1_cntl        = 'd0         ;
    std__pe28__lane10_strm1_data        = 'h1234_5678 ;
    std__pe28__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe28__lane11_strm0_cntl        = 'd0         ;
    std__pe28__lane11_strm0_data        = 'h1234_5678 ;
    std__pe28__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe28__lane11_strm1_cntl        = 'd0         ;
    std__pe28__lane11_strm1_data        = 'h1234_5678 ;
    std__pe28__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe28__lane12_strm0_cntl        = 'd0         ;
    std__pe28__lane12_strm0_data        = 'h1234_5678 ;
    std__pe28__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe28__lane12_strm1_cntl        = 'd0         ;
    std__pe28__lane12_strm1_data        = 'h1234_5678 ;
    std__pe28__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe28__lane13_strm0_cntl        = 'd0         ;
    std__pe28__lane13_strm0_data        = 'h1234_5678 ;
    std__pe28__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe28__lane13_strm1_cntl        = 'd0         ;
    std__pe28__lane13_strm1_data        = 'h1234_5678 ;
    std__pe28__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe28__lane14_strm0_cntl        = 'd0         ;
    std__pe28__lane14_strm0_data        = 'h1234_5678 ;
    std__pe28__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe28__lane14_strm1_cntl        = 'd0         ;
    std__pe28__lane14_strm1_data        = 'h1234_5678 ;
    std__pe28__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe28__lane15_strm0_cntl        = 'd0         ;
    std__pe28__lane15_strm0_data        = 'h1234_5678 ;
    std__pe28__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe28__lane15_strm1_cntl        = 'd0         ;
    std__pe28__lane15_strm1_data        = 'h1234_5678 ;
    std__pe28__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe28__lane16_strm0_cntl        = 'd0         ;
    std__pe28__lane16_strm0_data        = 'h1234_5678 ;
    std__pe28__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe28__lane16_strm1_cntl        = 'd0         ;
    std__pe28__lane16_strm1_data        = 'h1234_5678 ;
    std__pe28__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe28__lane17_strm0_cntl        = 'd0         ;
    std__pe28__lane17_strm0_data        = 'h1234_5678 ;
    std__pe28__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe28__lane17_strm1_cntl        = 'd0         ;
    std__pe28__lane17_strm1_data        = 'h1234_5678 ;
    std__pe28__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe28__lane18_strm0_cntl        = 'd0         ;
    std__pe28__lane18_strm0_data        = 'h1234_5678 ;
    std__pe28__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe28__lane18_strm1_cntl        = 'd0         ;
    std__pe28__lane18_strm1_data        = 'h1234_5678 ;
    std__pe28__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe28__lane19_strm0_cntl        = 'd0         ;
    std__pe28__lane19_strm0_data        = 'h1234_5678 ;
    std__pe28__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe28__lane19_strm1_cntl        = 'd0         ;
    std__pe28__lane19_strm1_data        = 'h1234_5678 ;
    std__pe28__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe28__lane20_strm0_cntl        = 'd0         ;
    std__pe28__lane20_strm0_data        = 'h1234_5678 ;
    std__pe28__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe28__lane20_strm1_cntl        = 'd0         ;
    std__pe28__lane20_strm1_data        = 'h1234_5678 ;
    std__pe28__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe28__lane21_strm0_cntl        = 'd0         ;
    std__pe28__lane21_strm0_data        = 'h1234_5678 ;
    std__pe28__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe28__lane21_strm1_cntl        = 'd0         ;
    std__pe28__lane21_strm1_data        = 'h1234_5678 ;
    std__pe28__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe28__lane22_strm0_cntl        = 'd0         ;
    std__pe28__lane22_strm0_data        = 'h1234_5678 ;
    std__pe28__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe28__lane22_strm1_cntl        = 'd0         ;
    std__pe28__lane22_strm1_data        = 'h1234_5678 ;
    std__pe28__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe28__lane23_strm0_cntl        = 'd0         ;
    std__pe28__lane23_strm0_data        = 'h1234_5678 ;
    std__pe28__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe28__lane23_strm1_cntl        = 'd0         ;
    std__pe28__lane23_strm1_data        = 'h1234_5678 ;
    std__pe28__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe28__lane24_strm0_cntl        = 'd0         ;
    std__pe28__lane24_strm0_data        = 'h1234_5678 ;
    std__pe28__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe28__lane24_strm1_cntl        = 'd0         ;
    std__pe28__lane24_strm1_data        = 'h1234_5678 ;
    std__pe28__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe28__lane25_strm0_cntl        = 'd0         ;
    std__pe28__lane25_strm0_data        = 'h1234_5678 ;
    std__pe28__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe28__lane25_strm1_cntl        = 'd0         ;
    std__pe28__lane25_strm1_data        = 'h1234_5678 ;
    std__pe28__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe28__lane26_strm0_cntl        = 'd0         ;
    std__pe28__lane26_strm0_data        = 'h1234_5678 ;
    std__pe28__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe28__lane26_strm1_cntl        = 'd0         ;
    std__pe28__lane26_strm1_data        = 'h1234_5678 ;
    std__pe28__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe28__lane27_strm0_cntl        = 'd0         ;
    std__pe28__lane27_strm0_data        = 'h1234_5678 ;
    std__pe28__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe28__lane27_strm1_cntl        = 'd0         ;
    std__pe28__lane27_strm1_data        = 'h1234_5678 ;
    std__pe28__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe28__lane28_strm0_cntl        = 'd0         ;
    std__pe28__lane28_strm0_data        = 'h1234_5678 ;
    std__pe28__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe28__lane28_strm1_cntl        = 'd0         ;
    std__pe28__lane28_strm1_data        = 'h1234_5678 ;
    std__pe28__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe28__lane29_strm0_cntl        = 'd0         ;
    std__pe28__lane29_strm0_data        = 'h1234_5678 ;
    std__pe28__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe28__lane29_strm1_cntl        = 'd0         ;
    std__pe28__lane29_strm1_data        = 'h1234_5678 ;
    std__pe28__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe28__lane30_strm0_cntl        = 'd0         ;
    std__pe28__lane30_strm0_data        = 'h1234_5678 ;
    std__pe28__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe28__lane30_strm1_cntl        = 'd0         ;
    std__pe28__lane30_strm1_data        = 'h1234_5678 ;
    std__pe28__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe28__lane31_strm0_cntl        = 'd0         ;
    std__pe28__lane31_strm0_data        = 'h1234_5678 ;
    std__pe28__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe28__lane31_strm1_cntl        = 'd0         ;
    std__pe28__lane31_strm1_data        = 'h1234_5678 ;
    std__pe28__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe29__lane0_strm0_cntl        = 'd0         ;
    std__pe29__lane0_strm0_data        = 'h1234_5678 ;
    std__pe29__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe29__lane0_strm1_cntl        = 'd0         ;
    std__pe29__lane0_strm1_data        = 'h1234_5678 ;
    std__pe29__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe29__lane1_strm0_cntl        = 'd0         ;
    std__pe29__lane1_strm0_data        = 'h1234_5678 ;
    std__pe29__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe29__lane1_strm1_cntl        = 'd0         ;
    std__pe29__lane1_strm1_data        = 'h1234_5678 ;
    std__pe29__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe29__lane2_strm0_cntl        = 'd0         ;
    std__pe29__lane2_strm0_data        = 'h1234_5678 ;
    std__pe29__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe29__lane2_strm1_cntl        = 'd0         ;
    std__pe29__lane2_strm1_data        = 'h1234_5678 ;
    std__pe29__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe29__lane3_strm0_cntl        = 'd0         ;
    std__pe29__lane3_strm0_data        = 'h1234_5678 ;
    std__pe29__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe29__lane3_strm1_cntl        = 'd0         ;
    std__pe29__lane3_strm1_data        = 'h1234_5678 ;
    std__pe29__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe29__lane4_strm0_cntl        = 'd0         ;
    std__pe29__lane4_strm0_data        = 'h1234_5678 ;
    std__pe29__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe29__lane4_strm1_cntl        = 'd0         ;
    std__pe29__lane4_strm1_data        = 'h1234_5678 ;
    std__pe29__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe29__lane5_strm0_cntl        = 'd0         ;
    std__pe29__lane5_strm0_data        = 'h1234_5678 ;
    std__pe29__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe29__lane5_strm1_cntl        = 'd0         ;
    std__pe29__lane5_strm1_data        = 'h1234_5678 ;
    std__pe29__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe29__lane6_strm0_cntl        = 'd0         ;
    std__pe29__lane6_strm0_data        = 'h1234_5678 ;
    std__pe29__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe29__lane6_strm1_cntl        = 'd0         ;
    std__pe29__lane6_strm1_data        = 'h1234_5678 ;
    std__pe29__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe29__lane7_strm0_cntl        = 'd0         ;
    std__pe29__lane7_strm0_data        = 'h1234_5678 ;
    std__pe29__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe29__lane7_strm1_cntl        = 'd0         ;
    std__pe29__lane7_strm1_data        = 'h1234_5678 ;
    std__pe29__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe29__lane8_strm0_cntl        = 'd0         ;
    std__pe29__lane8_strm0_data        = 'h1234_5678 ;
    std__pe29__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe29__lane8_strm1_cntl        = 'd0         ;
    std__pe29__lane8_strm1_data        = 'h1234_5678 ;
    std__pe29__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe29__lane9_strm0_cntl        = 'd0         ;
    std__pe29__lane9_strm0_data        = 'h1234_5678 ;
    std__pe29__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe29__lane9_strm1_cntl        = 'd0         ;
    std__pe29__lane9_strm1_data        = 'h1234_5678 ;
    std__pe29__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe29__lane10_strm0_cntl        = 'd0         ;
    std__pe29__lane10_strm0_data        = 'h1234_5678 ;
    std__pe29__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe29__lane10_strm1_cntl        = 'd0         ;
    std__pe29__lane10_strm1_data        = 'h1234_5678 ;
    std__pe29__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe29__lane11_strm0_cntl        = 'd0         ;
    std__pe29__lane11_strm0_data        = 'h1234_5678 ;
    std__pe29__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe29__lane11_strm1_cntl        = 'd0         ;
    std__pe29__lane11_strm1_data        = 'h1234_5678 ;
    std__pe29__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe29__lane12_strm0_cntl        = 'd0         ;
    std__pe29__lane12_strm0_data        = 'h1234_5678 ;
    std__pe29__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe29__lane12_strm1_cntl        = 'd0         ;
    std__pe29__lane12_strm1_data        = 'h1234_5678 ;
    std__pe29__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe29__lane13_strm0_cntl        = 'd0         ;
    std__pe29__lane13_strm0_data        = 'h1234_5678 ;
    std__pe29__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe29__lane13_strm1_cntl        = 'd0         ;
    std__pe29__lane13_strm1_data        = 'h1234_5678 ;
    std__pe29__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe29__lane14_strm0_cntl        = 'd0         ;
    std__pe29__lane14_strm0_data        = 'h1234_5678 ;
    std__pe29__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe29__lane14_strm1_cntl        = 'd0         ;
    std__pe29__lane14_strm1_data        = 'h1234_5678 ;
    std__pe29__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe29__lane15_strm0_cntl        = 'd0         ;
    std__pe29__lane15_strm0_data        = 'h1234_5678 ;
    std__pe29__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe29__lane15_strm1_cntl        = 'd0         ;
    std__pe29__lane15_strm1_data        = 'h1234_5678 ;
    std__pe29__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe29__lane16_strm0_cntl        = 'd0         ;
    std__pe29__lane16_strm0_data        = 'h1234_5678 ;
    std__pe29__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe29__lane16_strm1_cntl        = 'd0         ;
    std__pe29__lane16_strm1_data        = 'h1234_5678 ;
    std__pe29__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe29__lane17_strm0_cntl        = 'd0         ;
    std__pe29__lane17_strm0_data        = 'h1234_5678 ;
    std__pe29__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe29__lane17_strm1_cntl        = 'd0         ;
    std__pe29__lane17_strm1_data        = 'h1234_5678 ;
    std__pe29__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe29__lane18_strm0_cntl        = 'd0         ;
    std__pe29__lane18_strm0_data        = 'h1234_5678 ;
    std__pe29__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe29__lane18_strm1_cntl        = 'd0         ;
    std__pe29__lane18_strm1_data        = 'h1234_5678 ;
    std__pe29__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe29__lane19_strm0_cntl        = 'd0         ;
    std__pe29__lane19_strm0_data        = 'h1234_5678 ;
    std__pe29__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe29__lane19_strm1_cntl        = 'd0         ;
    std__pe29__lane19_strm1_data        = 'h1234_5678 ;
    std__pe29__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe29__lane20_strm0_cntl        = 'd0         ;
    std__pe29__lane20_strm0_data        = 'h1234_5678 ;
    std__pe29__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe29__lane20_strm1_cntl        = 'd0         ;
    std__pe29__lane20_strm1_data        = 'h1234_5678 ;
    std__pe29__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe29__lane21_strm0_cntl        = 'd0         ;
    std__pe29__lane21_strm0_data        = 'h1234_5678 ;
    std__pe29__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe29__lane21_strm1_cntl        = 'd0         ;
    std__pe29__lane21_strm1_data        = 'h1234_5678 ;
    std__pe29__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe29__lane22_strm0_cntl        = 'd0         ;
    std__pe29__lane22_strm0_data        = 'h1234_5678 ;
    std__pe29__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe29__lane22_strm1_cntl        = 'd0         ;
    std__pe29__lane22_strm1_data        = 'h1234_5678 ;
    std__pe29__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe29__lane23_strm0_cntl        = 'd0         ;
    std__pe29__lane23_strm0_data        = 'h1234_5678 ;
    std__pe29__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe29__lane23_strm1_cntl        = 'd0         ;
    std__pe29__lane23_strm1_data        = 'h1234_5678 ;
    std__pe29__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe29__lane24_strm0_cntl        = 'd0         ;
    std__pe29__lane24_strm0_data        = 'h1234_5678 ;
    std__pe29__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe29__lane24_strm1_cntl        = 'd0         ;
    std__pe29__lane24_strm1_data        = 'h1234_5678 ;
    std__pe29__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe29__lane25_strm0_cntl        = 'd0         ;
    std__pe29__lane25_strm0_data        = 'h1234_5678 ;
    std__pe29__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe29__lane25_strm1_cntl        = 'd0         ;
    std__pe29__lane25_strm1_data        = 'h1234_5678 ;
    std__pe29__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe29__lane26_strm0_cntl        = 'd0         ;
    std__pe29__lane26_strm0_data        = 'h1234_5678 ;
    std__pe29__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe29__lane26_strm1_cntl        = 'd0         ;
    std__pe29__lane26_strm1_data        = 'h1234_5678 ;
    std__pe29__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe29__lane27_strm0_cntl        = 'd0         ;
    std__pe29__lane27_strm0_data        = 'h1234_5678 ;
    std__pe29__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe29__lane27_strm1_cntl        = 'd0         ;
    std__pe29__lane27_strm1_data        = 'h1234_5678 ;
    std__pe29__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe29__lane28_strm0_cntl        = 'd0         ;
    std__pe29__lane28_strm0_data        = 'h1234_5678 ;
    std__pe29__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe29__lane28_strm1_cntl        = 'd0         ;
    std__pe29__lane28_strm1_data        = 'h1234_5678 ;
    std__pe29__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe29__lane29_strm0_cntl        = 'd0         ;
    std__pe29__lane29_strm0_data        = 'h1234_5678 ;
    std__pe29__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe29__lane29_strm1_cntl        = 'd0         ;
    std__pe29__lane29_strm1_data        = 'h1234_5678 ;
    std__pe29__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe29__lane30_strm0_cntl        = 'd0         ;
    std__pe29__lane30_strm0_data        = 'h1234_5678 ;
    std__pe29__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe29__lane30_strm1_cntl        = 'd0         ;
    std__pe29__lane30_strm1_data        = 'h1234_5678 ;
    std__pe29__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe29__lane31_strm0_cntl        = 'd0         ;
    std__pe29__lane31_strm0_data        = 'h1234_5678 ;
    std__pe29__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe29__lane31_strm1_cntl        = 'd0         ;
    std__pe29__lane31_strm1_data        = 'h1234_5678 ;
    std__pe29__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe30__lane0_strm0_cntl        = 'd0         ;
    std__pe30__lane0_strm0_data        = 'h1234_5678 ;
    std__pe30__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe30__lane0_strm1_cntl        = 'd0         ;
    std__pe30__lane0_strm1_data        = 'h1234_5678 ;
    std__pe30__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe30__lane1_strm0_cntl        = 'd0         ;
    std__pe30__lane1_strm0_data        = 'h1234_5678 ;
    std__pe30__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe30__lane1_strm1_cntl        = 'd0         ;
    std__pe30__lane1_strm1_data        = 'h1234_5678 ;
    std__pe30__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe30__lane2_strm0_cntl        = 'd0         ;
    std__pe30__lane2_strm0_data        = 'h1234_5678 ;
    std__pe30__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe30__lane2_strm1_cntl        = 'd0         ;
    std__pe30__lane2_strm1_data        = 'h1234_5678 ;
    std__pe30__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe30__lane3_strm0_cntl        = 'd0         ;
    std__pe30__lane3_strm0_data        = 'h1234_5678 ;
    std__pe30__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe30__lane3_strm1_cntl        = 'd0         ;
    std__pe30__lane3_strm1_data        = 'h1234_5678 ;
    std__pe30__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe30__lane4_strm0_cntl        = 'd0         ;
    std__pe30__lane4_strm0_data        = 'h1234_5678 ;
    std__pe30__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe30__lane4_strm1_cntl        = 'd0         ;
    std__pe30__lane4_strm1_data        = 'h1234_5678 ;
    std__pe30__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe30__lane5_strm0_cntl        = 'd0         ;
    std__pe30__lane5_strm0_data        = 'h1234_5678 ;
    std__pe30__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe30__lane5_strm1_cntl        = 'd0         ;
    std__pe30__lane5_strm1_data        = 'h1234_5678 ;
    std__pe30__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe30__lane6_strm0_cntl        = 'd0         ;
    std__pe30__lane6_strm0_data        = 'h1234_5678 ;
    std__pe30__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe30__lane6_strm1_cntl        = 'd0         ;
    std__pe30__lane6_strm1_data        = 'h1234_5678 ;
    std__pe30__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe30__lane7_strm0_cntl        = 'd0         ;
    std__pe30__lane7_strm0_data        = 'h1234_5678 ;
    std__pe30__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe30__lane7_strm1_cntl        = 'd0         ;
    std__pe30__lane7_strm1_data        = 'h1234_5678 ;
    std__pe30__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe30__lane8_strm0_cntl        = 'd0         ;
    std__pe30__lane8_strm0_data        = 'h1234_5678 ;
    std__pe30__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe30__lane8_strm1_cntl        = 'd0         ;
    std__pe30__lane8_strm1_data        = 'h1234_5678 ;
    std__pe30__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe30__lane9_strm0_cntl        = 'd0         ;
    std__pe30__lane9_strm0_data        = 'h1234_5678 ;
    std__pe30__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe30__lane9_strm1_cntl        = 'd0         ;
    std__pe30__lane9_strm1_data        = 'h1234_5678 ;
    std__pe30__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe30__lane10_strm0_cntl        = 'd0         ;
    std__pe30__lane10_strm0_data        = 'h1234_5678 ;
    std__pe30__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe30__lane10_strm1_cntl        = 'd0         ;
    std__pe30__lane10_strm1_data        = 'h1234_5678 ;
    std__pe30__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe30__lane11_strm0_cntl        = 'd0         ;
    std__pe30__lane11_strm0_data        = 'h1234_5678 ;
    std__pe30__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe30__lane11_strm1_cntl        = 'd0         ;
    std__pe30__lane11_strm1_data        = 'h1234_5678 ;
    std__pe30__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe30__lane12_strm0_cntl        = 'd0         ;
    std__pe30__lane12_strm0_data        = 'h1234_5678 ;
    std__pe30__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe30__lane12_strm1_cntl        = 'd0         ;
    std__pe30__lane12_strm1_data        = 'h1234_5678 ;
    std__pe30__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe30__lane13_strm0_cntl        = 'd0         ;
    std__pe30__lane13_strm0_data        = 'h1234_5678 ;
    std__pe30__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe30__lane13_strm1_cntl        = 'd0         ;
    std__pe30__lane13_strm1_data        = 'h1234_5678 ;
    std__pe30__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe30__lane14_strm0_cntl        = 'd0         ;
    std__pe30__lane14_strm0_data        = 'h1234_5678 ;
    std__pe30__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe30__lane14_strm1_cntl        = 'd0         ;
    std__pe30__lane14_strm1_data        = 'h1234_5678 ;
    std__pe30__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe30__lane15_strm0_cntl        = 'd0         ;
    std__pe30__lane15_strm0_data        = 'h1234_5678 ;
    std__pe30__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe30__lane15_strm1_cntl        = 'd0         ;
    std__pe30__lane15_strm1_data        = 'h1234_5678 ;
    std__pe30__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe30__lane16_strm0_cntl        = 'd0         ;
    std__pe30__lane16_strm0_data        = 'h1234_5678 ;
    std__pe30__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe30__lane16_strm1_cntl        = 'd0         ;
    std__pe30__lane16_strm1_data        = 'h1234_5678 ;
    std__pe30__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe30__lane17_strm0_cntl        = 'd0         ;
    std__pe30__lane17_strm0_data        = 'h1234_5678 ;
    std__pe30__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe30__lane17_strm1_cntl        = 'd0         ;
    std__pe30__lane17_strm1_data        = 'h1234_5678 ;
    std__pe30__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe30__lane18_strm0_cntl        = 'd0         ;
    std__pe30__lane18_strm0_data        = 'h1234_5678 ;
    std__pe30__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe30__lane18_strm1_cntl        = 'd0         ;
    std__pe30__lane18_strm1_data        = 'h1234_5678 ;
    std__pe30__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe30__lane19_strm0_cntl        = 'd0         ;
    std__pe30__lane19_strm0_data        = 'h1234_5678 ;
    std__pe30__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe30__lane19_strm1_cntl        = 'd0         ;
    std__pe30__lane19_strm1_data        = 'h1234_5678 ;
    std__pe30__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe30__lane20_strm0_cntl        = 'd0         ;
    std__pe30__lane20_strm0_data        = 'h1234_5678 ;
    std__pe30__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe30__lane20_strm1_cntl        = 'd0         ;
    std__pe30__lane20_strm1_data        = 'h1234_5678 ;
    std__pe30__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe30__lane21_strm0_cntl        = 'd0         ;
    std__pe30__lane21_strm0_data        = 'h1234_5678 ;
    std__pe30__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe30__lane21_strm1_cntl        = 'd0         ;
    std__pe30__lane21_strm1_data        = 'h1234_5678 ;
    std__pe30__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe30__lane22_strm0_cntl        = 'd0         ;
    std__pe30__lane22_strm0_data        = 'h1234_5678 ;
    std__pe30__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe30__lane22_strm1_cntl        = 'd0         ;
    std__pe30__lane22_strm1_data        = 'h1234_5678 ;
    std__pe30__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe30__lane23_strm0_cntl        = 'd0         ;
    std__pe30__lane23_strm0_data        = 'h1234_5678 ;
    std__pe30__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe30__lane23_strm1_cntl        = 'd0         ;
    std__pe30__lane23_strm1_data        = 'h1234_5678 ;
    std__pe30__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe30__lane24_strm0_cntl        = 'd0         ;
    std__pe30__lane24_strm0_data        = 'h1234_5678 ;
    std__pe30__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe30__lane24_strm1_cntl        = 'd0         ;
    std__pe30__lane24_strm1_data        = 'h1234_5678 ;
    std__pe30__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe30__lane25_strm0_cntl        = 'd0         ;
    std__pe30__lane25_strm0_data        = 'h1234_5678 ;
    std__pe30__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe30__lane25_strm1_cntl        = 'd0         ;
    std__pe30__lane25_strm1_data        = 'h1234_5678 ;
    std__pe30__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe30__lane26_strm0_cntl        = 'd0         ;
    std__pe30__lane26_strm0_data        = 'h1234_5678 ;
    std__pe30__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe30__lane26_strm1_cntl        = 'd0         ;
    std__pe30__lane26_strm1_data        = 'h1234_5678 ;
    std__pe30__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe30__lane27_strm0_cntl        = 'd0         ;
    std__pe30__lane27_strm0_data        = 'h1234_5678 ;
    std__pe30__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe30__lane27_strm1_cntl        = 'd0         ;
    std__pe30__lane27_strm1_data        = 'h1234_5678 ;
    std__pe30__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe30__lane28_strm0_cntl        = 'd0         ;
    std__pe30__lane28_strm0_data        = 'h1234_5678 ;
    std__pe30__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe30__lane28_strm1_cntl        = 'd0         ;
    std__pe30__lane28_strm1_data        = 'h1234_5678 ;
    std__pe30__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe30__lane29_strm0_cntl        = 'd0         ;
    std__pe30__lane29_strm0_data        = 'h1234_5678 ;
    std__pe30__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe30__lane29_strm1_cntl        = 'd0         ;
    std__pe30__lane29_strm1_data        = 'h1234_5678 ;
    std__pe30__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe30__lane30_strm0_cntl        = 'd0         ;
    std__pe30__lane30_strm0_data        = 'h1234_5678 ;
    std__pe30__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe30__lane30_strm1_cntl        = 'd0         ;
    std__pe30__lane30_strm1_data        = 'h1234_5678 ;
    std__pe30__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe30__lane31_strm0_cntl        = 'd0         ;
    std__pe30__lane31_strm0_data        = 'h1234_5678 ;
    std__pe30__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe30__lane31_strm1_cntl        = 'd0         ;
    std__pe30__lane31_strm1_data        = 'h1234_5678 ;
    std__pe30__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe31__lane0_strm0_cntl        = 'd0         ;
    std__pe31__lane0_strm0_data        = 'h1234_5678 ;
    std__pe31__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe31__lane0_strm1_cntl        = 'd0         ;
    std__pe31__lane0_strm1_data        = 'h1234_5678 ;
    std__pe31__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe31__lane1_strm0_cntl        = 'd0         ;
    std__pe31__lane1_strm0_data        = 'h1234_5678 ;
    std__pe31__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe31__lane1_strm1_cntl        = 'd0         ;
    std__pe31__lane1_strm1_data        = 'h1234_5678 ;
    std__pe31__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe31__lane2_strm0_cntl        = 'd0         ;
    std__pe31__lane2_strm0_data        = 'h1234_5678 ;
    std__pe31__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe31__lane2_strm1_cntl        = 'd0         ;
    std__pe31__lane2_strm1_data        = 'h1234_5678 ;
    std__pe31__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe31__lane3_strm0_cntl        = 'd0         ;
    std__pe31__lane3_strm0_data        = 'h1234_5678 ;
    std__pe31__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe31__lane3_strm1_cntl        = 'd0         ;
    std__pe31__lane3_strm1_data        = 'h1234_5678 ;
    std__pe31__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe31__lane4_strm0_cntl        = 'd0         ;
    std__pe31__lane4_strm0_data        = 'h1234_5678 ;
    std__pe31__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe31__lane4_strm1_cntl        = 'd0         ;
    std__pe31__lane4_strm1_data        = 'h1234_5678 ;
    std__pe31__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe31__lane5_strm0_cntl        = 'd0         ;
    std__pe31__lane5_strm0_data        = 'h1234_5678 ;
    std__pe31__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe31__lane5_strm1_cntl        = 'd0         ;
    std__pe31__lane5_strm1_data        = 'h1234_5678 ;
    std__pe31__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe31__lane6_strm0_cntl        = 'd0         ;
    std__pe31__lane6_strm0_data        = 'h1234_5678 ;
    std__pe31__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe31__lane6_strm1_cntl        = 'd0         ;
    std__pe31__lane6_strm1_data        = 'h1234_5678 ;
    std__pe31__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe31__lane7_strm0_cntl        = 'd0         ;
    std__pe31__lane7_strm0_data        = 'h1234_5678 ;
    std__pe31__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe31__lane7_strm1_cntl        = 'd0         ;
    std__pe31__lane7_strm1_data        = 'h1234_5678 ;
    std__pe31__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe31__lane8_strm0_cntl        = 'd0         ;
    std__pe31__lane8_strm0_data        = 'h1234_5678 ;
    std__pe31__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe31__lane8_strm1_cntl        = 'd0         ;
    std__pe31__lane8_strm1_data        = 'h1234_5678 ;
    std__pe31__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe31__lane9_strm0_cntl        = 'd0         ;
    std__pe31__lane9_strm0_data        = 'h1234_5678 ;
    std__pe31__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe31__lane9_strm1_cntl        = 'd0         ;
    std__pe31__lane9_strm1_data        = 'h1234_5678 ;
    std__pe31__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe31__lane10_strm0_cntl        = 'd0         ;
    std__pe31__lane10_strm0_data        = 'h1234_5678 ;
    std__pe31__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe31__lane10_strm1_cntl        = 'd0         ;
    std__pe31__lane10_strm1_data        = 'h1234_5678 ;
    std__pe31__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe31__lane11_strm0_cntl        = 'd0         ;
    std__pe31__lane11_strm0_data        = 'h1234_5678 ;
    std__pe31__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe31__lane11_strm1_cntl        = 'd0         ;
    std__pe31__lane11_strm1_data        = 'h1234_5678 ;
    std__pe31__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe31__lane12_strm0_cntl        = 'd0         ;
    std__pe31__lane12_strm0_data        = 'h1234_5678 ;
    std__pe31__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe31__lane12_strm1_cntl        = 'd0         ;
    std__pe31__lane12_strm1_data        = 'h1234_5678 ;
    std__pe31__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe31__lane13_strm0_cntl        = 'd0         ;
    std__pe31__lane13_strm0_data        = 'h1234_5678 ;
    std__pe31__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe31__lane13_strm1_cntl        = 'd0         ;
    std__pe31__lane13_strm1_data        = 'h1234_5678 ;
    std__pe31__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe31__lane14_strm0_cntl        = 'd0         ;
    std__pe31__lane14_strm0_data        = 'h1234_5678 ;
    std__pe31__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe31__lane14_strm1_cntl        = 'd0         ;
    std__pe31__lane14_strm1_data        = 'h1234_5678 ;
    std__pe31__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe31__lane15_strm0_cntl        = 'd0         ;
    std__pe31__lane15_strm0_data        = 'h1234_5678 ;
    std__pe31__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe31__lane15_strm1_cntl        = 'd0         ;
    std__pe31__lane15_strm1_data        = 'h1234_5678 ;
    std__pe31__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe31__lane16_strm0_cntl        = 'd0         ;
    std__pe31__lane16_strm0_data        = 'h1234_5678 ;
    std__pe31__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe31__lane16_strm1_cntl        = 'd0         ;
    std__pe31__lane16_strm1_data        = 'h1234_5678 ;
    std__pe31__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe31__lane17_strm0_cntl        = 'd0         ;
    std__pe31__lane17_strm0_data        = 'h1234_5678 ;
    std__pe31__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe31__lane17_strm1_cntl        = 'd0         ;
    std__pe31__lane17_strm1_data        = 'h1234_5678 ;
    std__pe31__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe31__lane18_strm0_cntl        = 'd0         ;
    std__pe31__lane18_strm0_data        = 'h1234_5678 ;
    std__pe31__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe31__lane18_strm1_cntl        = 'd0         ;
    std__pe31__lane18_strm1_data        = 'h1234_5678 ;
    std__pe31__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe31__lane19_strm0_cntl        = 'd0         ;
    std__pe31__lane19_strm0_data        = 'h1234_5678 ;
    std__pe31__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe31__lane19_strm1_cntl        = 'd0         ;
    std__pe31__lane19_strm1_data        = 'h1234_5678 ;
    std__pe31__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe31__lane20_strm0_cntl        = 'd0         ;
    std__pe31__lane20_strm0_data        = 'h1234_5678 ;
    std__pe31__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe31__lane20_strm1_cntl        = 'd0         ;
    std__pe31__lane20_strm1_data        = 'h1234_5678 ;
    std__pe31__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe31__lane21_strm0_cntl        = 'd0         ;
    std__pe31__lane21_strm0_data        = 'h1234_5678 ;
    std__pe31__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe31__lane21_strm1_cntl        = 'd0         ;
    std__pe31__lane21_strm1_data        = 'h1234_5678 ;
    std__pe31__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe31__lane22_strm0_cntl        = 'd0         ;
    std__pe31__lane22_strm0_data        = 'h1234_5678 ;
    std__pe31__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe31__lane22_strm1_cntl        = 'd0         ;
    std__pe31__lane22_strm1_data        = 'h1234_5678 ;
    std__pe31__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe31__lane23_strm0_cntl        = 'd0         ;
    std__pe31__lane23_strm0_data        = 'h1234_5678 ;
    std__pe31__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe31__lane23_strm1_cntl        = 'd0         ;
    std__pe31__lane23_strm1_data        = 'h1234_5678 ;
    std__pe31__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe31__lane24_strm0_cntl        = 'd0         ;
    std__pe31__lane24_strm0_data        = 'h1234_5678 ;
    std__pe31__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe31__lane24_strm1_cntl        = 'd0         ;
    std__pe31__lane24_strm1_data        = 'h1234_5678 ;
    std__pe31__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe31__lane25_strm0_cntl        = 'd0         ;
    std__pe31__lane25_strm0_data        = 'h1234_5678 ;
    std__pe31__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe31__lane25_strm1_cntl        = 'd0         ;
    std__pe31__lane25_strm1_data        = 'h1234_5678 ;
    std__pe31__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe31__lane26_strm0_cntl        = 'd0         ;
    std__pe31__lane26_strm0_data        = 'h1234_5678 ;
    std__pe31__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe31__lane26_strm1_cntl        = 'd0         ;
    std__pe31__lane26_strm1_data        = 'h1234_5678 ;
    std__pe31__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe31__lane27_strm0_cntl        = 'd0         ;
    std__pe31__lane27_strm0_data        = 'h1234_5678 ;
    std__pe31__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe31__lane27_strm1_cntl        = 'd0         ;
    std__pe31__lane27_strm1_data        = 'h1234_5678 ;
    std__pe31__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe31__lane28_strm0_cntl        = 'd0         ;
    std__pe31__lane28_strm0_data        = 'h1234_5678 ;
    std__pe31__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe31__lane28_strm1_cntl        = 'd0         ;
    std__pe31__lane28_strm1_data        = 'h1234_5678 ;
    std__pe31__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe31__lane29_strm0_cntl        = 'd0         ;
    std__pe31__lane29_strm0_data        = 'h1234_5678 ;
    std__pe31__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe31__lane29_strm1_cntl        = 'd0         ;
    std__pe31__lane29_strm1_data        = 'h1234_5678 ;
    std__pe31__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe31__lane30_strm0_cntl        = 'd0         ;
    std__pe31__lane30_strm0_data        = 'h1234_5678 ;
    std__pe31__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe31__lane30_strm1_cntl        = 'd0         ;
    std__pe31__lane30_strm1_data        = 'h1234_5678 ;
    std__pe31__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe31__lane31_strm0_cntl        = 'd0         ;
    std__pe31__lane31_strm0_data        = 'h1234_5678 ;
    std__pe31__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe31__lane31_strm1_cntl        = 'd0         ;
    std__pe31__lane31_strm1_data        = 'h1234_5678 ;
    std__pe31__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe32__lane0_strm0_cntl        = 'd0         ;
    std__pe32__lane0_strm0_data        = 'h1234_5678 ;
    std__pe32__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe32__lane0_strm1_cntl        = 'd0         ;
    std__pe32__lane0_strm1_data        = 'h1234_5678 ;
    std__pe32__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe32__lane1_strm0_cntl        = 'd0         ;
    std__pe32__lane1_strm0_data        = 'h1234_5678 ;
    std__pe32__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe32__lane1_strm1_cntl        = 'd0         ;
    std__pe32__lane1_strm1_data        = 'h1234_5678 ;
    std__pe32__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe32__lane2_strm0_cntl        = 'd0         ;
    std__pe32__lane2_strm0_data        = 'h1234_5678 ;
    std__pe32__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe32__lane2_strm1_cntl        = 'd0         ;
    std__pe32__lane2_strm1_data        = 'h1234_5678 ;
    std__pe32__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe32__lane3_strm0_cntl        = 'd0         ;
    std__pe32__lane3_strm0_data        = 'h1234_5678 ;
    std__pe32__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe32__lane3_strm1_cntl        = 'd0         ;
    std__pe32__lane3_strm1_data        = 'h1234_5678 ;
    std__pe32__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe32__lane4_strm0_cntl        = 'd0         ;
    std__pe32__lane4_strm0_data        = 'h1234_5678 ;
    std__pe32__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe32__lane4_strm1_cntl        = 'd0         ;
    std__pe32__lane4_strm1_data        = 'h1234_5678 ;
    std__pe32__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe32__lane5_strm0_cntl        = 'd0         ;
    std__pe32__lane5_strm0_data        = 'h1234_5678 ;
    std__pe32__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe32__lane5_strm1_cntl        = 'd0         ;
    std__pe32__lane5_strm1_data        = 'h1234_5678 ;
    std__pe32__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe32__lane6_strm0_cntl        = 'd0         ;
    std__pe32__lane6_strm0_data        = 'h1234_5678 ;
    std__pe32__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe32__lane6_strm1_cntl        = 'd0         ;
    std__pe32__lane6_strm1_data        = 'h1234_5678 ;
    std__pe32__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe32__lane7_strm0_cntl        = 'd0         ;
    std__pe32__lane7_strm0_data        = 'h1234_5678 ;
    std__pe32__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe32__lane7_strm1_cntl        = 'd0         ;
    std__pe32__lane7_strm1_data        = 'h1234_5678 ;
    std__pe32__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe32__lane8_strm0_cntl        = 'd0         ;
    std__pe32__lane8_strm0_data        = 'h1234_5678 ;
    std__pe32__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe32__lane8_strm1_cntl        = 'd0         ;
    std__pe32__lane8_strm1_data        = 'h1234_5678 ;
    std__pe32__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe32__lane9_strm0_cntl        = 'd0         ;
    std__pe32__lane9_strm0_data        = 'h1234_5678 ;
    std__pe32__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe32__lane9_strm1_cntl        = 'd0         ;
    std__pe32__lane9_strm1_data        = 'h1234_5678 ;
    std__pe32__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe32__lane10_strm0_cntl        = 'd0         ;
    std__pe32__lane10_strm0_data        = 'h1234_5678 ;
    std__pe32__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe32__lane10_strm1_cntl        = 'd0         ;
    std__pe32__lane10_strm1_data        = 'h1234_5678 ;
    std__pe32__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe32__lane11_strm0_cntl        = 'd0         ;
    std__pe32__lane11_strm0_data        = 'h1234_5678 ;
    std__pe32__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe32__lane11_strm1_cntl        = 'd0         ;
    std__pe32__lane11_strm1_data        = 'h1234_5678 ;
    std__pe32__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe32__lane12_strm0_cntl        = 'd0         ;
    std__pe32__lane12_strm0_data        = 'h1234_5678 ;
    std__pe32__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe32__lane12_strm1_cntl        = 'd0         ;
    std__pe32__lane12_strm1_data        = 'h1234_5678 ;
    std__pe32__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe32__lane13_strm0_cntl        = 'd0         ;
    std__pe32__lane13_strm0_data        = 'h1234_5678 ;
    std__pe32__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe32__lane13_strm1_cntl        = 'd0         ;
    std__pe32__lane13_strm1_data        = 'h1234_5678 ;
    std__pe32__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe32__lane14_strm0_cntl        = 'd0         ;
    std__pe32__lane14_strm0_data        = 'h1234_5678 ;
    std__pe32__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe32__lane14_strm1_cntl        = 'd0         ;
    std__pe32__lane14_strm1_data        = 'h1234_5678 ;
    std__pe32__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe32__lane15_strm0_cntl        = 'd0         ;
    std__pe32__lane15_strm0_data        = 'h1234_5678 ;
    std__pe32__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe32__lane15_strm1_cntl        = 'd0         ;
    std__pe32__lane15_strm1_data        = 'h1234_5678 ;
    std__pe32__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe32__lane16_strm0_cntl        = 'd0         ;
    std__pe32__lane16_strm0_data        = 'h1234_5678 ;
    std__pe32__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe32__lane16_strm1_cntl        = 'd0         ;
    std__pe32__lane16_strm1_data        = 'h1234_5678 ;
    std__pe32__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe32__lane17_strm0_cntl        = 'd0         ;
    std__pe32__lane17_strm0_data        = 'h1234_5678 ;
    std__pe32__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe32__lane17_strm1_cntl        = 'd0         ;
    std__pe32__lane17_strm1_data        = 'h1234_5678 ;
    std__pe32__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe32__lane18_strm0_cntl        = 'd0         ;
    std__pe32__lane18_strm0_data        = 'h1234_5678 ;
    std__pe32__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe32__lane18_strm1_cntl        = 'd0         ;
    std__pe32__lane18_strm1_data        = 'h1234_5678 ;
    std__pe32__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe32__lane19_strm0_cntl        = 'd0         ;
    std__pe32__lane19_strm0_data        = 'h1234_5678 ;
    std__pe32__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe32__lane19_strm1_cntl        = 'd0         ;
    std__pe32__lane19_strm1_data        = 'h1234_5678 ;
    std__pe32__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe32__lane20_strm0_cntl        = 'd0         ;
    std__pe32__lane20_strm0_data        = 'h1234_5678 ;
    std__pe32__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe32__lane20_strm1_cntl        = 'd0         ;
    std__pe32__lane20_strm1_data        = 'h1234_5678 ;
    std__pe32__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe32__lane21_strm0_cntl        = 'd0         ;
    std__pe32__lane21_strm0_data        = 'h1234_5678 ;
    std__pe32__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe32__lane21_strm1_cntl        = 'd0         ;
    std__pe32__lane21_strm1_data        = 'h1234_5678 ;
    std__pe32__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe32__lane22_strm0_cntl        = 'd0         ;
    std__pe32__lane22_strm0_data        = 'h1234_5678 ;
    std__pe32__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe32__lane22_strm1_cntl        = 'd0         ;
    std__pe32__lane22_strm1_data        = 'h1234_5678 ;
    std__pe32__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe32__lane23_strm0_cntl        = 'd0         ;
    std__pe32__lane23_strm0_data        = 'h1234_5678 ;
    std__pe32__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe32__lane23_strm1_cntl        = 'd0         ;
    std__pe32__lane23_strm1_data        = 'h1234_5678 ;
    std__pe32__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe32__lane24_strm0_cntl        = 'd0         ;
    std__pe32__lane24_strm0_data        = 'h1234_5678 ;
    std__pe32__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe32__lane24_strm1_cntl        = 'd0         ;
    std__pe32__lane24_strm1_data        = 'h1234_5678 ;
    std__pe32__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe32__lane25_strm0_cntl        = 'd0         ;
    std__pe32__lane25_strm0_data        = 'h1234_5678 ;
    std__pe32__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe32__lane25_strm1_cntl        = 'd0         ;
    std__pe32__lane25_strm1_data        = 'h1234_5678 ;
    std__pe32__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe32__lane26_strm0_cntl        = 'd0         ;
    std__pe32__lane26_strm0_data        = 'h1234_5678 ;
    std__pe32__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe32__lane26_strm1_cntl        = 'd0         ;
    std__pe32__lane26_strm1_data        = 'h1234_5678 ;
    std__pe32__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe32__lane27_strm0_cntl        = 'd0         ;
    std__pe32__lane27_strm0_data        = 'h1234_5678 ;
    std__pe32__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe32__lane27_strm1_cntl        = 'd0         ;
    std__pe32__lane27_strm1_data        = 'h1234_5678 ;
    std__pe32__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe32__lane28_strm0_cntl        = 'd0         ;
    std__pe32__lane28_strm0_data        = 'h1234_5678 ;
    std__pe32__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe32__lane28_strm1_cntl        = 'd0         ;
    std__pe32__lane28_strm1_data        = 'h1234_5678 ;
    std__pe32__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe32__lane29_strm0_cntl        = 'd0         ;
    std__pe32__lane29_strm0_data        = 'h1234_5678 ;
    std__pe32__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe32__lane29_strm1_cntl        = 'd0         ;
    std__pe32__lane29_strm1_data        = 'h1234_5678 ;
    std__pe32__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe32__lane30_strm0_cntl        = 'd0         ;
    std__pe32__lane30_strm0_data        = 'h1234_5678 ;
    std__pe32__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe32__lane30_strm1_cntl        = 'd0         ;
    std__pe32__lane30_strm1_data        = 'h1234_5678 ;
    std__pe32__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe32__lane31_strm0_cntl        = 'd0         ;
    std__pe32__lane31_strm0_data        = 'h1234_5678 ;
    std__pe32__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe32__lane31_strm1_cntl        = 'd0         ;
    std__pe32__lane31_strm1_data        = 'h1234_5678 ;
    std__pe32__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe33__lane0_strm0_cntl        = 'd0         ;
    std__pe33__lane0_strm0_data        = 'h1234_5678 ;
    std__pe33__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe33__lane0_strm1_cntl        = 'd0         ;
    std__pe33__lane0_strm1_data        = 'h1234_5678 ;
    std__pe33__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe33__lane1_strm0_cntl        = 'd0         ;
    std__pe33__lane1_strm0_data        = 'h1234_5678 ;
    std__pe33__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe33__lane1_strm1_cntl        = 'd0         ;
    std__pe33__lane1_strm1_data        = 'h1234_5678 ;
    std__pe33__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe33__lane2_strm0_cntl        = 'd0         ;
    std__pe33__lane2_strm0_data        = 'h1234_5678 ;
    std__pe33__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe33__lane2_strm1_cntl        = 'd0         ;
    std__pe33__lane2_strm1_data        = 'h1234_5678 ;
    std__pe33__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe33__lane3_strm0_cntl        = 'd0         ;
    std__pe33__lane3_strm0_data        = 'h1234_5678 ;
    std__pe33__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe33__lane3_strm1_cntl        = 'd0         ;
    std__pe33__lane3_strm1_data        = 'h1234_5678 ;
    std__pe33__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe33__lane4_strm0_cntl        = 'd0         ;
    std__pe33__lane4_strm0_data        = 'h1234_5678 ;
    std__pe33__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe33__lane4_strm1_cntl        = 'd0         ;
    std__pe33__lane4_strm1_data        = 'h1234_5678 ;
    std__pe33__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe33__lane5_strm0_cntl        = 'd0         ;
    std__pe33__lane5_strm0_data        = 'h1234_5678 ;
    std__pe33__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe33__lane5_strm1_cntl        = 'd0         ;
    std__pe33__lane5_strm1_data        = 'h1234_5678 ;
    std__pe33__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe33__lane6_strm0_cntl        = 'd0         ;
    std__pe33__lane6_strm0_data        = 'h1234_5678 ;
    std__pe33__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe33__lane6_strm1_cntl        = 'd0         ;
    std__pe33__lane6_strm1_data        = 'h1234_5678 ;
    std__pe33__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe33__lane7_strm0_cntl        = 'd0         ;
    std__pe33__lane7_strm0_data        = 'h1234_5678 ;
    std__pe33__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe33__lane7_strm1_cntl        = 'd0         ;
    std__pe33__lane7_strm1_data        = 'h1234_5678 ;
    std__pe33__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe33__lane8_strm0_cntl        = 'd0         ;
    std__pe33__lane8_strm0_data        = 'h1234_5678 ;
    std__pe33__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe33__lane8_strm1_cntl        = 'd0         ;
    std__pe33__lane8_strm1_data        = 'h1234_5678 ;
    std__pe33__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe33__lane9_strm0_cntl        = 'd0         ;
    std__pe33__lane9_strm0_data        = 'h1234_5678 ;
    std__pe33__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe33__lane9_strm1_cntl        = 'd0         ;
    std__pe33__lane9_strm1_data        = 'h1234_5678 ;
    std__pe33__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe33__lane10_strm0_cntl        = 'd0         ;
    std__pe33__lane10_strm0_data        = 'h1234_5678 ;
    std__pe33__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe33__lane10_strm1_cntl        = 'd0         ;
    std__pe33__lane10_strm1_data        = 'h1234_5678 ;
    std__pe33__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe33__lane11_strm0_cntl        = 'd0         ;
    std__pe33__lane11_strm0_data        = 'h1234_5678 ;
    std__pe33__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe33__lane11_strm1_cntl        = 'd0         ;
    std__pe33__lane11_strm1_data        = 'h1234_5678 ;
    std__pe33__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe33__lane12_strm0_cntl        = 'd0         ;
    std__pe33__lane12_strm0_data        = 'h1234_5678 ;
    std__pe33__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe33__lane12_strm1_cntl        = 'd0         ;
    std__pe33__lane12_strm1_data        = 'h1234_5678 ;
    std__pe33__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe33__lane13_strm0_cntl        = 'd0         ;
    std__pe33__lane13_strm0_data        = 'h1234_5678 ;
    std__pe33__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe33__lane13_strm1_cntl        = 'd0         ;
    std__pe33__lane13_strm1_data        = 'h1234_5678 ;
    std__pe33__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe33__lane14_strm0_cntl        = 'd0         ;
    std__pe33__lane14_strm0_data        = 'h1234_5678 ;
    std__pe33__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe33__lane14_strm1_cntl        = 'd0         ;
    std__pe33__lane14_strm1_data        = 'h1234_5678 ;
    std__pe33__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe33__lane15_strm0_cntl        = 'd0         ;
    std__pe33__lane15_strm0_data        = 'h1234_5678 ;
    std__pe33__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe33__lane15_strm1_cntl        = 'd0         ;
    std__pe33__lane15_strm1_data        = 'h1234_5678 ;
    std__pe33__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe33__lane16_strm0_cntl        = 'd0         ;
    std__pe33__lane16_strm0_data        = 'h1234_5678 ;
    std__pe33__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe33__lane16_strm1_cntl        = 'd0         ;
    std__pe33__lane16_strm1_data        = 'h1234_5678 ;
    std__pe33__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe33__lane17_strm0_cntl        = 'd0         ;
    std__pe33__lane17_strm0_data        = 'h1234_5678 ;
    std__pe33__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe33__lane17_strm1_cntl        = 'd0         ;
    std__pe33__lane17_strm1_data        = 'h1234_5678 ;
    std__pe33__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe33__lane18_strm0_cntl        = 'd0         ;
    std__pe33__lane18_strm0_data        = 'h1234_5678 ;
    std__pe33__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe33__lane18_strm1_cntl        = 'd0         ;
    std__pe33__lane18_strm1_data        = 'h1234_5678 ;
    std__pe33__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe33__lane19_strm0_cntl        = 'd0         ;
    std__pe33__lane19_strm0_data        = 'h1234_5678 ;
    std__pe33__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe33__lane19_strm1_cntl        = 'd0         ;
    std__pe33__lane19_strm1_data        = 'h1234_5678 ;
    std__pe33__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe33__lane20_strm0_cntl        = 'd0         ;
    std__pe33__lane20_strm0_data        = 'h1234_5678 ;
    std__pe33__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe33__lane20_strm1_cntl        = 'd0         ;
    std__pe33__lane20_strm1_data        = 'h1234_5678 ;
    std__pe33__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe33__lane21_strm0_cntl        = 'd0         ;
    std__pe33__lane21_strm0_data        = 'h1234_5678 ;
    std__pe33__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe33__lane21_strm1_cntl        = 'd0         ;
    std__pe33__lane21_strm1_data        = 'h1234_5678 ;
    std__pe33__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe33__lane22_strm0_cntl        = 'd0         ;
    std__pe33__lane22_strm0_data        = 'h1234_5678 ;
    std__pe33__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe33__lane22_strm1_cntl        = 'd0         ;
    std__pe33__lane22_strm1_data        = 'h1234_5678 ;
    std__pe33__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe33__lane23_strm0_cntl        = 'd0         ;
    std__pe33__lane23_strm0_data        = 'h1234_5678 ;
    std__pe33__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe33__lane23_strm1_cntl        = 'd0         ;
    std__pe33__lane23_strm1_data        = 'h1234_5678 ;
    std__pe33__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe33__lane24_strm0_cntl        = 'd0         ;
    std__pe33__lane24_strm0_data        = 'h1234_5678 ;
    std__pe33__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe33__lane24_strm1_cntl        = 'd0         ;
    std__pe33__lane24_strm1_data        = 'h1234_5678 ;
    std__pe33__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe33__lane25_strm0_cntl        = 'd0         ;
    std__pe33__lane25_strm0_data        = 'h1234_5678 ;
    std__pe33__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe33__lane25_strm1_cntl        = 'd0         ;
    std__pe33__lane25_strm1_data        = 'h1234_5678 ;
    std__pe33__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe33__lane26_strm0_cntl        = 'd0         ;
    std__pe33__lane26_strm0_data        = 'h1234_5678 ;
    std__pe33__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe33__lane26_strm1_cntl        = 'd0         ;
    std__pe33__lane26_strm1_data        = 'h1234_5678 ;
    std__pe33__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe33__lane27_strm0_cntl        = 'd0         ;
    std__pe33__lane27_strm0_data        = 'h1234_5678 ;
    std__pe33__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe33__lane27_strm1_cntl        = 'd0         ;
    std__pe33__lane27_strm1_data        = 'h1234_5678 ;
    std__pe33__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe33__lane28_strm0_cntl        = 'd0         ;
    std__pe33__lane28_strm0_data        = 'h1234_5678 ;
    std__pe33__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe33__lane28_strm1_cntl        = 'd0         ;
    std__pe33__lane28_strm1_data        = 'h1234_5678 ;
    std__pe33__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe33__lane29_strm0_cntl        = 'd0         ;
    std__pe33__lane29_strm0_data        = 'h1234_5678 ;
    std__pe33__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe33__lane29_strm1_cntl        = 'd0         ;
    std__pe33__lane29_strm1_data        = 'h1234_5678 ;
    std__pe33__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe33__lane30_strm0_cntl        = 'd0         ;
    std__pe33__lane30_strm0_data        = 'h1234_5678 ;
    std__pe33__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe33__lane30_strm1_cntl        = 'd0         ;
    std__pe33__lane30_strm1_data        = 'h1234_5678 ;
    std__pe33__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe33__lane31_strm0_cntl        = 'd0         ;
    std__pe33__lane31_strm0_data        = 'h1234_5678 ;
    std__pe33__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe33__lane31_strm1_cntl        = 'd0         ;
    std__pe33__lane31_strm1_data        = 'h1234_5678 ;
    std__pe33__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe34__lane0_strm0_cntl        = 'd0         ;
    std__pe34__lane0_strm0_data        = 'h1234_5678 ;
    std__pe34__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe34__lane0_strm1_cntl        = 'd0         ;
    std__pe34__lane0_strm1_data        = 'h1234_5678 ;
    std__pe34__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe34__lane1_strm0_cntl        = 'd0         ;
    std__pe34__lane1_strm0_data        = 'h1234_5678 ;
    std__pe34__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe34__lane1_strm1_cntl        = 'd0         ;
    std__pe34__lane1_strm1_data        = 'h1234_5678 ;
    std__pe34__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe34__lane2_strm0_cntl        = 'd0         ;
    std__pe34__lane2_strm0_data        = 'h1234_5678 ;
    std__pe34__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe34__lane2_strm1_cntl        = 'd0         ;
    std__pe34__lane2_strm1_data        = 'h1234_5678 ;
    std__pe34__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe34__lane3_strm0_cntl        = 'd0         ;
    std__pe34__lane3_strm0_data        = 'h1234_5678 ;
    std__pe34__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe34__lane3_strm1_cntl        = 'd0         ;
    std__pe34__lane3_strm1_data        = 'h1234_5678 ;
    std__pe34__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe34__lane4_strm0_cntl        = 'd0         ;
    std__pe34__lane4_strm0_data        = 'h1234_5678 ;
    std__pe34__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe34__lane4_strm1_cntl        = 'd0         ;
    std__pe34__lane4_strm1_data        = 'h1234_5678 ;
    std__pe34__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe34__lane5_strm0_cntl        = 'd0         ;
    std__pe34__lane5_strm0_data        = 'h1234_5678 ;
    std__pe34__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe34__lane5_strm1_cntl        = 'd0         ;
    std__pe34__lane5_strm1_data        = 'h1234_5678 ;
    std__pe34__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe34__lane6_strm0_cntl        = 'd0         ;
    std__pe34__lane6_strm0_data        = 'h1234_5678 ;
    std__pe34__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe34__lane6_strm1_cntl        = 'd0         ;
    std__pe34__lane6_strm1_data        = 'h1234_5678 ;
    std__pe34__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe34__lane7_strm0_cntl        = 'd0         ;
    std__pe34__lane7_strm0_data        = 'h1234_5678 ;
    std__pe34__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe34__lane7_strm1_cntl        = 'd0         ;
    std__pe34__lane7_strm1_data        = 'h1234_5678 ;
    std__pe34__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe34__lane8_strm0_cntl        = 'd0         ;
    std__pe34__lane8_strm0_data        = 'h1234_5678 ;
    std__pe34__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe34__lane8_strm1_cntl        = 'd0         ;
    std__pe34__lane8_strm1_data        = 'h1234_5678 ;
    std__pe34__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe34__lane9_strm0_cntl        = 'd0         ;
    std__pe34__lane9_strm0_data        = 'h1234_5678 ;
    std__pe34__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe34__lane9_strm1_cntl        = 'd0         ;
    std__pe34__lane9_strm1_data        = 'h1234_5678 ;
    std__pe34__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe34__lane10_strm0_cntl        = 'd0         ;
    std__pe34__lane10_strm0_data        = 'h1234_5678 ;
    std__pe34__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe34__lane10_strm1_cntl        = 'd0         ;
    std__pe34__lane10_strm1_data        = 'h1234_5678 ;
    std__pe34__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe34__lane11_strm0_cntl        = 'd0         ;
    std__pe34__lane11_strm0_data        = 'h1234_5678 ;
    std__pe34__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe34__lane11_strm1_cntl        = 'd0         ;
    std__pe34__lane11_strm1_data        = 'h1234_5678 ;
    std__pe34__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe34__lane12_strm0_cntl        = 'd0         ;
    std__pe34__lane12_strm0_data        = 'h1234_5678 ;
    std__pe34__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe34__lane12_strm1_cntl        = 'd0         ;
    std__pe34__lane12_strm1_data        = 'h1234_5678 ;
    std__pe34__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe34__lane13_strm0_cntl        = 'd0         ;
    std__pe34__lane13_strm0_data        = 'h1234_5678 ;
    std__pe34__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe34__lane13_strm1_cntl        = 'd0         ;
    std__pe34__lane13_strm1_data        = 'h1234_5678 ;
    std__pe34__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe34__lane14_strm0_cntl        = 'd0         ;
    std__pe34__lane14_strm0_data        = 'h1234_5678 ;
    std__pe34__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe34__lane14_strm1_cntl        = 'd0         ;
    std__pe34__lane14_strm1_data        = 'h1234_5678 ;
    std__pe34__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe34__lane15_strm0_cntl        = 'd0         ;
    std__pe34__lane15_strm0_data        = 'h1234_5678 ;
    std__pe34__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe34__lane15_strm1_cntl        = 'd0         ;
    std__pe34__lane15_strm1_data        = 'h1234_5678 ;
    std__pe34__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe34__lane16_strm0_cntl        = 'd0         ;
    std__pe34__lane16_strm0_data        = 'h1234_5678 ;
    std__pe34__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe34__lane16_strm1_cntl        = 'd0         ;
    std__pe34__lane16_strm1_data        = 'h1234_5678 ;
    std__pe34__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe34__lane17_strm0_cntl        = 'd0         ;
    std__pe34__lane17_strm0_data        = 'h1234_5678 ;
    std__pe34__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe34__lane17_strm1_cntl        = 'd0         ;
    std__pe34__lane17_strm1_data        = 'h1234_5678 ;
    std__pe34__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe34__lane18_strm0_cntl        = 'd0         ;
    std__pe34__lane18_strm0_data        = 'h1234_5678 ;
    std__pe34__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe34__lane18_strm1_cntl        = 'd0         ;
    std__pe34__lane18_strm1_data        = 'h1234_5678 ;
    std__pe34__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe34__lane19_strm0_cntl        = 'd0         ;
    std__pe34__lane19_strm0_data        = 'h1234_5678 ;
    std__pe34__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe34__lane19_strm1_cntl        = 'd0         ;
    std__pe34__lane19_strm1_data        = 'h1234_5678 ;
    std__pe34__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe34__lane20_strm0_cntl        = 'd0         ;
    std__pe34__lane20_strm0_data        = 'h1234_5678 ;
    std__pe34__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe34__lane20_strm1_cntl        = 'd0         ;
    std__pe34__lane20_strm1_data        = 'h1234_5678 ;
    std__pe34__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe34__lane21_strm0_cntl        = 'd0         ;
    std__pe34__lane21_strm0_data        = 'h1234_5678 ;
    std__pe34__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe34__lane21_strm1_cntl        = 'd0         ;
    std__pe34__lane21_strm1_data        = 'h1234_5678 ;
    std__pe34__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe34__lane22_strm0_cntl        = 'd0         ;
    std__pe34__lane22_strm0_data        = 'h1234_5678 ;
    std__pe34__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe34__lane22_strm1_cntl        = 'd0         ;
    std__pe34__lane22_strm1_data        = 'h1234_5678 ;
    std__pe34__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe34__lane23_strm0_cntl        = 'd0         ;
    std__pe34__lane23_strm0_data        = 'h1234_5678 ;
    std__pe34__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe34__lane23_strm1_cntl        = 'd0         ;
    std__pe34__lane23_strm1_data        = 'h1234_5678 ;
    std__pe34__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe34__lane24_strm0_cntl        = 'd0         ;
    std__pe34__lane24_strm0_data        = 'h1234_5678 ;
    std__pe34__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe34__lane24_strm1_cntl        = 'd0         ;
    std__pe34__lane24_strm1_data        = 'h1234_5678 ;
    std__pe34__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe34__lane25_strm0_cntl        = 'd0         ;
    std__pe34__lane25_strm0_data        = 'h1234_5678 ;
    std__pe34__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe34__lane25_strm1_cntl        = 'd0         ;
    std__pe34__lane25_strm1_data        = 'h1234_5678 ;
    std__pe34__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe34__lane26_strm0_cntl        = 'd0         ;
    std__pe34__lane26_strm0_data        = 'h1234_5678 ;
    std__pe34__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe34__lane26_strm1_cntl        = 'd0         ;
    std__pe34__lane26_strm1_data        = 'h1234_5678 ;
    std__pe34__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe34__lane27_strm0_cntl        = 'd0         ;
    std__pe34__lane27_strm0_data        = 'h1234_5678 ;
    std__pe34__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe34__lane27_strm1_cntl        = 'd0         ;
    std__pe34__lane27_strm1_data        = 'h1234_5678 ;
    std__pe34__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe34__lane28_strm0_cntl        = 'd0         ;
    std__pe34__lane28_strm0_data        = 'h1234_5678 ;
    std__pe34__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe34__lane28_strm1_cntl        = 'd0         ;
    std__pe34__lane28_strm1_data        = 'h1234_5678 ;
    std__pe34__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe34__lane29_strm0_cntl        = 'd0         ;
    std__pe34__lane29_strm0_data        = 'h1234_5678 ;
    std__pe34__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe34__lane29_strm1_cntl        = 'd0         ;
    std__pe34__lane29_strm1_data        = 'h1234_5678 ;
    std__pe34__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe34__lane30_strm0_cntl        = 'd0         ;
    std__pe34__lane30_strm0_data        = 'h1234_5678 ;
    std__pe34__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe34__lane30_strm1_cntl        = 'd0         ;
    std__pe34__lane30_strm1_data        = 'h1234_5678 ;
    std__pe34__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe34__lane31_strm0_cntl        = 'd0         ;
    std__pe34__lane31_strm0_data        = 'h1234_5678 ;
    std__pe34__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe34__lane31_strm1_cntl        = 'd0         ;
    std__pe34__lane31_strm1_data        = 'h1234_5678 ;
    std__pe34__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe35__lane0_strm0_cntl        = 'd0         ;
    std__pe35__lane0_strm0_data        = 'h1234_5678 ;
    std__pe35__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe35__lane0_strm1_cntl        = 'd0         ;
    std__pe35__lane0_strm1_data        = 'h1234_5678 ;
    std__pe35__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe35__lane1_strm0_cntl        = 'd0         ;
    std__pe35__lane1_strm0_data        = 'h1234_5678 ;
    std__pe35__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe35__lane1_strm1_cntl        = 'd0         ;
    std__pe35__lane1_strm1_data        = 'h1234_5678 ;
    std__pe35__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe35__lane2_strm0_cntl        = 'd0         ;
    std__pe35__lane2_strm0_data        = 'h1234_5678 ;
    std__pe35__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe35__lane2_strm1_cntl        = 'd0         ;
    std__pe35__lane2_strm1_data        = 'h1234_5678 ;
    std__pe35__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe35__lane3_strm0_cntl        = 'd0         ;
    std__pe35__lane3_strm0_data        = 'h1234_5678 ;
    std__pe35__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe35__lane3_strm1_cntl        = 'd0         ;
    std__pe35__lane3_strm1_data        = 'h1234_5678 ;
    std__pe35__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe35__lane4_strm0_cntl        = 'd0         ;
    std__pe35__lane4_strm0_data        = 'h1234_5678 ;
    std__pe35__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe35__lane4_strm1_cntl        = 'd0         ;
    std__pe35__lane4_strm1_data        = 'h1234_5678 ;
    std__pe35__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe35__lane5_strm0_cntl        = 'd0         ;
    std__pe35__lane5_strm0_data        = 'h1234_5678 ;
    std__pe35__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe35__lane5_strm1_cntl        = 'd0         ;
    std__pe35__lane5_strm1_data        = 'h1234_5678 ;
    std__pe35__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe35__lane6_strm0_cntl        = 'd0         ;
    std__pe35__lane6_strm0_data        = 'h1234_5678 ;
    std__pe35__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe35__lane6_strm1_cntl        = 'd0         ;
    std__pe35__lane6_strm1_data        = 'h1234_5678 ;
    std__pe35__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe35__lane7_strm0_cntl        = 'd0         ;
    std__pe35__lane7_strm0_data        = 'h1234_5678 ;
    std__pe35__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe35__lane7_strm1_cntl        = 'd0         ;
    std__pe35__lane7_strm1_data        = 'h1234_5678 ;
    std__pe35__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe35__lane8_strm0_cntl        = 'd0         ;
    std__pe35__lane8_strm0_data        = 'h1234_5678 ;
    std__pe35__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe35__lane8_strm1_cntl        = 'd0         ;
    std__pe35__lane8_strm1_data        = 'h1234_5678 ;
    std__pe35__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe35__lane9_strm0_cntl        = 'd0         ;
    std__pe35__lane9_strm0_data        = 'h1234_5678 ;
    std__pe35__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe35__lane9_strm1_cntl        = 'd0         ;
    std__pe35__lane9_strm1_data        = 'h1234_5678 ;
    std__pe35__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe35__lane10_strm0_cntl        = 'd0         ;
    std__pe35__lane10_strm0_data        = 'h1234_5678 ;
    std__pe35__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe35__lane10_strm1_cntl        = 'd0         ;
    std__pe35__lane10_strm1_data        = 'h1234_5678 ;
    std__pe35__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe35__lane11_strm0_cntl        = 'd0         ;
    std__pe35__lane11_strm0_data        = 'h1234_5678 ;
    std__pe35__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe35__lane11_strm1_cntl        = 'd0         ;
    std__pe35__lane11_strm1_data        = 'h1234_5678 ;
    std__pe35__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe35__lane12_strm0_cntl        = 'd0         ;
    std__pe35__lane12_strm0_data        = 'h1234_5678 ;
    std__pe35__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe35__lane12_strm1_cntl        = 'd0         ;
    std__pe35__lane12_strm1_data        = 'h1234_5678 ;
    std__pe35__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe35__lane13_strm0_cntl        = 'd0         ;
    std__pe35__lane13_strm0_data        = 'h1234_5678 ;
    std__pe35__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe35__lane13_strm1_cntl        = 'd0         ;
    std__pe35__lane13_strm1_data        = 'h1234_5678 ;
    std__pe35__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe35__lane14_strm0_cntl        = 'd0         ;
    std__pe35__lane14_strm0_data        = 'h1234_5678 ;
    std__pe35__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe35__lane14_strm1_cntl        = 'd0         ;
    std__pe35__lane14_strm1_data        = 'h1234_5678 ;
    std__pe35__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe35__lane15_strm0_cntl        = 'd0         ;
    std__pe35__lane15_strm0_data        = 'h1234_5678 ;
    std__pe35__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe35__lane15_strm1_cntl        = 'd0         ;
    std__pe35__lane15_strm1_data        = 'h1234_5678 ;
    std__pe35__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe35__lane16_strm0_cntl        = 'd0         ;
    std__pe35__lane16_strm0_data        = 'h1234_5678 ;
    std__pe35__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe35__lane16_strm1_cntl        = 'd0         ;
    std__pe35__lane16_strm1_data        = 'h1234_5678 ;
    std__pe35__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe35__lane17_strm0_cntl        = 'd0         ;
    std__pe35__lane17_strm0_data        = 'h1234_5678 ;
    std__pe35__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe35__lane17_strm1_cntl        = 'd0         ;
    std__pe35__lane17_strm1_data        = 'h1234_5678 ;
    std__pe35__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe35__lane18_strm0_cntl        = 'd0         ;
    std__pe35__lane18_strm0_data        = 'h1234_5678 ;
    std__pe35__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe35__lane18_strm1_cntl        = 'd0         ;
    std__pe35__lane18_strm1_data        = 'h1234_5678 ;
    std__pe35__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe35__lane19_strm0_cntl        = 'd0         ;
    std__pe35__lane19_strm0_data        = 'h1234_5678 ;
    std__pe35__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe35__lane19_strm1_cntl        = 'd0         ;
    std__pe35__lane19_strm1_data        = 'h1234_5678 ;
    std__pe35__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe35__lane20_strm0_cntl        = 'd0         ;
    std__pe35__lane20_strm0_data        = 'h1234_5678 ;
    std__pe35__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe35__lane20_strm1_cntl        = 'd0         ;
    std__pe35__lane20_strm1_data        = 'h1234_5678 ;
    std__pe35__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe35__lane21_strm0_cntl        = 'd0         ;
    std__pe35__lane21_strm0_data        = 'h1234_5678 ;
    std__pe35__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe35__lane21_strm1_cntl        = 'd0         ;
    std__pe35__lane21_strm1_data        = 'h1234_5678 ;
    std__pe35__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe35__lane22_strm0_cntl        = 'd0         ;
    std__pe35__lane22_strm0_data        = 'h1234_5678 ;
    std__pe35__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe35__lane22_strm1_cntl        = 'd0         ;
    std__pe35__lane22_strm1_data        = 'h1234_5678 ;
    std__pe35__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe35__lane23_strm0_cntl        = 'd0         ;
    std__pe35__lane23_strm0_data        = 'h1234_5678 ;
    std__pe35__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe35__lane23_strm1_cntl        = 'd0         ;
    std__pe35__lane23_strm1_data        = 'h1234_5678 ;
    std__pe35__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe35__lane24_strm0_cntl        = 'd0         ;
    std__pe35__lane24_strm0_data        = 'h1234_5678 ;
    std__pe35__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe35__lane24_strm1_cntl        = 'd0         ;
    std__pe35__lane24_strm1_data        = 'h1234_5678 ;
    std__pe35__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe35__lane25_strm0_cntl        = 'd0         ;
    std__pe35__lane25_strm0_data        = 'h1234_5678 ;
    std__pe35__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe35__lane25_strm1_cntl        = 'd0         ;
    std__pe35__lane25_strm1_data        = 'h1234_5678 ;
    std__pe35__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe35__lane26_strm0_cntl        = 'd0         ;
    std__pe35__lane26_strm0_data        = 'h1234_5678 ;
    std__pe35__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe35__lane26_strm1_cntl        = 'd0         ;
    std__pe35__lane26_strm1_data        = 'h1234_5678 ;
    std__pe35__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe35__lane27_strm0_cntl        = 'd0         ;
    std__pe35__lane27_strm0_data        = 'h1234_5678 ;
    std__pe35__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe35__lane27_strm1_cntl        = 'd0         ;
    std__pe35__lane27_strm1_data        = 'h1234_5678 ;
    std__pe35__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe35__lane28_strm0_cntl        = 'd0         ;
    std__pe35__lane28_strm0_data        = 'h1234_5678 ;
    std__pe35__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe35__lane28_strm1_cntl        = 'd0         ;
    std__pe35__lane28_strm1_data        = 'h1234_5678 ;
    std__pe35__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe35__lane29_strm0_cntl        = 'd0         ;
    std__pe35__lane29_strm0_data        = 'h1234_5678 ;
    std__pe35__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe35__lane29_strm1_cntl        = 'd0         ;
    std__pe35__lane29_strm1_data        = 'h1234_5678 ;
    std__pe35__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe35__lane30_strm0_cntl        = 'd0         ;
    std__pe35__lane30_strm0_data        = 'h1234_5678 ;
    std__pe35__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe35__lane30_strm1_cntl        = 'd0         ;
    std__pe35__lane30_strm1_data        = 'h1234_5678 ;
    std__pe35__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe35__lane31_strm0_cntl        = 'd0         ;
    std__pe35__lane31_strm0_data        = 'h1234_5678 ;
    std__pe35__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe35__lane31_strm1_cntl        = 'd0         ;
    std__pe35__lane31_strm1_data        = 'h1234_5678 ;
    std__pe35__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe36__lane0_strm0_cntl        = 'd0         ;
    std__pe36__lane0_strm0_data        = 'h1234_5678 ;
    std__pe36__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe36__lane0_strm1_cntl        = 'd0         ;
    std__pe36__lane0_strm1_data        = 'h1234_5678 ;
    std__pe36__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe36__lane1_strm0_cntl        = 'd0         ;
    std__pe36__lane1_strm0_data        = 'h1234_5678 ;
    std__pe36__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe36__lane1_strm1_cntl        = 'd0         ;
    std__pe36__lane1_strm1_data        = 'h1234_5678 ;
    std__pe36__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe36__lane2_strm0_cntl        = 'd0         ;
    std__pe36__lane2_strm0_data        = 'h1234_5678 ;
    std__pe36__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe36__lane2_strm1_cntl        = 'd0         ;
    std__pe36__lane2_strm1_data        = 'h1234_5678 ;
    std__pe36__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe36__lane3_strm0_cntl        = 'd0         ;
    std__pe36__lane3_strm0_data        = 'h1234_5678 ;
    std__pe36__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe36__lane3_strm1_cntl        = 'd0         ;
    std__pe36__lane3_strm1_data        = 'h1234_5678 ;
    std__pe36__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe36__lane4_strm0_cntl        = 'd0         ;
    std__pe36__lane4_strm0_data        = 'h1234_5678 ;
    std__pe36__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe36__lane4_strm1_cntl        = 'd0         ;
    std__pe36__lane4_strm1_data        = 'h1234_5678 ;
    std__pe36__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe36__lane5_strm0_cntl        = 'd0         ;
    std__pe36__lane5_strm0_data        = 'h1234_5678 ;
    std__pe36__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe36__lane5_strm1_cntl        = 'd0         ;
    std__pe36__lane5_strm1_data        = 'h1234_5678 ;
    std__pe36__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe36__lane6_strm0_cntl        = 'd0         ;
    std__pe36__lane6_strm0_data        = 'h1234_5678 ;
    std__pe36__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe36__lane6_strm1_cntl        = 'd0         ;
    std__pe36__lane6_strm1_data        = 'h1234_5678 ;
    std__pe36__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe36__lane7_strm0_cntl        = 'd0         ;
    std__pe36__lane7_strm0_data        = 'h1234_5678 ;
    std__pe36__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe36__lane7_strm1_cntl        = 'd0         ;
    std__pe36__lane7_strm1_data        = 'h1234_5678 ;
    std__pe36__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe36__lane8_strm0_cntl        = 'd0         ;
    std__pe36__lane8_strm0_data        = 'h1234_5678 ;
    std__pe36__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe36__lane8_strm1_cntl        = 'd0         ;
    std__pe36__lane8_strm1_data        = 'h1234_5678 ;
    std__pe36__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe36__lane9_strm0_cntl        = 'd0         ;
    std__pe36__lane9_strm0_data        = 'h1234_5678 ;
    std__pe36__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe36__lane9_strm1_cntl        = 'd0         ;
    std__pe36__lane9_strm1_data        = 'h1234_5678 ;
    std__pe36__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe36__lane10_strm0_cntl        = 'd0         ;
    std__pe36__lane10_strm0_data        = 'h1234_5678 ;
    std__pe36__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe36__lane10_strm1_cntl        = 'd0         ;
    std__pe36__lane10_strm1_data        = 'h1234_5678 ;
    std__pe36__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe36__lane11_strm0_cntl        = 'd0         ;
    std__pe36__lane11_strm0_data        = 'h1234_5678 ;
    std__pe36__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe36__lane11_strm1_cntl        = 'd0         ;
    std__pe36__lane11_strm1_data        = 'h1234_5678 ;
    std__pe36__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe36__lane12_strm0_cntl        = 'd0         ;
    std__pe36__lane12_strm0_data        = 'h1234_5678 ;
    std__pe36__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe36__lane12_strm1_cntl        = 'd0         ;
    std__pe36__lane12_strm1_data        = 'h1234_5678 ;
    std__pe36__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe36__lane13_strm0_cntl        = 'd0         ;
    std__pe36__lane13_strm0_data        = 'h1234_5678 ;
    std__pe36__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe36__lane13_strm1_cntl        = 'd0         ;
    std__pe36__lane13_strm1_data        = 'h1234_5678 ;
    std__pe36__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe36__lane14_strm0_cntl        = 'd0         ;
    std__pe36__lane14_strm0_data        = 'h1234_5678 ;
    std__pe36__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe36__lane14_strm1_cntl        = 'd0         ;
    std__pe36__lane14_strm1_data        = 'h1234_5678 ;
    std__pe36__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe36__lane15_strm0_cntl        = 'd0         ;
    std__pe36__lane15_strm0_data        = 'h1234_5678 ;
    std__pe36__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe36__lane15_strm1_cntl        = 'd0         ;
    std__pe36__lane15_strm1_data        = 'h1234_5678 ;
    std__pe36__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe36__lane16_strm0_cntl        = 'd0         ;
    std__pe36__lane16_strm0_data        = 'h1234_5678 ;
    std__pe36__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe36__lane16_strm1_cntl        = 'd0         ;
    std__pe36__lane16_strm1_data        = 'h1234_5678 ;
    std__pe36__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe36__lane17_strm0_cntl        = 'd0         ;
    std__pe36__lane17_strm0_data        = 'h1234_5678 ;
    std__pe36__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe36__lane17_strm1_cntl        = 'd0         ;
    std__pe36__lane17_strm1_data        = 'h1234_5678 ;
    std__pe36__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe36__lane18_strm0_cntl        = 'd0         ;
    std__pe36__lane18_strm0_data        = 'h1234_5678 ;
    std__pe36__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe36__lane18_strm1_cntl        = 'd0         ;
    std__pe36__lane18_strm1_data        = 'h1234_5678 ;
    std__pe36__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe36__lane19_strm0_cntl        = 'd0         ;
    std__pe36__lane19_strm0_data        = 'h1234_5678 ;
    std__pe36__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe36__lane19_strm1_cntl        = 'd0         ;
    std__pe36__lane19_strm1_data        = 'h1234_5678 ;
    std__pe36__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe36__lane20_strm0_cntl        = 'd0         ;
    std__pe36__lane20_strm0_data        = 'h1234_5678 ;
    std__pe36__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe36__lane20_strm1_cntl        = 'd0         ;
    std__pe36__lane20_strm1_data        = 'h1234_5678 ;
    std__pe36__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe36__lane21_strm0_cntl        = 'd0         ;
    std__pe36__lane21_strm0_data        = 'h1234_5678 ;
    std__pe36__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe36__lane21_strm1_cntl        = 'd0         ;
    std__pe36__lane21_strm1_data        = 'h1234_5678 ;
    std__pe36__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe36__lane22_strm0_cntl        = 'd0         ;
    std__pe36__lane22_strm0_data        = 'h1234_5678 ;
    std__pe36__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe36__lane22_strm1_cntl        = 'd0         ;
    std__pe36__lane22_strm1_data        = 'h1234_5678 ;
    std__pe36__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe36__lane23_strm0_cntl        = 'd0         ;
    std__pe36__lane23_strm0_data        = 'h1234_5678 ;
    std__pe36__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe36__lane23_strm1_cntl        = 'd0         ;
    std__pe36__lane23_strm1_data        = 'h1234_5678 ;
    std__pe36__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe36__lane24_strm0_cntl        = 'd0         ;
    std__pe36__lane24_strm0_data        = 'h1234_5678 ;
    std__pe36__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe36__lane24_strm1_cntl        = 'd0         ;
    std__pe36__lane24_strm1_data        = 'h1234_5678 ;
    std__pe36__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe36__lane25_strm0_cntl        = 'd0         ;
    std__pe36__lane25_strm0_data        = 'h1234_5678 ;
    std__pe36__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe36__lane25_strm1_cntl        = 'd0         ;
    std__pe36__lane25_strm1_data        = 'h1234_5678 ;
    std__pe36__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe36__lane26_strm0_cntl        = 'd0         ;
    std__pe36__lane26_strm0_data        = 'h1234_5678 ;
    std__pe36__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe36__lane26_strm1_cntl        = 'd0         ;
    std__pe36__lane26_strm1_data        = 'h1234_5678 ;
    std__pe36__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe36__lane27_strm0_cntl        = 'd0         ;
    std__pe36__lane27_strm0_data        = 'h1234_5678 ;
    std__pe36__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe36__lane27_strm1_cntl        = 'd0         ;
    std__pe36__lane27_strm1_data        = 'h1234_5678 ;
    std__pe36__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe36__lane28_strm0_cntl        = 'd0         ;
    std__pe36__lane28_strm0_data        = 'h1234_5678 ;
    std__pe36__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe36__lane28_strm1_cntl        = 'd0         ;
    std__pe36__lane28_strm1_data        = 'h1234_5678 ;
    std__pe36__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe36__lane29_strm0_cntl        = 'd0         ;
    std__pe36__lane29_strm0_data        = 'h1234_5678 ;
    std__pe36__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe36__lane29_strm1_cntl        = 'd0         ;
    std__pe36__lane29_strm1_data        = 'h1234_5678 ;
    std__pe36__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe36__lane30_strm0_cntl        = 'd0         ;
    std__pe36__lane30_strm0_data        = 'h1234_5678 ;
    std__pe36__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe36__lane30_strm1_cntl        = 'd0         ;
    std__pe36__lane30_strm1_data        = 'h1234_5678 ;
    std__pe36__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe36__lane31_strm0_cntl        = 'd0         ;
    std__pe36__lane31_strm0_data        = 'h1234_5678 ;
    std__pe36__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe36__lane31_strm1_cntl        = 'd0         ;
    std__pe36__lane31_strm1_data        = 'h1234_5678 ;
    std__pe36__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe37__lane0_strm0_cntl        = 'd0         ;
    std__pe37__lane0_strm0_data        = 'h1234_5678 ;
    std__pe37__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe37__lane0_strm1_cntl        = 'd0         ;
    std__pe37__lane0_strm1_data        = 'h1234_5678 ;
    std__pe37__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe37__lane1_strm0_cntl        = 'd0         ;
    std__pe37__lane1_strm0_data        = 'h1234_5678 ;
    std__pe37__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe37__lane1_strm1_cntl        = 'd0         ;
    std__pe37__lane1_strm1_data        = 'h1234_5678 ;
    std__pe37__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe37__lane2_strm0_cntl        = 'd0         ;
    std__pe37__lane2_strm0_data        = 'h1234_5678 ;
    std__pe37__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe37__lane2_strm1_cntl        = 'd0         ;
    std__pe37__lane2_strm1_data        = 'h1234_5678 ;
    std__pe37__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe37__lane3_strm0_cntl        = 'd0         ;
    std__pe37__lane3_strm0_data        = 'h1234_5678 ;
    std__pe37__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe37__lane3_strm1_cntl        = 'd0         ;
    std__pe37__lane3_strm1_data        = 'h1234_5678 ;
    std__pe37__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe37__lane4_strm0_cntl        = 'd0         ;
    std__pe37__lane4_strm0_data        = 'h1234_5678 ;
    std__pe37__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe37__lane4_strm1_cntl        = 'd0         ;
    std__pe37__lane4_strm1_data        = 'h1234_5678 ;
    std__pe37__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe37__lane5_strm0_cntl        = 'd0         ;
    std__pe37__lane5_strm0_data        = 'h1234_5678 ;
    std__pe37__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe37__lane5_strm1_cntl        = 'd0         ;
    std__pe37__lane5_strm1_data        = 'h1234_5678 ;
    std__pe37__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe37__lane6_strm0_cntl        = 'd0         ;
    std__pe37__lane6_strm0_data        = 'h1234_5678 ;
    std__pe37__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe37__lane6_strm1_cntl        = 'd0         ;
    std__pe37__lane6_strm1_data        = 'h1234_5678 ;
    std__pe37__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe37__lane7_strm0_cntl        = 'd0         ;
    std__pe37__lane7_strm0_data        = 'h1234_5678 ;
    std__pe37__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe37__lane7_strm1_cntl        = 'd0         ;
    std__pe37__lane7_strm1_data        = 'h1234_5678 ;
    std__pe37__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe37__lane8_strm0_cntl        = 'd0         ;
    std__pe37__lane8_strm0_data        = 'h1234_5678 ;
    std__pe37__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe37__lane8_strm1_cntl        = 'd0         ;
    std__pe37__lane8_strm1_data        = 'h1234_5678 ;
    std__pe37__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe37__lane9_strm0_cntl        = 'd0         ;
    std__pe37__lane9_strm0_data        = 'h1234_5678 ;
    std__pe37__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe37__lane9_strm1_cntl        = 'd0         ;
    std__pe37__lane9_strm1_data        = 'h1234_5678 ;
    std__pe37__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe37__lane10_strm0_cntl        = 'd0         ;
    std__pe37__lane10_strm0_data        = 'h1234_5678 ;
    std__pe37__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe37__lane10_strm1_cntl        = 'd0         ;
    std__pe37__lane10_strm1_data        = 'h1234_5678 ;
    std__pe37__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe37__lane11_strm0_cntl        = 'd0         ;
    std__pe37__lane11_strm0_data        = 'h1234_5678 ;
    std__pe37__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe37__lane11_strm1_cntl        = 'd0         ;
    std__pe37__lane11_strm1_data        = 'h1234_5678 ;
    std__pe37__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe37__lane12_strm0_cntl        = 'd0         ;
    std__pe37__lane12_strm0_data        = 'h1234_5678 ;
    std__pe37__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe37__lane12_strm1_cntl        = 'd0         ;
    std__pe37__lane12_strm1_data        = 'h1234_5678 ;
    std__pe37__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe37__lane13_strm0_cntl        = 'd0         ;
    std__pe37__lane13_strm0_data        = 'h1234_5678 ;
    std__pe37__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe37__lane13_strm1_cntl        = 'd0         ;
    std__pe37__lane13_strm1_data        = 'h1234_5678 ;
    std__pe37__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe37__lane14_strm0_cntl        = 'd0         ;
    std__pe37__lane14_strm0_data        = 'h1234_5678 ;
    std__pe37__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe37__lane14_strm1_cntl        = 'd0         ;
    std__pe37__lane14_strm1_data        = 'h1234_5678 ;
    std__pe37__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe37__lane15_strm0_cntl        = 'd0         ;
    std__pe37__lane15_strm0_data        = 'h1234_5678 ;
    std__pe37__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe37__lane15_strm1_cntl        = 'd0         ;
    std__pe37__lane15_strm1_data        = 'h1234_5678 ;
    std__pe37__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe37__lane16_strm0_cntl        = 'd0         ;
    std__pe37__lane16_strm0_data        = 'h1234_5678 ;
    std__pe37__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe37__lane16_strm1_cntl        = 'd0         ;
    std__pe37__lane16_strm1_data        = 'h1234_5678 ;
    std__pe37__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe37__lane17_strm0_cntl        = 'd0         ;
    std__pe37__lane17_strm0_data        = 'h1234_5678 ;
    std__pe37__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe37__lane17_strm1_cntl        = 'd0         ;
    std__pe37__lane17_strm1_data        = 'h1234_5678 ;
    std__pe37__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe37__lane18_strm0_cntl        = 'd0         ;
    std__pe37__lane18_strm0_data        = 'h1234_5678 ;
    std__pe37__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe37__lane18_strm1_cntl        = 'd0         ;
    std__pe37__lane18_strm1_data        = 'h1234_5678 ;
    std__pe37__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe37__lane19_strm0_cntl        = 'd0         ;
    std__pe37__lane19_strm0_data        = 'h1234_5678 ;
    std__pe37__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe37__lane19_strm1_cntl        = 'd0         ;
    std__pe37__lane19_strm1_data        = 'h1234_5678 ;
    std__pe37__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe37__lane20_strm0_cntl        = 'd0         ;
    std__pe37__lane20_strm0_data        = 'h1234_5678 ;
    std__pe37__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe37__lane20_strm1_cntl        = 'd0         ;
    std__pe37__lane20_strm1_data        = 'h1234_5678 ;
    std__pe37__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe37__lane21_strm0_cntl        = 'd0         ;
    std__pe37__lane21_strm0_data        = 'h1234_5678 ;
    std__pe37__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe37__lane21_strm1_cntl        = 'd0         ;
    std__pe37__lane21_strm1_data        = 'h1234_5678 ;
    std__pe37__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe37__lane22_strm0_cntl        = 'd0         ;
    std__pe37__lane22_strm0_data        = 'h1234_5678 ;
    std__pe37__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe37__lane22_strm1_cntl        = 'd0         ;
    std__pe37__lane22_strm1_data        = 'h1234_5678 ;
    std__pe37__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe37__lane23_strm0_cntl        = 'd0         ;
    std__pe37__lane23_strm0_data        = 'h1234_5678 ;
    std__pe37__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe37__lane23_strm1_cntl        = 'd0         ;
    std__pe37__lane23_strm1_data        = 'h1234_5678 ;
    std__pe37__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe37__lane24_strm0_cntl        = 'd0         ;
    std__pe37__lane24_strm0_data        = 'h1234_5678 ;
    std__pe37__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe37__lane24_strm1_cntl        = 'd0         ;
    std__pe37__lane24_strm1_data        = 'h1234_5678 ;
    std__pe37__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe37__lane25_strm0_cntl        = 'd0         ;
    std__pe37__lane25_strm0_data        = 'h1234_5678 ;
    std__pe37__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe37__lane25_strm1_cntl        = 'd0         ;
    std__pe37__lane25_strm1_data        = 'h1234_5678 ;
    std__pe37__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe37__lane26_strm0_cntl        = 'd0         ;
    std__pe37__lane26_strm0_data        = 'h1234_5678 ;
    std__pe37__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe37__lane26_strm1_cntl        = 'd0         ;
    std__pe37__lane26_strm1_data        = 'h1234_5678 ;
    std__pe37__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe37__lane27_strm0_cntl        = 'd0         ;
    std__pe37__lane27_strm0_data        = 'h1234_5678 ;
    std__pe37__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe37__lane27_strm1_cntl        = 'd0         ;
    std__pe37__lane27_strm1_data        = 'h1234_5678 ;
    std__pe37__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe37__lane28_strm0_cntl        = 'd0         ;
    std__pe37__lane28_strm0_data        = 'h1234_5678 ;
    std__pe37__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe37__lane28_strm1_cntl        = 'd0         ;
    std__pe37__lane28_strm1_data        = 'h1234_5678 ;
    std__pe37__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe37__lane29_strm0_cntl        = 'd0         ;
    std__pe37__lane29_strm0_data        = 'h1234_5678 ;
    std__pe37__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe37__lane29_strm1_cntl        = 'd0         ;
    std__pe37__lane29_strm1_data        = 'h1234_5678 ;
    std__pe37__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe37__lane30_strm0_cntl        = 'd0         ;
    std__pe37__lane30_strm0_data        = 'h1234_5678 ;
    std__pe37__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe37__lane30_strm1_cntl        = 'd0         ;
    std__pe37__lane30_strm1_data        = 'h1234_5678 ;
    std__pe37__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe37__lane31_strm0_cntl        = 'd0         ;
    std__pe37__lane31_strm0_data        = 'h1234_5678 ;
    std__pe37__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe37__lane31_strm1_cntl        = 'd0         ;
    std__pe37__lane31_strm1_data        = 'h1234_5678 ;
    std__pe37__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe38__lane0_strm0_cntl        = 'd0         ;
    std__pe38__lane0_strm0_data        = 'h1234_5678 ;
    std__pe38__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe38__lane0_strm1_cntl        = 'd0         ;
    std__pe38__lane0_strm1_data        = 'h1234_5678 ;
    std__pe38__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe38__lane1_strm0_cntl        = 'd0         ;
    std__pe38__lane1_strm0_data        = 'h1234_5678 ;
    std__pe38__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe38__lane1_strm1_cntl        = 'd0         ;
    std__pe38__lane1_strm1_data        = 'h1234_5678 ;
    std__pe38__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe38__lane2_strm0_cntl        = 'd0         ;
    std__pe38__lane2_strm0_data        = 'h1234_5678 ;
    std__pe38__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe38__lane2_strm1_cntl        = 'd0         ;
    std__pe38__lane2_strm1_data        = 'h1234_5678 ;
    std__pe38__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe38__lane3_strm0_cntl        = 'd0         ;
    std__pe38__lane3_strm0_data        = 'h1234_5678 ;
    std__pe38__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe38__lane3_strm1_cntl        = 'd0         ;
    std__pe38__lane3_strm1_data        = 'h1234_5678 ;
    std__pe38__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe38__lane4_strm0_cntl        = 'd0         ;
    std__pe38__lane4_strm0_data        = 'h1234_5678 ;
    std__pe38__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe38__lane4_strm1_cntl        = 'd0         ;
    std__pe38__lane4_strm1_data        = 'h1234_5678 ;
    std__pe38__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe38__lane5_strm0_cntl        = 'd0         ;
    std__pe38__lane5_strm0_data        = 'h1234_5678 ;
    std__pe38__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe38__lane5_strm1_cntl        = 'd0         ;
    std__pe38__lane5_strm1_data        = 'h1234_5678 ;
    std__pe38__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe38__lane6_strm0_cntl        = 'd0         ;
    std__pe38__lane6_strm0_data        = 'h1234_5678 ;
    std__pe38__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe38__lane6_strm1_cntl        = 'd0         ;
    std__pe38__lane6_strm1_data        = 'h1234_5678 ;
    std__pe38__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe38__lane7_strm0_cntl        = 'd0         ;
    std__pe38__lane7_strm0_data        = 'h1234_5678 ;
    std__pe38__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe38__lane7_strm1_cntl        = 'd0         ;
    std__pe38__lane7_strm1_data        = 'h1234_5678 ;
    std__pe38__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe38__lane8_strm0_cntl        = 'd0         ;
    std__pe38__lane8_strm0_data        = 'h1234_5678 ;
    std__pe38__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe38__lane8_strm1_cntl        = 'd0         ;
    std__pe38__lane8_strm1_data        = 'h1234_5678 ;
    std__pe38__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe38__lane9_strm0_cntl        = 'd0         ;
    std__pe38__lane9_strm0_data        = 'h1234_5678 ;
    std__pe38__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe38__lane9_strm1_cntl        = 'd0         ;
    std__pe38__lane9_strm1_data        = 'h1234_5678 ;
    std__pe38__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe38__lane10_strm0_cntl        = 'd0         ;
    std__pe38__lane10_strm0_data        = 'h1234_5678 ;
    std__pe38__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe38__lane10_strm1_cntl        = 'd0         ;
    std__pe38__lane10_strm1_data        = 'h1234_5678 ;
    std__pe38__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe38__lane11_strm0_cntl        = 'd0         ;
    std__pe38__lane11_strm0_data        = 'h1234_5678 ;
    std__pe38__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe38__lane11_strm1_cntl        = 'd0         ;
    std__pe38__lane11_strm1_data        = 'h1234_5678 ;
    std__pe38__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe38__lane12_strm0_cntl        = 'd0         ;
    std__pe38__lane12_strm0_data        = 'h1234_5678 ;
    std__pe38__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe38__lane12_strm1_cntl        = 'd0         ;
    std__pe38__lane12_strm1_data        = 'h1234_5678 ;
    std__pe38__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe38__lane13_strm0_cntl        = 'd0         ;
    std__pe38__lane13_strm0_data        = 'h1234_5678 ;
    std__pe38__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe38__lane13_strm1_cntl        = 'd0         ;
    std__pe38__lane13_strm1_data        = 'h1234_5678 ;
    std__pe38__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe38__lane14_strm0_cntl        = 'd0         ;
    std__pe38__lane14_strm0_data        = 'h1234_5678 ;
    std__pe38__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe38__lane14_strm1_cntl        = 'd0         ;
    std__pe38__lane14_strm1_data        = 'h1234_5678 ;
    std__pe38__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe38__lane15_strm0_cntl        = 'd0         ;
    std__pe38__lane15_strm0_data        = 'h1234_5678 ;
    std__pe38__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe38__lane15_strm1_cntl        = 'd0         ;
    std__pe38__lane15_strm1_data        = 'h1234_5678 ;
    std__pe38__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe38__lane16_strm0_cntl        = 'd0         ;
    std__pe38__lane16_strm0_data        = 'h1234_5678 ;
    std__pe38__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe38__lane16_strm1_cntl        = 'd0         ;
    std__pe38__lane16_strm1_data        = 'h1234_5678 ;
    std__pe38__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe38__lane17_strm0_cntl        = 'd0         ;
    std__pe38__lane17_strm0_data        = 'h1234_5678 ;
    std__pe38__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe38__lane17_strm1_cntl        = 'd0         ;
    std__pe38__lane17_strm1_data        = 'h1234_5678 ;
    std__pe38__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe38__lane18_strm0_cntl        = 'd0         ;
    std__pe38__lane18_strm0_data        = 'h1234_5678 ;
    std__pe38__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe38__lane18_strm1_cntl        = 'd0         ;
    std__pe38__lane18_strm1_data        = 'h1234_5678 ;
    std__pe38__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe38__lane19_strm0_cntl        = 'd0         ;
    std__pe38__lane19_strm0_data        = 'h1234_5678 ;
    std__pe38__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe38__lane19_strm1_cntl        = 'd0         ;
    std__pe38__lane19_strm1_data        = 'h1234_5678 ;
    std__pe38__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe38__lane20_strm0_cntl        = 'd0         ;
    std__pe38__lane20_strm0_data        = 'h1234_5678 ;
    std__pe38__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe38__lane20_strm1_cntl        = 'd0         ;
    std__pe38__lane20_strm1_data        = 'h1234_5678 ;
    std__pe38__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe38__lane21_strm0_cntl        = 'd0         ;
    std__pe38__lane21_strm0_data        = 'h1234_5678 ;
    std__pe38__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe38__lane21_strm1_cntl        = 'd0         ;
    std__pe38__lane21_strm1_data        = 'h1234_5678 ;
    std__pe38__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe38__lane22_strm0_cntl        = 'd0         ;
    std__pe38__lane22_strm0_data        = 'h1234_5678 ;
    std__pe38__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe38__lane22_strm1_cntl        = 'd0         ;
    std__pe38__lane22_strm1_data        = 'h1234_5678 ;
    std__pe38__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe38__lane23_strm0_cntl        = 'd0         ;
    std__pe38__lane23_strm0_data        = 'h1234_5678 ;
    std__pe38__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe38__lane23_strm1_cntl        = 'd0         ;
    std__pe38__lane23_strm1_data        = 'h1234_5678 ;
    std__pe38__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe38__lane24_strm0_cntl        = 'd0         ;
    std__pe38__lane24_strm0_data        = 'h1234_5678 ;
    std__pe38__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe38__lane24_strm1_cntl        = 'd0         ;
    std__pe38__lane24_strm1_data        = 'h1234_5678 ;
    std__pe38__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe38__lane25_strm0_cntl        = 'd0         ;
    std__pe38__lane25_strm0_data        = 'h1234_5678 ;
    std__pe38__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe38__lane25_strm1_cntl        = 'd0         ;
    std__pe38__lane25_strm1_data        = 'h1234_5678 ;
    std__pe38__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe38__lane26_strm0_cntl        = 'd0         ;
    std__pe38__lane26_strm0_data        = 'h1234_5678 ;
    std__pe38__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe38__lane26_strm1_cntl        = 'd0         ;
    std__pe38__lane26_strm1_data        = 'h1234_5678 ;
    std__pe38__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe38__lane27_strm0_cntl        = 'd0         ;
    std__pe38__lane27_strm0_data        = 'h1234_5678 ;
    std__pe38__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe38__lane27_strm1_cntl        = 'd0         ;
    std__pe38__lane27_strm1_data        = 'h1234_5678 ;
    std__pe38__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe38__lane28_strm0_cntl        = 'd0         ;
    std__pe38__lane28_strm0_data        = 'h1234_5678 ;
    std__pe38__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe38__lane28_strm1_cntl        = 'd0         ;
    std__pe38__lane28_strm1_data        = 'h1234_5678 ;
    std__pe38__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe38__lane29_strm0_cntl        = 'd0         ;
    std__pe38__lane29_strm0_data        = 'h1234_5678 ;
    std__pe38__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe38__lane29_strm1_cntl        = 'd0         ;
    std__pe38__lane29_strm1_data        = 'h1234_5678 ;
    std__pe38__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe38__lane30_strm0_cntl        = 'd0         ;
    std__pe38__lane30_strm0_data        = 'h1234_5678 ;
    std__pe38__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe38__lane30_strm1_cntl        = 'd0         ;
    std__pe38__lane30_strm1_data        = 'h1234_5678 ;
    std__pe38__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe38__lane31_strm0_cntl        = 'd0         ;
    std__pe38__lane31_strm0_data        = 'h1234_5678 ;
    std__pe38__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe38__lane31_strm1_cntl        = 'd0         ;
    std__pe38__lane31_strm1_data        = 'h1234_5678 ;
    std__pe38__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe39__lane0_strm0_cntl        = 'd0         ;
    std__pe39__lane0_strm0_data        = 'h1234_5678 ;
    std__pe39__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe39__lane0_strm1_cntl        = 'd0         ;
    std__pe39__lane0_strm1_data        = 'h1234_5678 ;
    std__pe39__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe39__lane1_strm0_cntl        = 'd0         ;
    std__pe39__lane1_strm0_data        = 'h1234_5678 ;
    std__pe39__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe39__lane1_strm1_cntl        = 'd0         ;
    std__pe39__lane1_strm1_data        = 'h1234_5678 ;
    std__pe39__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe39__lane2_strm0_cntl        = 'd0         ;
    std__pe39__lane2_strm0_data        = 'h1234_5678 ;
    std__pe39__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe39__lane2_strm1_cntl        = 'd0         ;
    std__pe39__lane2_strm1_data        = 'h1234_5678 ;
    std__pe39__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe39__lane3_strm0_cntl        = 'd0         ;
    std__pe39__lane3_strm0_data        = 'h1234_5678 ;
    std__pe39__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe39__lane3_strm1_cntl        = 'd0         ;
    std__pe39__lane3_strm1_data        = 'h1234_5678 ;
    std__pe39__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe39__lane4_strm0_cntl        = 'd0         ;
    std__pe39__lane4_strm0_data        = 'h1234_5678 ;
    std__pe39__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe39__lane4_strm1_cntl        = 'd0         ;
    std__pe39__lane4_strm1_data        = 'h1234_5678 ;
    std__pe39__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe39__lane5_strm0_cntl        = 'd0         ;
    std__pe39__lane5_strm0_data        = 'h1234_5678 ;
    std__pe39__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe39__lane5_strm1_cntl        = 'd0         ;
    std__pe39__lane5_strm1_data        = 'h1234_5678 ;
    std__pe39__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe39__lane6_strm0_cntl        = 'd0         ;
    std__pe39__lane6_strm0_data        = 'h1234_5678 ;
    std__pe39__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe39__lane6_strm1_cntl        = 'd0         ;
    std__pe39__lane6_strm1_data        = 'h1234_5678 ;
    std__pe39__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe39__lane7_strm0_cntl        = 'd0         ;
    std__pe39__lane7_strm0_data        = 'h1234_5678 ;
    std__pe39__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe39__lane7_strm1_cntl        = 'd0         ;
    std__pe39__lane7_strm1_data        = 'h1234_5678 ;
    std__pe39__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe39__lane8_strm0_cntl        = 'd0         ;
    std__pe39__lane8_strm0_data        = 'h1234_5678 ;
    std__pe39__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe39__lane8_strm1_cntl        = 'd0         ;
    std__pe39__lane8_strm1_data        = 'h1234_5678 ;
    std__pe39__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe39__lane9_strm0_cntl        = 'd0         ;
    std__pe39__lane9_strm0_data        = 'h1234_5678 ;
    std__pe39__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe39__lane9_strm1_cntl        = 'd0         ;
    std__pe39__lane9_strm1_data        = 'h1234_5678 ;
    std__pe39__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe39__lane10_strm0_cntl        = 'd0         ;
    std__pe39__lane10_strm0_data        = 'h1234_5678 ;
    std__pe39__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe39__lane10_strm1_cntl        = 'd0         ;
    std__pe39__lane10_strm1_data        = 'h1234_5678 ;
    std__pe39__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe39__lane11_strm0_cntl        = 'd0         ;
    std__pe39__lane11_strm0_data        = 'h1234_5678 ;
    std__pe39__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe39__lane11_strm1_cntl        = 'd0         ;
    std__pe39__lane11_strm1_data        = 'h1234_5678 ;
    std__pe39__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe39__lane12_strm0_cntl        = 'd0         ;
    std__pe39__lane12_strm0_data        = 'h1234_5678 ;
    std__pe39__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe39__lane12_strm1_cntl        = 'd0         ;
    std__pe39__lane12_strm1_data        = 'h1234_5678 ;
    std__pe39__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe39__lane13_strm0_cntl        = 'd0         ;
    std__pe39__lane13_strm0_data        = 'h1234_5678 ;
    std__pe39__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe39__lane13_strm1_cntl        = 'd0         ;
    std__pe39__lane13_strm1_data        = 'h1234_5678 ;
    std__pe39__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe39__lane14_strm0_cntl        = 'd0         ;
    std__pe39__lane14_strm0_data        = 'h1234_5678 ;
    std__pe39__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe39__lane14_strm1_cntl        = 'd0         ;
    std__pe39__lane14_strm1_data        = 'h1234_5678 ;
    std__pe39__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe39__lane15_strm0_cntl        = 'd0         ;
    std__pe39__lane15_strm0_data        = 'h1234_5678 ;
    std__pe39__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe39__lane15_strm1_cntl        = 'd0         ;
    std__pe39__lane15_strm1_data        = 'h1234_5678 ;
    std__pe39__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe39__lane16_strm0_cntl        = 'd0         ;
    std__pe39__lane16_strm0_data        = 'h1234_5678 ;
    std__pe39__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe39__lane16_strm1_cntl        = 'd0         ;
    std__pe39__lane16_strm1_data        = 'h1234_5678 ;
    std__pe39__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe39__lane17_strm0_cntl        = 'd0         ;
    std__pe39__lane17_strm0_data        = 'h1234_5678 ;
    std__pe39__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe39__lane17_strm1_cntl        = 'd0         ;
    std__pe39__lane17_strm1_data        = 'h1234_5678 ;
    std__pe39__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe39__lane18_strm0_cntl        = 'd0         ;
    std__pe39__lane18_strm0_data        = 'h1234_5678 ;
    std__pe39__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe39__lane18_strm1_cntl        = 'd0         ;
    std__pe39__lane18_strm1_data        = 'h1234_5678 ;
    std__pe39__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe39__lane19_strm0_cntl        = 'd0         ;
    std__pe39__lane19_strm0_data        = 'h1234_5678 ;
    std__pe39__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe39__lane19_strm1_cntl        = 'd0         ;
    std__pe39__lane19_strm1_data        = 'h1234_5678 ;
    std__pe39__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe39__lane20_strm0_cntl        = 'd0         ;
    std__pe39__lane20_strm0_data        = 'h1234_5678 ;
    std__pe39__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe39__lane20_strm1_cntl        = 'd0         ;
    std__pe39__lane20_strm1_data        = 'h1234_5678 ;
    std__pe39__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe39__lane21_strm0_cntl        = 'd0         ;
    std__pe39__lane21_strm0_data        = 'h1234_5678 ;
    std__pe39__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe39__lane21_strm1_cntl        = 'd0         ;
    std__pe39__lane21_strm1_data        = 'h1234_5678 ;
    std__pe39__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe39__lane22_strm0_cntl        = 'd0         ;
    std__pe39__lane22_strm0_data        = 'h1234_5678 ;
    std__pe39__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe39__lane22_strm1_cntl        = 'd0         ;
    std__pe39__lane22_strm1_data        = 'h1234_5678 ;
    std__pe39__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe39__lane23_strm0_cntl        = 'd0         ;
    std__pe39__lane23_strm0_data        = 'h1234_5678 ;
    std__pe39__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe39__lane23_strm1_cntl        = 'd0         ;
    std__pe39__lane23_strm1_data        = 'h1234_5678 ;
    std__pe39__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe39__lane24_strm0_cntl        = 'd0         ;
    std__pe39__lane24_strm0_data        = 'h1234_5678 ;
    std__pe39__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe39__lane24_strm1_cntl        = 'd0         ;
    std__pe39__lane24_strm1_data        = 'h1234_5678 ;
    std__pe39__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe39__lane25_strm0_cntl        = 'd0         ;
    std__pe39__lane25_strm0_data        = 'h1234_5678 ;
    std__pe39__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe39__lane25_strm1_cntl        = 'd0         ;
    std__pe39__lane25_strm1_data        = 'h1234_5678 ;
    std__pe39__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe39__lane26_strm0_cntl        = 'd0         ;
    std__pe39__lane26_strm0_data        = 'h1234_5678 ;
    std__pe39__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe39__lane26_strm1_cntl        = 'd0         ;
    std__pe39__lane26_strm1_data        = 'h1234_5678 ;
    std__pe39__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe39__lane27_strm0_cntl        = 'd0         ;
    std__pe39__lane27_strm0_data        = 'h1234_5678 ;
    std__pe39__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe39__lane27_strm1_cntl        = 'd0         ;
    std__pe39__lane27_strm1_data        = 'h1234_5678 ;
    std__pe39__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe39__lane28_strm0_cntl        = 'd0         ;
    std__pe39__lane28_strm0_data        = 'h1234_5678 ;
    std__pe39__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe39__lane28_strm1_cntl        = 'd0         ;
    std__pe39__lane28_strm1_data        = 'h1234_5678 ;
    std__pe39__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe39__lane29_strm0_cntl        = 'd0         ;
    std__pe39__lane29_strm0_data        = 'h1234_5678 ;
    std__pe39__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe39__lane29_strm1_cntl        = 'd0         ;
    std__pe39__lane29_strm1_data        = 'h1234_5678 ;
    std__pe39__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe39__lane30_strm0_cntl        = 'd0         ;
    std__pe39__lane30_strm0_data        = 'h1234_5678 ;
    std__pe39__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe39__lane30_strm1_cntl        = 'd0         ;
    std__pe39__lane30_strm1_data        = 'h1234_5678 ;
    std__pe39__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe39__lane31_strm0_cntl        = 'd0         ;
    std__pe39__lane31_strm0_data        = 'h1234_5678 ;
    std__pe39__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe39__lane31_strm1_cntl        = 'd0         ;
    std__pe39__lane31_strm1_data        = 'h1234_5678 ;
    std__pe39__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe40__lane0_strm0_cntl        = 'd0         ;
    std__pe40__lane0_strm0_data        = 'h1234_5678 ;
    std__pe40__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe40__lane0_strm1_cntl        = 'd0         ;
    std__pe40__lane0_strm1_data        = 'h1234_5678 ;
    std__pe40__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe40__lane1_strm0_cntl        = 'd0         ;
    std__pe40__lane1_strm0_data        = 'h1234_5678 ;
    std__pe40__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe40__lane1_strm1_cntl        = 'd0         ;
    std__pe40__lane1_strm1_data        = 'h1234_5678 ;
    std__pe40__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe40__lane2_strm0_cntl        = 'd0         ;
    std__pe40__lane2_strm0_data        = 'h1234_5678 ;
    std__pe40__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe40__lane2_strm1_cntl        = 'd0         ;
    std__pe40__lane2_strm1_data        = 'h1234_5678 ;
    std__pe40__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe40__lane3_strm0_cntl        = 'd0         ;
    std__pe40__lane3_strm0_data        = 'h1234_5678 ;
    std__pe40__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe40__lane3_strm1_cntl        = 'd0         ;
    std__pe40__lane3_strm1_data        = 'h1234_5678 ;
    std__pe40__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe40__lane4_strm0_cntl        = 'd0         ;
    std__pe40__lane4_strm0_data        = 'h1234_5678 ;
    std__pe40__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe40__lane4_strm1_cntl        = 'd0         ;
    std__pe40__lane4_strm1_data        = 'h1234_5678 ;
    std__pe40__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe40__lane5_strm0_cntl        = 'd0         ;
    std__pe40__lane5_strm0_data        = 'h1234_5678 ;
    std__pe40__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe40__lane5_strm1_cntl        = 'd0         ;
    std__pe40__lane5_strm1_data        = 'h1234_5678 ;
    std__pe40__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe40__lane6_strm0_cntl        = 'd0         ;
    std__pe40__lane6_strm0_data        = 'h1234_5678 ;
    std__pe40__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe40__lane6_strm1_cntl        = 'd0         ;
    std__pe40__lane6_strm1_data        = 'h1234_5678 ;
    std__pe40__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe40__lane7_strm0_cntl        = 'd0         ;
    std__pe40__lane7_strm0_data        = 'h1234_5678 ;
    std__pe40__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe40__lane7_strm1_cntl        = 'd0         ;
    std__pe40__lane7_strm1_data        = 'h1234_5678 ;
    std__pe40__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe40__lane8_strm0_cntl        = 'd0         ;
    std__pe40__lane8_strm0_data        = 'h1234_5678 ;
    std__pe40__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe40__lane8_strm1_cntl        = 'd0         ;
    std__pe40__lane8_strm1_data        = 'h1234_5678 ;
    std__pe40__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe40__lane9_strm0_cntl        = 'd0         ;
    std__pe40__lane9_strm0_data        = 'h1234_5678 ;
    std__pe40__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe40__lane9_strm1_cntl        = 'd0         ;
    std__pe40__lane9_strm1_data        = 'h1234_5678 ;
    std__pe40__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe40__lane10_strm0_cntl        = 'd0         ;
    std__pe40__lane10_strm0_data        = 'h1234_5678 ;
    std__pe40__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe40__lane10_strm1_cntl        = 'd0         ;
    std__pe40__lane10_strm1_data        = 'h1234_5678 ;
    std__pe40__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe40__lane11_strm0_cntl        = 'd0         ;
    std__pe40__lane11_strm0_data        = 'h1234_5678 ;
    std__pe40__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe40__lane11_strm1_cntl        = 'd0         ;
    std__pe40__lane11_strm1_data        = 'h1234_5678 ;
    std__pe40__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe40__lane12_strm0_cntl        = 'd0         ;
    std__pe40__lane12_strm0_data        = 'h1234_5678 ;
    std__pe40__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe40__lane12_strm1_cntl        = 'd0         ;
    std__pe40__lane12_strm1_data        = 'h1234_5678 ;
    std__pe40__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe40__lane13_strm0_cntl        = 'd0         ;
    std__pe40__lane13_strm0_data        = 'h1234_5678 ;
    std__pe40__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe40__lane13_strm1_cntl        = 'd0         ;
    std__pe40__lane13_strm1_data        = 'h1234_5678 ;
    std__pe40__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe40__lane14_strm0_cntl        = 'd0         ;
    std__pe40__lane14_strm0_data        = 'h1234_5678 ;
    std__pe40__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe40__lane14_strm1_cntl        = 'd0         ;
    std__pe40__lane14_strm1_data        = 'h1234_5678 ;
    std__pe40__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe40__lane15_strm0_cntl        = 'd0         ;
    std__pe40__lane15_strm0_data        = 'h1234_5678 ;
    std__pe40__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe40__lane15_strm1_cntl        = 'd0         ;
    std__pe40__lane15_strm1_data        = 'h1234_5678 ;
    std__pe40__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe40__lane16_strm0_cntl        = 'd0         ;
    std__pe40__lane16_strm0_data        = 'h1234_5678 ;
    std__pe40__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe40__lane16_strm1_cntl        = 'd0         ;
    std__pe40__lane16_strm1_data        = 'h1234_5678 ;
    std__pe40__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe40__lane17_strm0_cntl        = 'd0         ;
    std__pe40__lane17_strm0_data        = 'h1234_5678 ;
    std__pe40__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe40__lane17_strm1_cntl        = 'd0         ;
    std__pe40__lane17_strm1_data        = 'h1234_5678 ;
    std__pe40__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe40__lane18_strm0_cntl        = 'd0         ;
    std__pe40__lane18_strm0_data        = 'h1234_5678 ;
    std__pe40__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe40__lane18_strm1_cntl        = 'd0         ;
    std__pe40__lane18_strm1_data        = 'h1234_5678 ;
    std__pe40__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe40__lane19_strm0_cntl        = 'd0         ;
    std__pe40__lane19_strm0_data        = 'h1234_5678 ;
    std__pe40__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe40__lane19_strm1_cntl        = 'd0         ;
    std__pe40__lane19_strm1_data        = 'h1234_5678 ;
    std__pe40__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe40__lane20_strm0_cntl        = 'd0         ;
    std__pe40__lane20_strm0_data        = 'h1234_5678 ;
    std__pe40__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe40__lane20_strm1_cntl        = 'd0         ;
    std__pe40__lane20_strm1_data        = 'h1234_5678 ;
    std__pe40__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe40__lane21_strm0_cntl        = 'd0         ;
    std__pe40__lane21_strm0_data        = 'h1234_5678 ;
    std__pe40__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe40__lane21_strm1_cntl        = 'd0         ;
    std__pe40__lane21_strm1_data        = 'h1234_5678 ;
    std__pe40__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe40__lane22_strm0_cntl        = 'd0         ;
    std__pe40__lane22_strm0_data        = 'h1234_5678 ;
    std__pe40__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe40__lane22_strm1_cntl        = 'd0         ;
    std__pe40__lane22_strm1_data        = 'h1234_5678 ;
    std__pe40__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe40__lane23_strm0_cntl        = 'd0         ;
    std__pe40__lane23_strm0_data        = 'h1234_5678 ;
    std__pe40__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe40__lane23_strm1_cntl        = 'd0         ;
    std__pe40__lane23_strm1_data        = 'h1234_5678 ;
    std__pe40__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe40__lane24_strm0_cntl        = 'd0         ;
    std__pe40__lane24_strm0_data        = 'h1234_5678 ;
    std__pe40__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe40__lane24_strm1_cntl        = 'd0         ;
    std__pe40__lane24_strm1_data        = 'h1234_5678 ;
    std__pe40__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe40__lane25_strm0_cntl        = 'd0         ;
    std__pe40__lane25_strm0_data        = 'h1234_5678 ;
    std__pe40__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe40__lane25_strm1_cntl        = 'd0         ;
    std__pe40__lane25_strm1_data        = 'h1234_5678 ;
    std__pe40__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe40__lane26_strm0_cntl        = 'd0         ;
    std__pe40__lane26_strm0_data        = 'h1234_5678 ;
    std__pe40__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe40__lane26_strm1_cntl        = 'd0         ;
    std__pe40__lane26_strm1_data        = 'h1234_5678 ;
    std__pe40__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe40__lane27_strm0_cntl        = 'd0         ;
    std__pe40__lane27_strm0_data        = 'h1234_5678 ;
    std__pe40__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe40__lane27_strm1_cntl        = 'd0         ;
    std__pe40__lane27_strm1_data        = 'h1234_5678 ;
    std__pe40__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe40__lane28_strm0_cntl        = 'd0         ;
    std__pe40__lane28_strm0_data        = 'h1234_5678 ;
    std__pe40__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe40__lane28_strm1_cntl        = 'd0         ;
    std__pe40__lane28_strm1_data        = 'h1234_5678 ;
    std__pe40__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe40__lane29_strm0_cntl        = 'd0         ;
    std__pe40__lane29_strm0_data        = 'h1234_5678 ;
    std__pe40__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe40__lane29_strm1_cntl        = 'd0         ;
    std__pe40__lane29_strm1_data        = 'h1234_5678 ;
    std__pe40__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe40__lane30_strm0_cntl        = 'd0         ;
    std__pe40__lane30_strm0_data        = 'h1234_5678 ;
    std__pe40__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe40__lane30_strm1_cntl        = 'd0         ;
    std__pe40__lane30_strm1_data        = 'h1234_5678 ;
    std__pe40__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe40__lane31_strm0_cntl        = 'd0         ;
    std__pe40__lane31_strm0_data        = 'h1234_5678 ;
    std__pe40__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe40__lane31_strm1_cntl        = 'd0         ;
    std__pe40__lane31_strm1_data        = 'h1234_5678 ;
    std__pe40__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe41__lane0_strm0_cntl        = 'd0         ;
    std__pe41__lane0_strm0_data        = 'h1234_5678 ;
    std__pe41__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe41__lane0_strm1_cntl        = 'd0         ;
    std__pe41__lane0_strm1_data        = 'h1234_5678 ;
    std__pe41__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe41__lane1_strm0_cntl        = 'd0         ;
    std__pe41__lane1_strm0_data        = 'h1234_5678 ;
    std__pe41__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe41__lane1_strm1_cntl        = 'd0         ;
    std__pe41__lane1_strm1_data        = 'h1234_5678 ;
    std__pe41__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe41__lane2_strm0_cntl        = 'd0         ;
    std__pe41__lane2_strm0_data        = 'h1234_5678 ;
    std__pe41__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe41__lane2_strm1_cntl        = 'd0         ;
    std__pe41__lane2_strm1_data        = 'h1234_5678 ;
    std__pe41__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe41__lane3_strm0_cntl        = 'd0         ;
    std__pe41__lane3_strm0_data        = 'h1234_5678 ;
    std__pe41__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe41__lane3_strm1_cntl        = 'd0         ;
    std__pe41__lane3_strm1_data        = 'h1234_5678 ;
    std__pe41__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe41__lane4_strm0_cntl        = 'd0         ;
    std__pe41__lane4_strm0_data        = 'h1234_5678 ;
    std__pe41__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe41__lane4_strm1_cntl        = 'd0         ;
    std__pe41__lane4_strm1_data        = 'h1234_5678 ;
    std__pe41__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe41__lane5_strm0_cntl        = 'd0         ;
    std__pe41__lane5_strm0_data        = 'h1234_5678 ;
    std__pe41__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe41__lane5_strm1_cntl        = 'd0         ;
    std__pe41__lane5_strm1_data        = 'h1234_5678 ;
    std__pe41__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe41__lane6_strm0_cntl        = 'd0         ;
    std__pe41__lane6_strm0_data        = 'h1234_5678 ;
    std__pe41__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe41__lane6_strm1_cntl        = 'd0         ;
    std__pe41__lane6_strm1_data        = 'h1234_5678 ;
    std__pe41__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe41__lane7_strm0_cntl        = 'd0         ;
    std__pe41__lane7_strm0_data        = 'h1234_5678 ;
    std__pe41__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe41__lane7_strm1_cntl        = 'd0         ;
    std__pe41__lane7_strm1_data        = 'h1234_5678 ;
    std__pe41__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe41__lane8_strm0_cntl        = 'd0         ;
    std__pe41__lane8_strm0_data        = 'h1234_5678 ;
    std__pe41__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe41__lane8_strm1_cntl        = 'd0         ;
    std__pe41__lane8_strm1_data        = 'h1234_5678 ;
    std__pe41__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe41__lane9_strm0_cntl        = 'd0         ;
    std__pe41__lane9_strm0_data        = 'h1234_5678 ;
    std__pe41__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe41__lane9_strm1_cntl        = 'd0         ;
    std__pe41__lane9_strm1_data        = 'h1234_5678 ;
    std__pe41__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe41__lane10_strm0_cntl        = 'd0         ;
    std__pe41__lane10_strm0_data        = 'h1234_5678 ;
    std__pe41__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe41__lane10_strm1_cntl        = 'd0         ;
    std__pe41__lane10_strm1_data        = 'h1234_5678 ;
    std__pe41__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe41__lane11_strm0_cntl        = 'd0         ;
    std__pe41__lane11_strm0_data        = 'h1234_5678 ;
    std__pe41__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe41__lane11_strm1_cntl        = 'd0         ;
    std__pe41__lane11_strm1_data        = 'h1234_5678 ;
    std__pe41__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe41__lane12_strm0_cntl        = 'd0         ;
    std__pe41__lane12_strm0_data        = 'h1234_5678 ;
    std__pe41__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe41__lane12_strm1_cntl        = 'd0         ;
    std__pe41__lane12_strm1_data        = 'h1234_5678 ;
    std__pe41__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe41__lane13_strm0_cntl        = 'd0         ;
    std__pe41__lane13_strm0_data        = 'h1234_5678 ;
    std__pe41__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe41__lane13_strm1_cntl        = 'd0         ;
    std__pe41__lane13_strm1_data        = 'h1234_5678 ;
    std__pe41__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe41__lane14_strm0_cntl        = 'd0         ;
    std__pe41__lane14_strm0_data        = 'h1234_5678 ;
    std__pe41__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe41__lane14_strm1_cntl        = 'd0         ;
    std__pe41__lane14_strm1_data        = 'h1234_5678 ;
    std__pe41__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe41__lane15_strm0_cntl        = 'd0         ;
    std__pe41__lane15_strm0_data        = 'h1234_5678 ;
    std__pe41__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe41__lane15_strm1_cntl        = 'd0         ;
    std__pe41__lane15_strm1_data        = 'h1234_5678 ;
    std__pe41__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe41__lane16_strm0_cntl        = 'd0         ;
    std__pe41__lane16_strm0_data        = 'h1234_5678 ;
    std__pe41__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe41__lane16_strm1_cntl        = 'd0         ;
    std__pe41__lane16_strm1_data        = 'h1234_5678 ;
    std__pe41__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe41__lane17_strm0_cntl        = 'd0         ;
    std__pe41__lane17_strm0_data        = 'h1234_5678 ;
    std__pe41__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe41__lane17_strm1_cntl        = 'd0         ;
    std__pe41__lane17_strm1_data        = 'h1234_5678 ;
    std__pe41__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe41__lane18_strm0_cntl        = 'd0         ;
    std__pe41__lane18_strm0_data        = 'h1234_5678 ;
    std__pe41__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe41__lane18_strm1_cntl        = 'd0         ;
    std__pe41__lane18_strm1_data        = 'h1234_5678 ;
    std__pe41__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe41__lane19_strm0_cntl        = 'd0         ;
    std__pe41__lane19_strm0_data        = 'h1234_5678 ;
    std__pe41__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe41__lane19_strm1_cntl        = 'd0         ;
    std__pe41__lane19_strm1_data        = 'h1234_5678 ;
    std__pe41__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe41__lane20_strm0_cntl        = 'd0         ;
    std__pe41__lane20_strm0_data        = 'h1234_5678 ;
    std__pe41__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe41__lane20_strm1_cntl        = 'd0         ;
    std__pe41__lane20_strm1_data        = 'h1234_5678 ;
    std__pe41__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe41__lane21_strm0_cntl        = 'd0         ;
    std__pe41__lane21_strm0_data        = 'h1234_5678 ;
    std__pe41__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe41__lane21_strm1_cntl        = 'd0         ;
    std__pe41__lane21_strm1_data        = 'h1234_5678 ;
    std__pe41__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe41__lane22_strm0_cntl        = 'd0         ;
    std__pe41__lane22_strm0_data        = 'h1234_5678 ;
    std__pe41__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe41__lane22_strm1_cntl        = 'd0         ;
    std__pe41__lane22_strm1_data        = 'h1234_5678 ;
    std__pe41__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe41__lane23_strm0_cntl        = 'd0         ;
    std__pe41__lane23_strm0_data        = 'h1234_5678 ;
    std__pe41__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe41__lane23_strm1_cntl        = 'd0         ;
    std__pe41__lane23_strm1_data        = 'h1234_5678 ;
    std__pe41__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe41__lane24_strm0_cntl        = 'd0         ;
    std__pe41__lane24_strm0_data        = 'h1234_5678 ;
    std__pe41__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe41__lane24_strm1_cntl        = 'd0         ;
    std__pe41__lane24_strm1_data        = 'h1234_5678 ;
    std__pe41__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe41__lane25_strm0_cntl        = 'd0         ;
    std__pe41__lane25_strm0_data        = 'h1234_5678 ;
    std__pe41__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe41__lane25_strm1_cntl        = 'd0         ;
    std__pe41__lane25_strm1_data        = 'h1234_5678 ;
    std__pe41__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe41__lane26_strm0_cntl        = 'd0         ;
    std__pe41__lane26_strm0_data        = 'h1234_5678 ;
    std__pe41__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe41__lane26_strm1_cntl        = 'd0         ;
    std__pe41__lane26_strm1_data        = 'h1234_5678 ;
    std__pe41__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe41__lane27_strm0_cntl        = 'd0         ;
    std__pe41__lane27_strm0_data        = 'h1234_5678 ;
    std__pe41__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe41__lane27_strm1_cntl        = 'd0         ;
    std__pe41__lane27_strm1_data        = 'h1234_5678 ;
    std__pe41__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe41__lane28_strm0_cntl        = 'd0         ;
    std__pe41__lane28_strm0_data        = 'h1234_5678 ;
    std__pe41__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe41__lane28_strm1_cntl        = 'd0         ;
    std__pe41__lane28_strm1_data        = 'h1234_5678 ;
    std__pe41__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe41__lane29_strm0_cntl        = 'd0         ;
    std__pe41__lane29_strm0_data        = 'h1234_5678 ;
    std__pe41__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe41__lane29_strm1_cntl        = 'd0         ;
    std__pe41__lane29_strm1_data        = 'h1234_5678 ;
    std__pe41__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe41__lane30_strm0_cntl        = 'd0         ;
    std__pe41__lane30_strm0_data        = 'h1234_5678 ;
    std__pe41__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe41__lane30_strm1_cntl        = 'd0         ;
    std__pe41__lane30_strm1_data        = 'h1234_5678 ;
    std__pe41__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe41__lane31_strm0_cntl        = 'd0         ;
    std__pe41__lane31_strm0_data        = 'h1234_5678 ;
    std__pe41__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe41__lane31_strm1_cntl        = 'd0         ;
    std__pe41__lane31_strm1_data        = 'h1234_5678 ;
    std__pe41__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe42__lane0_strm0_cntl        = 'd0         ;
    std__pe42__lane0_strm0_data        = 'h1234_5678 ;
    std__pe42__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe42__lane0_strm1_cntl        = 'd0         ;
    std__pe42__lane0_strm1_data        = 'h1234_5678 ;
    std__pe42__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe42__lane1_strm0_cntl        = 'd0         ;
    std__pe42__lane1_strm0_data        = 'h1234_5678 ;
    std__pe42__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe42__lane1_strm1_cntl        = 'd0         ;
    std__pe42__lane1_strm1_data        = 'h1234_5678 ;
    std__pe42__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe42__lane2_strm0_cntl        = 'd0         ;
    std__pe42__lane2_strm0_data        = 'h1234_5678 ;
    std__pe42__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe42__lane2_strm1_cntl        = 'd0         ;
    std__pe42__lane2_strm1_data        = 'h1234_5678 ;
    std__pe42__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe42__lane3_strm0_cntl        = 'd0         ;
    std__pe42__lane3_strm0_data        = 'h1234_5678 ;
    std__pe42__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe42__lane3_strm1_cntl        = 'd0         ;
    std__pe42__lane3_strm1_data        = 'h1234_5678 ;
    std__pe42__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe42__lane4_strm0_cntl        = 'd0         ;
    std__pe42__lane4_strm0_data        = 'h1234_5678 ;
    std__pe42__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe42__lane4_strm1_cntl        = 'd0         ;
    std__pe42__lane4_strm1_data        = 'h1234_5678 ;
    std__pe42__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe42__lane5_strm0_cntl        = 'd0         ;
    std__pe42__lane5_strm0_data        = 'h1234_5678 ;
    std__pe42__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe42__lane5_strm1_cntl        = 'd0         ;
    std__pe42__lane5_strm1_data        = 'h1234_5678 ;
    std__pe42__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe42__lane6_strm0_cntl        = 'd0         ;
    std__pe42__lane6_strm0_data        = 'h1234_5678 ;
    std__pe42__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe42__lane6_strm1_cntl        = 'd0         ;
    std__pe42__lane6_strm1_data        = 'h1234_5678 ;
    std__pe42__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe42__lane7_strm0_cntl        = 'd0         ;
    std__pe42__lane7_strm0_data        = 'h1234_5678 ;
    std__pe42__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe42__lane7_strm1_cntl        = 'd0         ;
    std__pe42__lane7_strm1_data        = 'h1234_5678 ;
    std__pe42__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe42__lane8_strm0_cntl        = 'd0         ;
    std__pe42__lane8_strm0_data        = 'h1234_5678 ;
    std__pe42__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe42__lane8_strm1_cntl        = 'd0         ;
    std__pe42__lane8_strm1_data        = 'h1234_5678 ;
    std__pe42__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe42__lane9_strm0_cntl        = 'd0         ;
    std__pe42__lane9_strm0_data        = 'h1234_5678 ;
    std__pe42__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe42__lane9_strm1_cntl        = 'd0         ;
    std__pe42__lane9_strm1_data        = 'h1234_5678 ;
    std__pe42__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe42__lane10_strm0_cntl        = 'd0         ;
    std__pe42__lane10_strm0_data        = 'h1234_5678 ;
    std__pe42__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe42__lane10_strm1_cntl        = 'd0         ;
    std__pe42__lane10_strm1_data        = 'h1234_5678 ;
    std__pe42__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe42__lane11_strm0_cntl        = 'd0         ;
    std__pe42__lane11_strm0_data        = 'h1234_5678 ;
    std__pe42__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe42__lane11_strm1_cntl        = 'd0         ;
    std__pe42__lane11_strm1_data        = 'h1234_5678 ;
    std__pe42__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe42__lane12_strm0_cntl        = 'd0         ;
    std__pe42__lane12_strm0_data        = 'h1234_5678 ;
    std__pe42__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe42__lane12_strm1_cntl        = 'd0         ;
    std__pe42__lane12_strm1_data        = 'h1234_5678 ;
    std__pe42__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe42__lane13_strm0_cntl        = 'd0         ;
    std__pe42__lane13_strm0_data        = 'h1234_5678 ;
    std__pe42__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe42__lane13_strm1_cntl        = 'd0         ;
    std__pe42__lane13_strm1_data        = 'h1234_5678 ;
    std__pe42__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe42__lane14_strm0_cntl        = 'd0         ;
    std__pe42__lane14_strm0_data        = 'h1234_5678 ;
    std__pe42__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe42__lane14_strm1_cntl        = 'd0         ;
    std__pe42__lane14_strm1_data        = 'h1234_5678 ;
    std__pe42__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe42__lane15_strm0_cntl        = 'd0         ;
    std__pe42__lane15_strm0_data        = 'h1234_5678 ;
    std__pe42__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe42__lane15_strm1_cntl        = 'd0         ;
    std__pe42__lane15_strm1_data        = 'h1234_5678 ;
    std__pe42__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe42__lane16_strm0_cntl        = 'd0         ;
    std__pe42__lane16_strm0_data        = 'h1234_5678 ;
    std__pe42__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe42__lane16_strm1_cntl        = 'd0         ;
    std__pe42__lane16_strm1_data        = 'h1234_5678 ;
    std__pe42__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe42__lane17_strm0_cntl        = 'd0         ;
    std__pe42__lane17_strm0_data        = 'h1234_5678 ;
    std__pe42__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe42__lane17_strm1_cntl        = 'd0         ;
    std__pe42__lane17_strm1_data        = 'h1234_5678 ;
    std__pe42__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe42__lane18_strm0_cntl        = 'd0         ;
    std__pe42__lane18_strm0_data        = 'h1234_5678 ;
    std__pe42__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe42__lane18_strm1_cntl        = 'd0         ;
    std__pe42__lane18_strm1_data        = 'h1234_5678 ;
    std__pe42__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe42__lane19_strm0_cntl        = 'd0         ;
    std__pe42__lane19_strm0_data        = 'h1234_5678 ;
    std__pe42__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe42__lane19_strm1_cntl        = 'd0         ;
    std__pe42__lane19_strm1_data        = 'h1234_5678 ;
    std__pe42__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe42__lane20_strm0_cntl        = 'd0         ;
    std__pe42__lane20_strm0_data        = 'h1234_5678 ;
    std__pe42__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe42__lane20_strm1_cntl        = 'd0         ;
    std__pe42__lane20_strm1_data        = 'h1234_5678 ;
    std__pe42__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe42__lane21_strm0_cntl        = 'd0         ;
    std__pe42__lane21_strm0_data        = 'h1234_5678 ;
    std__pe42__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe42__lane21_strm1_cntl        = 'd0         ;
    std__pe42__lane21_strm1_data        = 'h1234_5678 ;
    std__pe42__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe42__lane22_strm0_cntl        = 'd0         ;
    std__pe42__lane22_strm0_data        = 'h1234_5678 ;
    std__pe42__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe42__lane22_strm1_cntl        = 'd0         ;
    std__pe42__lane22_strm1_data        = 'h1234_5678 ;
    std__pe42__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe42__lane23_strm0_cntl        = 'd0         ;
    std__pe42__lane23_strm0_data        = 'h1234_5678 ;
    std__pe42__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe42__lane23_strm1_cntl        = 'd0         ;
    std__pe42__lane23_strm1_data        = 'h1234_5678 ;
    std__pe42__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe42__lane24_strm0_cntl        = 'd0         ;
    std__pe42__lane24_strm0_data        = 'h1234_5678 ;
    std__pe42__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe42__lane24_strm1_cntl        = 'd0         ;
    std__pe42__lane24_strm1_data        = 'h1234_5678 ;
    std__pe42__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe42__lane25_strm0_cntl        = 'd0         ;
    std__pe42__lane25_strm0_data        = 'h1234_5678 ;
    std__pe42__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe42__lane25_strm1_cntl        = 'd0         ;
    std__pe42__lane25_strm1_data        = 'h1234_5678 ;
    std__pe42__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe42__lane26_strm0_cntl        = 'd0         ;
    std__pe42__lane26_strm0_data        = 'h1234_5678 ;
    std__pe42__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe42__lane26_strm1_cntl        = 'd0         ;
    std__pe42__lane26_strm1_data        = 'h1234_5678 ;
    std__pe42__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe42__lane27_strm0_cntl        = 'd0         ;
    std__pe42__lane27_strm0_data        = 'h1234_5678 ;
    std__pe42__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe42__lane27_strm1_cntl        = 'd0         ;
    std__pe42__lane27_strm1_data        = 'h1234_5678 ;
    std__pe42__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe42__lane28_strm0_cntl        = 'd0         ;
    std__pe42__lane28_strm0_data        = 'h1234_5678 ;
    std__pe42__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe42__lane28_strm1_cntl        = 'd0         ;
    std__pe42__lane28_strm1_data        = 'h1234_5678 ;
    std__pe42__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe42__lane29_strm0_cntl        = 'd0         ;
    std__pe42__lane29_strm0_data        = 'h1234_5678 ;
    std__pe42__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe42__lane29_strm1_cntl        = 'd0         ;
    std__pe42__lane29_strm1_data        = 'h1234_5678 ;
    std__pe42__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe42__lane30_strm0_cntl        = 'd0         ;
    std__pe42__lane30_strm0_data        = 'h1234_5678 ;
    std__pe42__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe42__lane30_strm1_cntl        = 'd0         ;
    std__pe42__lane30_strm1_data        = 'h1234_5678 ;
    std__pe42__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe42__lane31_strm0_cntl        = 'd0         ;
    std__pe42__lane31_strm0_data        = 'h1234_5678 ;
    std__pe42__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe42__lane31_strm1_cntl        = 'd0         ;
    std__pe42__lane31_strm1_data        = 'h1234_5678 ;
    std__pe42__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe43__lane0_strm0_cntl        = 'd0         ;
    std__pe43__lane0_strm0_data        = 'h1234_5678 ;
    std__pe43__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe43__lane0_strm1_cntl        = 'd0         ;
    std__pe43__lane0_strm1_data        = 'h1234_5678 ;
    std__pe43__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe43__lane1_strm0_cntl        = 'd0         ;
    std__pe43__lane1_strm0_data        = 'h1234_5678 ;
    std__pe43__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe43__lane1_strm1_cntl        = 'd0         ;
    std__pe43__lane1_strm1_data        = 'h1234_5678 ;
    std__pe43__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe43__lane2_strm0_cntl        = 'd0         ;
    std__pe43__lane2_strm0_data        = 'h1234_5678 ;
    std__pe43__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe43__lane2_strm1_cntl        = 'd0         ;
    std__pe43__lane2_strm1_data        = 'h1234_5678 ;
    std__pe43__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe43__lane3_strm0_cntl        = 'd0         ;
    std__pe43__lane3_strm0_data        = 'h1234_5678 ;
    std__pe43__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe43__lane3_strm1_cntl        = 'd0         ;
    std__pe43__lane3_strm1_data        = 'h1234_5678 ;
    std__pe43__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe43__lane4_strm0_cntl        = 'd0         ;
    std__pe43__lane4_strm0_data        = 'h1234_5678 ;
    std__pe43__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe43__lane4_strm1_cntl        = 'd0         ;
    std__pe43__lane4_strm1_data        = 'h1234_5678 ;
    std__pe43__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe43__lane5_strm0_cntl        = 'd0         ;
    std__pe43__lane5_strm0_data        = 'h1234_5678 ;
    std__pe43__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe43__lane5_strm1_cntl        = 'd0         ;
    std__pe43__lane5_strm1_data        = 'h1234_5678 ;
    std__pe43__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe43__lane6_strm0_cntl        = 'd0         ;
    std__pe43__lane6_strm0_data        = 'h1234_5678 ;
    std__pe43__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe43__lane6_strm1_cntl        = 'd0         ;
    std__pe43__lane6_strm1_data        = 'h1234_5678 ;
    std__pe43__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe43__lane7_strm0_cntl        = 'd0         ;
    std__pe43__lane7_strm0_data        = 'h1234_5678 ;
    std__pe43__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe43__lane7_strm1_cntl        = 'd0         ;
    std__pe43__lane7_strm1_data        = 'h1234_5678 ;
    std__pe43__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe43__lane8_strm0_cntl        = 'd0         ;
    std__pe43__lane8_strm0_data        = 'h1234_5678 ;
    std__pe43__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe43__lane8_strm1_cntl        = 'd0         ;
    std__pe43__lane8_strm1_data        = 'h1234_5678 ;
    std__pe43__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe43__lane9_strm0_cntl        = 'd0         ;
    std__pe43__lane9_strm0_data        = 'h1234_5678 ;
    std__pe43__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe43__lane9_strm1_cntl        = 'd0         ;
    std__pe43__lane9_strm1_data        = 'h1234_5678 ;
    std__pe43__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe43__lane10_strm0_cntl        = 'd0         ;
    std__pe43__lane10_strm0_data        = 'h1234_5678 ;
    std__pe43__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe43__lane10_strm1_cntl        = 'd0         ;
    std__pe43__lane10_strm1_data        = 'h1234_5678 ;
    std__pe43__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe43__lane11_strm0_cntl        = 'd0         ;
    std__pe43__lane11_strm0_data        = 'h1234_5678 ;
    std__pe43__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe43__lane11_strm1_cntl        = 'd0         ;
    std__pe43__lane11_strm1_data        = 'h1234_5678 ;
    std__pe43__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe43__lane12_strm0_cntl        = 'd0         ;
    std__pe43__lane12_strm0_data        = 'h1234_5678 ;
    std__pe43__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe43__lane12_strm1_cntl        = 'd0         ;
    std__pe43__lane12_strm1_data        = 'h1234_5678 ;
    std__pe43__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe43__lane13_strm0_cntl        = 'd0         ;
    std__pe43__lane13_strm0_data        = 'h1234_5678 ;
    std__pe43__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe43__lane13_strm1_cntl        = 'd0         ;
    std__pe43__lane13_strm1_data        = 'h1234_5678 ;
    std__pe43__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe43__lane14_strm0_cntl        = 'd0         ;
    std__pe43__lane14_strm0_data        = 'h1234_5678 ;
    std__pe43__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe43__lane14_strm1_cntl        = 'd0         ;
    std__pe43__lane14_strm1_data        = 'h1234_5678 ;
    std__pe43__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe43__lane15_strm0_cntl        = 'd0         ;
    std__pe43__lane15_strm0_data        = 'h1234_5678 ;
    std__pe43__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe43__lane15_strm1_cntl        = 'd0         ;
    std__pe43__lane15_strm1_data        = 'h1234_5678 ;
    std__pe43__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe43__lane16_strm0_cntl        = 'd0         ;
    std__pe43__lane16_strm0_data        = 'h1234_5678 ;
    std__pe43__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe43__lane16_strm1_cntl        = 'd0         ;
    std__pe43__lane16_strm1_data        = 'h1234_5678 ;
    std__pe43__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe43__lane17_strm0_cntl        = 'd0         ;
    std__pe43__lane17_strm0_data        = 'h1234_5678 ;
    std__pe43__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe43__lane17_strm1_cntl        = 'd0         ;
    std__pe43__lane17_strm1_data        = 'h1234_5678 ;
    std__pe43__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe43__lane18_strm0_cntl        = 'd0         ;
    std__pe43__lane18_strm0_data        = 'h1234_5678 ;
    std__pe43__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe43__lane18_strm1_cntl        = 'd0         ;
    std__pe43__lane18_strm1_data        = 'h1234_5678 ;
    std__pe43__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe43__lane19_strm0_cntl        = 'd0         ;
    std__pe43__lane19_strm0_data        = 'h1234_5678 ;
    std__pe43__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe43__lane19_strm1_cntl        = 'd0         ;
    std__pe43__lane19_strm1_data        = 'h1234_5678 ;
    std__pe43__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe43__lane20_strm0_cntl        = 'd0         ;
    std__pe43__lane20_strm0_data        = 'h1234_5678 ;
    std__pe43__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe43__lane20_strm1_cntl        = 'd0         ;
    std__pe43__lane20_strm1_data        = 'h1234_5678 ;
    std__pe43__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe43__lane21_strm0_cntl        = 'd0         ;
    std__pe43__lane21_strm0_data        = 'h1234_5678 ;
    std__pe43__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe43__lane21_strm1_cntl        = 'd0         ;
    std__pe43__lane21_strm1_data        = 'h1234_5678 ;
    std__pe43__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe43__lane22_strm0_cntl        = 'd0         ;
    std__pe43__lane22_strm0_data        = 'h1234_5678 ;
    std__pe43__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe43__lane22_strm1_cntl        = 'd0         ;
    std__pe43__lane22_strm1_data        = 'h1234_5678 ;
    std__pe43__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe43__lane23_strm0_cntl        = 'd0         ;
    std__pe43__lane23_strm0_data        = 'h1234_5678 ;
    std__pe43__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe43__lane23_strm1_cntl        = 'd0         ;
    std__pe43__lane23_strm1_data        = 'h1234_5678 ;
    std__pe43__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe43__lane24_strm0_cntl        = 'd0         ;
    std__pe43__lane24_strm0_data        = 'h1234_5678 ;
    std__pe43__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe43__lane24_strm1_cntl        = 'd0         ;
    std__pe43__lane24_strm1_data        = 'h1234_5678 ;
    std__pe43__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe43__lane25_strm0_cntl        = 'd0         ;
    std__pe43__lane25_strm0_data        = 'h1234_5678 ;
    std__pe43__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe43__lane25_strm1_cntl        = 'd0         ;
    std__pe43__lane25_strm1_data        = 'h1234_5678 ;
    std__pe43__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe43__lane26_strm0_cntl        = 'd0         ;
    std__pe43__lane26_strm0_data        = 'h1234_5678 ;
    std__pe43__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe43__lane26_strm1_cntl        = 'd0         ;
    std__pe43__lane26_strm1_data        = 'h1234_5678 ;
    std__pe43__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe43__lane27_strm0_cntl        = 'd0         ;
    std__pe43__lane27_strm0_data        = 'h1234_5678 ;
    std__pe43__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe43__lane27_strm1_cntl        = 'd0         ;
    std__pe43__lane27_strm1_data        = 'h1234_5678 ;
    std__pe43__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe43__lane28_strm0_cntl        = 'd0         ;
    std__pe43__lane28_strm0_data        = 'h1234_5678 ;
    std__pe43__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe43__lane28_strm1_cntl        = 'd0         ;
    std__pe43__lane28_strm1_data        = 'h1234_5678 ;
    std__pe43__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe43__lane29_strm0_cntl        = 'd0         ;
    std__pe43__lane29_strm0_data        = 'h1234_5678 ;
    std__pe43__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe43__lane29_strm1_cntl        = 'd0         ;
    std__pe43__lane29_strm1_data        = 'h1234_5678 ;
    std__pe43__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe43__lane30_strm0_cntl        = 'd0         ;
    std__pe43__lane30_strm0_data        = 'h1234_5678 ;
    std__pe43__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe43__lane30_strm1_cntl        = 'd0         ;
    std__pe43__lane30_strm1_data        = 'h1234_5678 ;
    std__pe43__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe43__lane31_strm0_cntl        = 'd0         ;
    std__pe43__lane31_strm0_data        = 'h1234_5678 ;
    std__pe43__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe43__lane31_strm1_cntl        = 'd0         ;
    std__pe43__lane31_strm1_data        = 'h1234_5678 ;
    std__pe43__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe44__lane0_strm0_cntl        = 'd0         ;
    std__pe44__lane0_strm0_data        = 'h1234_5678 ;
    std__pe44__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe44__lane0_strm1_cntl        = 'd0         ;
    std__pe44__lane0_strm1_data        = 'h1234_5678 ;
    std__pe44__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe44__lane1_strm0_cntl        = 'd0         ;
    std__pe44__lane1_strm0_data        = 'h1234_5678 ;
    std__pe44__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe44__lane1_strm1_cntl        = 'd0         ;
    std__pe44__lane1_strm1_data        = 'h1234_5678 ;
    std__pe44__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe44__lane2_strm0_cntl        = 'd0         ;
    std__pe44__lane2_strm0_data        = 'h1234_5678 ;
    std__pe44__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe44__lane2_strm1_cntl        = 'd0         ;
    std__pe44__lane2_strm1_data        = 'h1234_5678 ;
    std__pe44__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe44__lane3_strm0_cntl        = 'd0         ;
    std__pe44__lane3_strm0_data        = 'h1234_5678 ;
    std__pe44__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe44__lane3_strm1_cntl        = 'd0         ;
    std__pe44__lane3_strm1_data        = 'h1234_5678 ;
    std__pe44__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe44__lane4_strm0_cntl        = 'd0         ;
    std__pe44__lane4_strm0_data        = 'h1234_5678 ;
    std__pe44__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe44__lane4_strm1_cntl        = 'd0         ;
    std__pe44__lane4_strm1_data        = 'h1234_5678 ;
    std__pe44__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe44__lane5_strm0_cntl        = 'd0         ;
    std__pe44__lane5_strm0_data        = 'h1234_5678 ;
    std__pe44__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe44__lane5_strm1_cntl        = 'd0         ;
    std__pe44__lane5_strm1_data        = 'h1234_5678 ;
    std__pe44__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe44__lane6_strm0_cntl        = 'd0         ;
    std__pe44__lane6_strm0_data        = 'h1234_5678 ;
    std__pe44__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe44__lane6_strm1_cntl        = 'd0         ;
    std__pe44__lane6_strm1_data        = 'h1234_5678 ;
    std__pe44__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe44__lane7_strm0_cntl        = 'd0         ;
    std__pe44__lane7_strm0_data        = 'h1234_5678 ;
    std__pe44__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe44__lane7_strm1_cntl        = 'd0         ;
    std__pe44__lane7_strm1_data        = 'h1234_5678 ;
    std__pe44__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe44__lane8_strm0_cntl        = 'd0         ;
    std__pe44__lane8_strm0_data        = 'h1234_5678 ;
    std__pe44__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe44__lane8_strm1_cntl        = 'd0         ;
    std__pe44__lane8_strm1_data        = 'h1234_5678 ;
    std__pe44__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe44__lane9_strm0_cntl        = 'd0         ;
    std__pe44__lane9_strm0_data        = 'h1234_5678 ;
    std__pe44__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe44__lane9_strm1_cntl        = 'd0         ;
    std__pe44__lane9_strm1_data        = 'h1234_5678 ;
    std__pe44__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe44__lane10_strm0_cntl        = 'd0         ;
    std__pe44__lane10_strm0_data        = 'h1234_5678 ;
    std__pe44__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe44__lane10_strm1_cntl        = 'd0         ;
    std__pe44__lane10_strm1_data        = 'h1234_5678 ;
    std__pe44__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe44__lane11_strm0_cntl        = 'd0         ;
    std__pe44__lane11_strm0_data        = 'h1234_5678 ;
    std__pe44__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe44__lane11_strm1_cntl        = 'd0         ;
    std__pe44__lane11_strm1_data        = 'h1234_5678 ;
    std__pe44__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe44__lane12_strm0_cntl        = 'd0         ;
    std__pe44__lane12_strm0_data        = 'h1234_5678 ;
    std__pe44__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe44__lane12_strm1_cntl        = 'd0         ;
    std__pe44__lane12_strm1_data        = 'h1234_5678 ;
    std__pe44__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe44__lane13_strm0_cntl        = 'd0         ;
    std__pe44__lane13_strm0_data        = 'h1234_5678 ;
    std__pe44__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe44__lane13_strm1_cntl        = 'd0         ;
    std__pe44__lane13_strm1_data        = 'h1234_5678 ;
    std__pe44__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe44__lane14_strm0_cntl        = 'd0         ;
    std__pe44__lane14_strm0_data        = 'h1234_5678 ;
    std__pe44__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe44__lane14_strm1_cntl        = 'd0         ;
    std__pe44__lane14_strm1_data        = 'h1234_5678 ;
    std__pe44__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe44__lane15_strm0_cntl        = 'd0         ;
    std__pe44__lane15_strm0_data        = 'h1234_5678 ;
    std__pe44__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe44__lane15_strm1_cntl        = 'd0         ;
    std__pe44__lane15_strm1_data        = 'h1234_5678 ;
    std__pe44__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe44__lane16_strm0_cntl        = 'd0         ;
    std__pe44__lane16_strm0_data        = 'h1234_5678 ;
    std__pe44__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe44__lane16_strm1_cntl        = 'd0         ;
    std__pe44__lane16_strm1_data        = 'h1234_5678 ;
    std__pe44__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe44__lane17_strm0_cntl        = 'd0         ;
    std__pe44__lane17_strm0_data        = 'h1234_5678 ;
    std__pe44__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe44__lane17_strm1_cntl        = 'd0         ;
    std__pe44__lane17_strm1_data        = 'h1234_5678 ;
    std__pe44__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe44__lane18_strm0_cntl        = 'd0         ;
    std__pe44__lane18_strm0_data        = 'h1234_5678 ;
    std__pe44__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe44__lane18_strm1_cntl        = 'd0         ;
    std__pe44__lane18_strm1_data        = 'h1234_5678 ;
    std__pe44__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe44__lane19_strm0_cntl        = 'd0         ;
    std__pe44__lane19_strm0_data        = 'h1234_5678 ;
    std__pe44__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe44__lane19_strm1_cntl        = 'd0         ;
    std__pe44__lane19_strm1_data        = 'h1234_5678 ;
    std__pe44__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe44__lane20_strm0_cntl        = 'd0         ;
    std__pe44__lane20_strm0_data        = 'h1234_5678 ;
    std__pe44__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe44__lane20_strm1_cntl        = 'd0         ;
    std__pe44__lane20_strm1_data        = 'h1234_5678 ;
    std__pe44__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe44__lane21_strm0_cntl        = 'd0         ;
    std__pe44__lane21_strm0_data        = 'h1234_5678 ;
    std__pe44__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe44__lane21_strm1_cntl        = 'd0         ;
    std__pe44__lane21_strm1_data        = 'h1234_5678 ;
    std__pe44__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe44__lane22_strm0_cntl        = 'd0         ;
    std__pe44__lane22_strm0_data        = 'h1234_5678 ;
    std__pe44__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe44__lane22_strm1_cntl        = 'd0         ;
    std__pe44__lane22_strm1_data        = 'h1234_5678 ;
    std__pe44__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe44__lane23_strm0_cntl        = 'd0         ;
    std__pe44__lane23_strm0_data        = 'h1234_5678 ;
    std__pe44__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe44__lane23_strm1_cntl        = 'd0         ;
    std__pe44__lane23_strm1_data        = 'h1234_5678 ;
    std__pe44__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe44__lane24_strm0_cntl        = 'd0         ;
    std__pe44__lane24_strm0_data        = 'h1234_5678 ;
    std__pe44__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe44__lane24_strm1_cntl        = 'd0         ;
    std__pe44__lane24_strm1_data        = 'h1234_5678 ;
    std__pe44__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe44__lane25_strm0_cntl        = 'd0         ;
    std__pe44__lane25_strm0_data        = 'h1234_5678 ;
    std__pe44__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe44__lane25_strm1_cntl        = 'd0         ;
    std__pe44__lane25_strm1_data        = 'h1234_5678 ;
    std__pe44__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe44__lane26_strm0_cntl        = 'd0         ;
    std__pe44__lane26_strm0_data        = 'h1234_5678 ;
    std__pe44__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe44__lane26_strm1_cntl        = 'd0         ;
    std__pe44__lane26_strm1_data        = 'h1234_5678 ;
    std__pe44__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe44__lane27_strm0_cntl        = 'd0         ;
    std__pe44__lane27_strm0_data        = 'h1234_5678 ;
    std__pe44__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe44__lane27_strm1_cntl        = 'd0         ;
    std__pe44__lane27_strm1_data        = 'h1234_5678 ;
    std__pe44__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe44__lane28_strm0_cntl        = 'd0         ;
    std__pe44__lane28_strm0_data        = 'h1234_5678 ;
    std__pe44__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe44__lane28_strm1_cntl        = 'd0         ;
    std__pe44__lane28_strm1_data        = 'h1234_5678 ;
    std__pe44__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe44__lane29_strm0_cntl        = 'd0         ;
    std__pe44__lane29_strm0_data        = 'h1234_5678 ;
    std__pe44__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe44__lane29_strm1_cntl        = 'd0         ;
    std__pe44__lane29_strm1_data        = 'h1234_5678 ;
    std__pe44__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe44__lane30_strm0_cntl        = 'd0         ;
    std__pe44__lane30_strm0_data        = 'h1234_5678 ;
    std__pe44__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe44__lane30_strm1_cntl        = 'd0         ;
    std__pe44__lane30_strm1_data        = 'h1234_5678 ;
    std__pe44__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe44__lane31_strm0_cntl        = 'd0         ;
    std__pe44__lane31_strm0_data        = 'h1234_5678 ;
    std__pe44__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe44__lane31_strm1_cntl        = 'd0         ;
    std__pe44__lane31_strm1_data        = 'h1234_5678 ;
    std__pe44__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe45__lane0_strm0_cntl        = 'd0         ;
    std__pe45__lane0_strm0_data        = 'h1234_5678 ;
    std__pe45__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe45__lane0_strm1_cntl        = 'd0         ;
    std__pe45__lane0_strm1_data        = 'h1234_5678 ;
    std__pe45__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe45__lane1_strm0_cntl        = 'd0         ;
    std__pe45__lane1_strm0_data        = 'h1234_5678 ;
    std__pe45__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe45__lane1_strm1_cntl        = 'd0         ;
    std__pe45__lane1_strm1_data        = 'h1234_5678 ;
    std__pe45__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe45__lane2_strm0_cntl        = 'd0         ;
    std__pe45__lane2_strm0_data        = 'h1234_5678 ;
    std__pe45__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe45__lane2_strm1_cntl        = 'd0         ;
    std__pe45__lane2_strm1_data        = 'h1234_5678 ;
    std__pe45__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe45__lane3_strm0_cntl        = 'd0         ;
    std__pe45__lane3_strm0_data        = 'h1234_5678 ;
    std__pe45__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe45__lane3_strm1_cntl        = 'd0         ;
    std__pe45__lane3_strm1_data        = 'h1234_5678 ;
    std__pe45__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe45__lane4_strm0_cntl        = 'd0         ;
    std__pe45__lane4_strm0_data        = 'h1234_5678 ;
    std__pe45__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe45__lane4_strm1_cntl        = 'd0         ;
    std__pe45__lane4_strm1_data        = 'h1234_5678 ;
    std__pe45__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe45__lane5_strm0_cntl        = 'd0         ;
    std__pe45__lane5_strm0_data        = 'h1234_5678 ;
    std__pe45__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe45__lane5_strm1_cntl        = 'd0         ;
    std__pe45__lane5_strm1_data        = 'h1234_5678 ;
    std__pe45__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe45__lane6_strm0_cntl        = 'd0         ;
    std__pe45__lane6_strm0_data        = 'h1234_5678 ;
    std__pe45__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe45__lane6_strm1_cntl        = 'd0         ;
    std__pe45__lane6_strm1_data        = 'h1234_5678 ;
    std__pe45__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe45__lane7_strm0_cntl        = 'd0         ;
    std__pe45__lane7_strm0_data        = 'h1234_5678 ;
    std__pe45__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe45__lane7_strm1_cntl        = 'd0         ;
    std__pe45__lane7_strm1_data        = 'h1234_5678 ;
    std__pe45__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe45__lane8_strm0_cntl        = 'd0         ;
    std__pe45__lane8_strm0_data        = 'h1234_5678 ;
    std__pe45__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe45__lane8_strm1_cntl        = 'd0         ;
    std__pe45__lane8_strm1_data        = 'h1234_5678 ;
    std__pe45__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe45__lane9_strm0_cntl        = 'd0         ;
    std__pe45__lane9_strm0_data        = 'h1234_5678 ;
    std__pe45__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe45__lane9_strm1_cntl        = 'd0         ;
    std__pe45__lane9_strm1_data        = 'h1234_5678 ;
    std__pe45__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe45__lane10_strm0_cntl        = 'd0         ;
    std__pe45__lane10_strm0_data        = 'h1234_5678 ;
    std__pe45__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe45__lane10_strm1_cntl        = 'd0         ;
    std__pe45__lane10_strm1_data        = 'h1234_5678 ;
    std__pe45__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe45__lane11_strm0_cntl        = 'd0         ;
    std__pe45__lane11_strm0_data        = 'h1234_5678 ;
    std__pe45__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe45__lane11_strm1_cntl        = 'd0         ;
    std__pe45__lane11_strm1_data        = 'h1234_5678 ;
    std__pe45__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe45__lane12_strm0_cntl        = 'd0         ;
    std__pe45__lane12_strm0_data        = 'h1234_5678 ;
    std__pe45__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe45__lane12_strm1_cntl        = 'd0         ;
    std__pe45__lane12_strm1_data        = 'h1234_5678 ;
    std__pe45__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe45__lane13_strm0_cntl        = 'd0         ;
    std__pe45__lane13_strm0_data        = 'h1234_5678 ;
    std__pe45__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe45__lane13_strm1_cntl        = 'd0         ;
    std__pe45__lane13_strm1_data        = 'h1234_5678 ;
    std__pe45__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe45__lane14_strm0_cntl        = 'd0         ;
    std__pe45__lane14_strm0_data        = 'h1234_5678 ;
    std__pe45__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe45__lane14_strm1_cntl        = 'd0         ;
    std__pe45__lane14_strm1_data        = 'h1234_5678 ;
    std__pe45__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe45__lane15_strm0_cntl        = 'd0         ;
    std__pe45__lane15_strm0_data        = 'h1234_5678 ;
    std__pe45__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe45__lane15_strm1_cntl        = 'd0         ;
    std__pe45__lane15_strm1_data        = 'h1234_5678 ;
    std__pe45__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe45__lane16_strm0_cntl        = 'd0         ;
    std__pe45__lane16_strm0_data        = 'h1234_5678 ;
    std__pe45__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe45__lane16_strm1_cntl        = 'd0         ;
    std__pe45__lane16_strm1_data        = 'h1234_5678 ;
    std__pe45__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe45__lane17_strm0_cntl        = 'd0         ;
    std__pe45__lane17_strm0_data        = 'h1234_5678 ;
    std__pe45__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe45__lane17_strm1_cntl        = 'd0         ;
    std__pe45__lane17_strm1_data        = 'h1234_5678 ;
    std__pe45__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe45__lane18_strm0_cntl        = 'd0         ;
    std__pe45__lane18_strm0_data        = 'h1234_5678 ;
    std__pe45__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe45__lane18_strm1_cntl        = 'd0         ;
    std__pe45__lane18_strm1_data        = 'h1234_5678 ;
    std__pe45__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe45__lane19_strm0_cntl        = 'd0         ;
    std__pe45__lane19_strm0_data        = 'h1234_5678 ;
    std__pe45__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe45__lane19_strm1_cntl        = 'd0         ;
    std__pe45__lane19_strm1_data        = 'h1234_5678 ;
    std__pe45__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe45__lane20_strm0_cntl        = 'd0         ;
    std__pe45__lane20_strm0_data        = 'h1234_5678 ;
    std__pe45__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe45__lane20_strm1_cntl        = 'd0         ;
    std__pe45__lane20_strm1_data        = 'h1234_5678 ;
    std__pe45__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe45__lane21_strm0_cntl        = 'd0         ;
    std__pe45__lane21_strm0_data        = 'h1234_5678 ;
    std__pe45__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe45__lane21_strm1_cntl        = 'd0         ;
    std__pe45__lane21_strm1_data        = 'h1234_5678 ;
    std__pe45__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe45__lane22_strm0_cntl        = 'd0         ;
    std__pe45__lane22_strm0_data        = 'h1234_5678 ;
    std__pe45__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe45__lane22_strm1_cntl        = 'd0         ;
    std__pe45__lane22_strm1_data        = 'h1234_5678 ;
    std__pe45__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe45__lane23_strm0_cntl        = 'd0         ;
    std__pe45__lane23_strm0_data        = 'h1234_5678 ;
    std__pe45__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe45__lane23_strm1_cntl        = 'd0         ;
    std__pe45__lane23_strm1_data        = 'h1234_5678 ;
    std__pe45__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe45__lane24_strm0_cntl        = 'd0         ;
    std__pe45__lane24_strm0_data        = 'h1234_5678 ;
    std__pe45__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe45__lane24_strm1_cntl        = 'd0         ;
    std__pe45__lane24_strm1_data        = 'h1234_5678 ;
    std__pe45__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe45__lane25_strm0_cntl        = 'd0         ;
    std__pe45__lane25_strm0_data        = 'h1234_5678 ;
    std__pe45__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe45__lane25_strm1_cntl        = 'd0         ;
    std__pe45__lane25_strm1_data        = 'h1234_5678 ;
    std__pe45__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe45__lane26_strm0_cntl        = 'd0         ;
    std__pe45__lane26_strm0_data        = 'h1234_5678 ;
    std__pe45__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe45__lane26_strm1_cntl        = 'd0         ;
    std__pe45__lane26_strm1_data        = 'h1234_5678 ;
    std__pe45__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe45__lane27_strm0_cntl        = 'd0         ;
    std__pe45__lane27_strm0_data        = 'h1234_5678 ;
    std__pe45__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe45__lane27_strm1_cntl        = 'd0         ;
    std__pe45__lane27_strm1_data        = 'h1234_5678 ;
    std__pe45__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe45__lane28_strm0_cntl        = 'd0         ;
    std__pe45__lane28_strm0_data        = 'h1234_5678 ;
    std__pe45__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe45__lane28_strm1_cntl        = 'd0         ;
    std__pe45__lane28_strm1_data        = 'h1234_5678 ;
    std__pe45__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe45__lane29_strm0_cntl        = 'd0         ;
    std__pe45__lane29_strm0_data        = 'h1234_5678 ;
    std__pe45__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe45__lane29_strm1_cntl        = 'd0         ;
    std__pe45__lane29_strm1_data        = 'h1234_5678 ;
    std__pe45__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe45__lane30_strm0_cntl        = 'd0         ;
    std__pe45__lane30_strm0_data        = 'h1234_5678 ;
    std__pe45__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe45__lane30_strm1_cntl        = 'd0         ;
    std__pe45__lane30_strm1_data        = 'h1234_5678 ;
    std__pe45__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe45__lane31_strm0_cntl        = 'd0         ;
    std__pe45__lane31_strm0_data        = 'h1234_5678 ;
    std__pe45__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe45__lane31_strm1_cntl        = 'd0         ;
    std__pe45__lane31_strm1_data        = 'h1234_5678 ;
    std__pe45__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe46__lane0_strm0_cntl        = 'd0         ;
    std__pe46__lane0_strm0_data        = 'h1234_5678 ;
    std__pe46__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe46__lane0_strm1_cntl        = 'd0         ;
    std__pe46__lane0_strm1_data        = 'h1234_5678 ;
    std__pe46__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe46__lane1_strm0_cntl        = 'd0         ;
    std__pe46__lane1_strm0_data        = 'h1234_5678 ;
    std__pe46__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe46__lane1_strm1_cntl        = 'd0         ;
    std__pe46__lane1_strm1_data        = 'h1234_5678 ;
    std__pe46__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe46__lane2_strm0_cntl        = 'd0         ;
    std__pe46__lane2_strm0_data        = 'h1234_5678 ;
    std__pe46__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe46__lane2_strm1_cntl        = 'd0         ;
    std__pe46__lane2_strm1_data        = 'h1234_5678 ;
    std__pe46__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe46__lane3_strm0_cntl        = 'd0         ;
    std__pe46__lane3_strm0_data        = 'h1234_5678 ;
    std__pe46__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe46__lane3_strm1_cntl        = 'd0         ;
    std__pe46__lane3_strm1_data        = 'h1234_5678 ;
    std__pe46__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe46__lane4_strm0_cntl        = 'd0         ;
    std__pe46__lane4_strm0_data        = 'h1234_5678 ;
    std__pe46__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe46__lane4_strm1_cntl        = 'd0         ;
    std__pe46__lane4_strm1_data        = 'h1234_5678 ;
    std__pe46__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe46__lane5_strm0_cntl        = 'd0         ;
    std__pe46__lane5_strm0_data        = 'h1234_5678 ;
    std__pe46__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe46__lane5_strm1_cntl        = 'd0         ;
    std__pe46__lane5_strm1_data        = 'h1234_5678 ;
    std__pe46__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe46__lane6_strm0_cntl        = 'd0         ;
    std__pe46__lane6_strm0_data        = 'h1234_5678 ;
    std__pe46__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe46__lane6_strm1_cntl        = 'd0         ;
    std__pe46__lane6_strm1_data        = 'h1234_5678 ;
    std__pe46__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe46__lane7_strm0_cntl        = 'd0         ;
    std__pe46__lane7_strm0_data        = 'h1234_5678 ;
    std__pe46__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe46__lane7_strm1_cntl        = 'd0         ;
    std__pe46__lane7_strm1_data        = 'h1234_5678 ;
    std__pe46__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe46__lane8_strm0_cntl        = 'd0         ;
    std__pe46__lane8_strm0_data        = 'h1234_5678 ;
    std__pe46__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe46__lane8_strm1_cntl        = 'd0         ;
    std__pe46__lane8_strm1_data        = 'h1234_5678 ;
    std__pe46__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe46__lane9_strm0_cntl        = 'd0         ;
    std__pe46__lane9_strm0_data        = 'h1234_5678 ;
    std__pe46__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe46__lane9_strm1_cntl        = 'd0         ;
    std__pe46__lane9_strm1_data        = 'h1234_5678 ;
    std__pe46__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe46__lane10_strm0_cntl        = 'd0         ;
    std__pe46__lane10_strm0_data        = 'h1234_5678 ;
    std__pe46__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe46__lane10_strm1_cntl        = 'd0         ;
    std__pe46__lane10_strm1_data        = 'h1234_5678 ;
    std__pe46__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe46__lane11_strm0_cntl        = 'd0         ;
    std__pe46__lane11_strm0_data        = 'h1234_5678 ;
    std__pe46__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe46__lane11_strm1_cntl        = 'd0         ;
    std__pe46__lane11_strm1_data        = 'h1234_5678 ;
    std__pe46__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe46__lane12_strm0_cntl        = 'd0         ;
    std__pe46__lane12_strm0_data        = 'h1234_5678 ;
    std__pe46__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe46__lane12_strm1_cntl        = 'd0         ;
    std__pe46__lane12_strm1_data        = 'h1234_5678 ;
    std__pe46__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe46__lane13_strm0_cntl        = 'd0         ;
    std__pe46__lane13_strm0_data        = 'h1234_5678 ;
    std__pe46__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe46__lane13_strm1_cntl        = 'd0         ;
    std__pe46__lane13_strm1_data        = 'h1234_5678 ;
    std__pe46__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe46__lane14_strm0_cntl        = 'd0         ;
    std__pe46__lane14_strm0_data        = 'h1234_5678 ;
    std__pe46__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe46__lane14_strm1_cntl        = 'd0         ;
    std__pe46__lane14_strm1_data        = 'h1234_5678 ;
    std__pe46__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe46__lane15_strm0_cntl        = 'd0         ;
    std__pe46__lane15_strm0_data        = 'h1234_5678 ;
    std__pe46__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe46__lane15_strm1_cntl        = 'd0         ;
    std__pe46__lane15_strm1_data        = 'h1234_5678 ;
    std__pe46__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe46__lane16_strm0_cntl        = 'd0         ;
    std__pe46__lane16_strm0_data        = 'h1234_5678 ;
    std__pe46__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe46__lane16_strm1_cntl        = 'd0         ;
    std__pe46__lane16_strm1_data        = 'h1234_5678 ;
    std__pe46__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe46__lane17_strm0_cntl        = 'd0         ;
    std__pe46__lane17_strm0_data        = 'h1234_5678 ;
    std__pe46__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe46__lane17_strm1_cntl        = 'd0         ;
    std__pe46__lane17_strm1_data        = 'h1234_5678 ;
    std__pe46__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe46__lane18_strm0_cntl        = 'd0         ;
    std__pe46__lane18_strm0_data        = 'h1234_5678 ;
    std__pe46__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe46__lane18_strm1_cntl        = 'd0         ;
    std__pe46__lane18_strm1_data        = 'h1234_5678 ;
    std__pe46__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe46__lane19_strm0_cntl        = 'd0         ;
    std__pe46__lane19_strm0_data        = 'h1234_5678 ;
    std__pe46__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe46__lane19_strm1_cntl        = 'd0         ;
    std__pe46__lane19_strm1_data        = 'h1234_5678 ;
    std__pe46__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe46__lane20_strm0_cntl        = 'd0         ;
    std__pe46__lane20_strm0_data        = 'h1234_5678 ;
    std__pe46__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe46__lane20_strm1_cntl        = 'd0         ;
    std__pe46__lane20_strm1_data        = 'h1234_5678 ;
    std__pe46__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe46__lane21_strm0_cntl        = 'd0         ;
    std__pe46__lane21_strm0_data        = 'h1234_5678 ;
    std__pe46__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe46__lane21_strm1_cntl        = 'd0         ;
    std__pe46__lane21_strm1_data        = 'h1234_5678 ;
    std__pe46__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe46__lane22_strm0_cntl        = 'd0         ;
    std__pe46__lane22_strm0_data        = 'h1234_5678 ;
    std__pe46__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe46__lane22_strm1_cntl        = 'd0         ;
    std__pe46__lane22_strm1_data        = 'h1234_5678 ;
    std__pe46__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe46__lane23_strm0_cntl        = 'd0         ;
    std__pe46__lane23_strm0_data        = 'h1234_5678 ;
    std__pe46__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe46__lane23_strm1_cntl        = 'd0         ;
    std__pe46__lane23_strm1_data        = 'h1234_5678 ;
    std__pe46__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe46__lane24_strm0_cntl        = 'd0         ;
    std__pe46__lane24_strm0_data        = 'h1234_5678 ;
    std__pe46__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe46__lane24_strm1_cntl        = 'd0         ;
    std__pe46__lane24_strm1_data        = 'h1234_5678 ;
    std__pe46__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe46__lane25_strm0_cntl        = 'd0         ;
    std__pe46__lane25_strm0_data        = 'h1234_5678 ;
    std__pe46__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe46__lane25_strm1_cntl        = 'd0         ;
    std__pe46__lane25_strm1_data        = 'h1234_5678 ;
    std__pe46__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe46__lane26_strm0_cntl        = 'd0         ;
    std__pe46__lane26_strm0_data        = 'h1234_5678 ;
    std__pe46__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe46__lane26_strm1_cntl        = 'd0         ;
    std__pe46__lane26_strm1_data        = 'h1234_5678 ;
    std__pe46__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe46__lane27_strm0_cntl        = 'd0         ;
    std__pe46__lane27_strm0_data        = 'h1234_5678 ;
    std__pe46__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe46__lane27_strm1_cntl        = 'd0         ;
    std__pe46__lane27_strm1_data        = 'h1234_5678 ;
    std__pe46__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe46__lane28_strm0_cntl        = 'd0         ;
    std__pe46__lane28_strm0_data        = 'h1234_5678 ;
    std__pe46__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe46__lane28_strm1_cntl        = 'd0         ;
    std__pe46__lane28_strm1_data        = 'h1234_5678 ;
    std__pe46__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe46__lane29_strm0_cntl        = 'd0         ;
    std__pe46__lane29_strm0_data        = 'h1234_5678 ;
    std__pe46__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe46__lane29_strm1_cntl        = 'd0         ;
    std__pe46__lane29_strm1_data        = 'h1234_5678 ;
    std__pe46__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe46__lane30_strm0_cntl        = 'd0         ;
    std__pe46__lane30_strm0_data        = 'h1234_5678 ;
    std__pe46__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe46__lane30_strm1_cntl        = 'd0         ;
    std__pe46__lane30_strm1_data        = 'h1234_5678 ;
    std__pe46__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe46__lane31_strm0_cntl        = 'd0         ;
    std__pe46__lane31_strm0_data        = 'h1234_5678 ;
    std__pe46__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe46__lane31_strm1_cntl        = 'd0         ;
    std__pe46__lane31_strm1_data        = 'h1234_5678 ;
    std__pe46__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe47__lane0_strm0_cntl        = 'd0         ;
    std__pe47__lane0_strm0_data        = 'h1234_5678 ;
    std__pe47__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe47__lane0_strm1_cntl        = 'd0         ;
    std__pe47__lane0_strm1_data        = 'h1234_5678 ;
    std__pe47__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe47__lane1_strm0_cntl        = 'd0         ;
    std__pe47__lane1_strm0_data        = 'h1234_5678 ;
    std__pe47__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe47__lane1_strm1_cntl        = 'd0         ;
    std__pe47__lane1_strm1_data        = 'h1234_5678 ;
    std__pe47__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe47__lane2_strm0_cntl        = 'd0         ;
    std__pe47__lane2_strm0_data        = 'h1234_5678 ;
    std__pe47__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe47__lane2_strm1_cntl        = 'd0         ;
    std__pe47__lane2_strm1_data        = 'h1234_5678 ;
    std__pe47__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe47__lane3_strm0_cntl        = 'd0         ;
    std__pe47__lane3_strm0_data        = 'h1234_5678 ;
    std__pe47__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe47__lane3_strm1_cntl        = 'd0         ;
    std__pe47__lane3_strm1_data        = 'h1234_5678 ;
    std__pe47__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe47__lane4_strm0_cntl        = 'd0         ;
    std__pe47__lane4_strm0_data        = 'h1234_5678 ;
    std__pe47__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe47__lane4_strm1_cntl        = 'd0         ;
    std__pe47__lane4_strm1_data        = 'h1234_5678 ;
    std__pe47__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe47__lane5_strm0_cntl        = 'd0         ;
    std__pe47__lane5_strm0_data        = 'h1234_5678 ;
    std__pe47__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe47__lane5_strm1_cntl        = 'd0         ;
    std__pe47__lane5_strm1_data        = 'h1234_5678 ;
    std__pe47__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe47__lane6_strm0_cntl        = 'd0         ;
    std__pe47__lane6_strm0_data        = 'h1234_5678 ;
    std__pe47__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe47__lane6_strm1_cntl        = 'd0         ;
    std__pe47__lane6_strm1_data        = 'h1234_5678 ;
    std__pe47__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe47__lane7_strm0_cntl        = 'd0         ;
    std__pe47__lane7_strm0_data        = 'h1234_5678 ;
    std__pe47__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe47__lane7_strm1_cntl        = 'd0         ;
    std__pe47__lane7_strm1_data        = 'h1234_5678 ;
    std__pe47__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe47__lane8_strm0_cntl        = 'd0         ;
    std__pe47__lane8_strm0_data        = 'h1234_5678 ;
    std__pe47__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe47__lane8_strm1_cntl        = 'd0         ;
    std__pe47__lane8_strm1_data        = 'h1234_5678 ;
    std__pe47__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe47__lane9_strm0_cntl        = 'd0         ;
    std__pe47__lane9_strm0_data        = 'h1234_5678 ;
    std__pe47__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe47__lane9_strm1_cntl        = 'd0         ;
    std__pe47__lane9_strm1_data        = 'h1234_5678 ;
    std__pe47__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe47__lane10_strm0_cntl        = 'd0         ;
    std__pe47__lane10_strm0_data        = 'h1234_5678 ;
    std__pe47__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe47__lane10_strm1_cntl        = 'd0         ;
    std__pe47__lane10_strm1_data        = 'h1234_5678 ;
    std__pe47__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe47__lane11_strm0_cntl        = 'd0         ;
    std__pe47__lane11_strm0_data        = 'h1234_5678 ;
    std__pe47__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe47__lane11_strm1_cntl        = 'd0         ;
    std__pe47__lane11_strm1_data        = 'h1234_5678 ;
    std__pe47__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe47__lane12_strm0_cntl        = 'd0         ;
    std__pe47__lane12_strm0_data        = 'h1234_5678 ;
    std__pe47__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe47__lane12_strm1_cntl        = 'd0         ;
    std__pe47__lane12_strm1_data        = 'h1234_5678 ;
    std__pe47__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe47__lane13_strm0_cntl        = 'd0         ;
    std__pe47__lane13_strm0_data        = 'h1234_5678 ;
    std__pe47__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe47__lane13_strm1_cntl        = 'd0         ;
    std__pe47__lane13_strm1_data        = 'h1234_5678 ;
    std__pe47__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe47__lane14_strm0_cntl        = 'd0         ;
    std__pe47__lane14_strm0_data        = 'h1234_5678 ;
    std__pe47__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe47__lane14_strm1_cntl        = 'd0         ;
    std__pe47__lane14_strm1_data        = 'h1234_5678 ;
    std__pe47__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe47__lane15_strm0_cntl        = 'd0         ;
    std__pe47__lane15_strm0_data        = 'h1234_5678 ;
    std__pe47__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe47__lane15_strm1_cntl        = 'd0         ;
    std__pe47__lane15_strm1_data        = 'h1234_5678 ;
    std__pe47__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe47__lane16_strm0_cntl        = 'd0         ;
    std__pe47__lane16_strm0_data        = 'h1234_5678 ;
    std__pe47__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe47__lane16_strm1_cntl        = 'd0         ;
    std__pe47__lane16_strm1_data        = 'h1234_5678 ;
    std__pe47__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe47__lane17_strm0_cntl        = 'd0         ;
    std__pe47__lane17_strm0_data        = 'h1234_5678 ;
    std__pe47__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe47__lane17_strm1_cntl        = 'd0         ;
    std__pe47__lane17_strm1_data        = 'h1234_5678 ;
    std__pe47__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe47__lane18_strm0_cntl        = 'd0         ;
    std__pe47__lane18_strm0_data        = 'h1234_5678 ;
    std__pe47__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe47__lane18_strm1_cntl        = 'd0         ;
    std__pe47__lane18_strm1_data        = 'h1234_5678 ;
    std__pe47__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe47__lane19_strm0_cntl        = 'd0         ;
    std__pe47__lane19_strm0_data        = 'h1234_5678 ;
    std__pe47__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe47__lane19_strm1_cntl        = 'd0         ;
    std__pe47__lane19_strm1_data        = 'h1234_5678 ;
    std__pe47__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe47__lane20_strm0_cntl        = 'd0         ;
    std__pe47__lane20_strm0_data        = 'h1234_5678 ;
    std__pe47__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe47__lane20_strm1_cntl        = 'd0         ;
    std__pe47__lane20_strm1_data        = 'h1234_5678 ;
    std__pe47__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe47__lane21_strm0_cntl        = 'd0         ;
    std__pe47__lane21_strm0_data        = 'h1234_5678 ;
    std__pe47__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe47__lane21_strm1_cntl        = 'd0         ;
    std__pe47__lane21_strm1_data        = 'h1234_5678 ;
    std__pe47__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe47__lane22_strm0_cntl        = 'd0         ;
    std__pe47__lane22_strm0_data        = 'h1234_5678 ;
    std__pe47__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe47__lane22_strm1_cntl        = 'd0         ;
    std__pe47__lane22_strm1_data        = 'h1234_5678 ;
    std__pe47__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe47__lane23_strm0_cntl        = 'd0         ;
    std__pe47__lane23_strm0_data        = 'h1234_5678 ;
    std__pe47__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe47__lane23_strm1_cntl        = 'd0         ;
    std__pe47__lane23_strm1_data        = 'h1234_5678 ;
    std__pe47__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe47__lane24_strm0_cntl        = 'd0         ;
    std__pe47__lane24_strm0_data        = 'h1234_5678 ;
    std__pe47__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe47__lane24_strm1_cntl        = 'd0         ;
    std__pe47__lane24_strm1_data        = 'h1234_5678 ;
    std__pe47__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe47__lane25_strm0_cntl        = 'd0         ;
    std__pe47__lane25_strm0_data        = 'h1234_5678 ;
    std__pe47__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe47__lane25_strm1_cntl        = 'd0         ;
    std__pe47__lane25_strm1_data        = 'h1234_5678 ;
    std__pe47__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe47__lane26_strm0_cntl        = 'd0         ;
    std__pe47__lane26_strm0_data        = 'h1234_5678 ;
    std__pe47__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe47__lane26_strm1_cntl        = 'd0         ;
    std__pe47__lane26_strm1_data        = 'h1234_5678 ;
    std__pe47__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe47__lane27_strm0_cntl        = 'd0         ;
    std__pe47__lane27_strm0_data        = 'h1234_5678 ;
    std__pe47__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe47__lane27_strm1_cntl        = 'd0         ;
    std__pe47__lane27_strm1_data        = 'h1234_5678 ;
    std__pe47__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe47__lane28_strm0_cntl        = 'd0         ;
    std__pe47__lane28_strm0_data        = 'h1234_5678 ;
    std__pe47__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe47__lane28_strm1_cntl        = 'd0         ;
    std__pe47__lane28_strm1_data        = 'h1234_5678 ;
    std__pe47__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe47__lane29_strm0_cntl        = 'd0         ;
    std__pe47__lane29_strm0_data        = 'h1234_5678 ;
    std__pe47__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe47__lane29_strm1_cntl        = 'd0         ;
    std__pe47__lane29_strm1_data        = 'h1234_5678 ;
    std__pe47__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe47__lane30_strm0_cntl        = 'd0         ;
    std__pe47__lane30_strm0_data        = 'h1234_5678 ;
    std__pe47__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe47__lane30_strm1_cntl        = 'd0         ;
    std__pe47__lane30_strm1_data        = 'h1234_5678 ;
    std__pe47__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe47__lane31_strm0_cntl        = 'd0         ;
    std__pe47__lane31_strm0_data        = 'h1234_5678 ;
    std__pe47__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe47__lane31_strm1_cntl        = 'd0         ;
    std__pe47__lane31_strm1_data        = 'h1234_5678 ;
    std__pe47__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe48__lane0_strm0_cntl        = 'd0         ;
    std__pe48__lane0_strm0_data        = 'h1234_5678 ;
    std__pe48__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe48__lane0_strm1_cntl        = 'd0         ;
    std__pe48__lane0_strm1_data        = 'h1234_5678 ;
    std__pe48__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe48__lane1_strm0_cntl        = 'd0         ;
    std__pe48__lane1_strm0_data        = 'h1234_5678 ;
    std__pe48__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe48__lane1_strm1_cntl        = 'd0         ;
    std__pe48__lane1_strm1_data        = 'h1234_5678 ;
    std__pe48__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe48__lane2_strm0_cntl        = 'd0         ;
    std__pe48__lane2_strm0_data        = 'h1234_5678 ;
    std__pe48__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe48__lane2_strm1_cntl        = 'd0         ;
    std__pe48__lane2_strm1_data        = 'h1234_5678 ;
    std__pe48__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe48__lane3_strm0_cntl        = 'd0         ;
    std__pe48__lane3_strm0_data        = 'h1234_5678 ;
    std__pe48__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe48__lane3_strm1_cntl        = 'd0         ;
    std__pe48__lane3_strm1_data        = 'h1234_5678 ;
    std__pe48__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe48__lane4_strm0_cntl        = 'd0         ;
    std__pe48__lane4_strm0_data        = 'h1234_5678 ;
    std__pe48__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe48__lane4_strm1_cntl        = 'd0         ;
    std__pe48__lane4_strm1_data        = 'h1234_5678 ;
    std__pe48__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe48__lane5_strm0_cntl        = 'd0         ;
    std__pe48__lane5_strm0_data        = 'h1234_5678 ;
    std__pe48__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe48__lane5_strm1_cntl        = 'd0         ;
    std__pe48__lane5_strm1_data        = 'h1234_5678 ;
    std__pe48__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe48__lane6_strm0_cntl        = 'd0         ;
    std__pe48__lane6_strm0_data        = 'h1234_5678 ;
    std__pe48__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe48__lane6_strm1_cntl        = 'd0         ;
    std__pe48__lane6_strm1_data        = 'h1234_5678 ;
    std__pe48__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe48__lane7_strm0_cntl        = 'd0         ;
    std__pe48__lane7_strm0_data        = 'h1234_5678 ;
    std__pe48__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe48__lane7_strm1_cntl        = 'd0         ;
    std__pe48__lane7_strm1_data        = 'h1234_5678 ;
    std__pe48__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe48__lane8_strm0_cntl        = 'd0         ;
    std__pe48__lane8_strm0_data        = 'h1234_5678 ;
    std__pe48__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe48__lane8_strm1_cntl        = 'd0         ;
    std__pe48__lane8_strm1_data        = 'h1234_5678 ;
    std__pe48__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe48__lane9_strm0_cntl        = 'd0         ;
    std__pe48__lane9_strm0_data        = 'h1234_5678 ;
    std__pe48__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe48__lane9_strm1_cntl        = 'd0         ;
    std__pe48__lane9_strm1_data        = 'h1234_5678 ;
    std__pe48__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe48__lane10_strm0_cntl        = 'd0         ;
    std__pe48__lane10_strm0_data        = 'h1234_5678 ;
    std__pe48__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe48__lane10_strm1_cntl        = 'd0         ;
    std__pe48__lane10_strm1_data        = 'h1234_5678 ;
    std__pe48__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe48__lane11_strm0_cntl        = 'd0         ;
    std__pe48__lane11_strm0_data        = 'h1234_5678 ;
    std__pe48__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe48__lane11_strm1_cntl        = 'd0         ;
    std__pe48__lane11_strm1_data        = 'h1234_5678 ;
    std__pe48__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe48__lane12_strm0_cntl        = 'd0         ;
    std__pe48__lane12_strm0_data        = 'h1234_5678 ;
    std__pe48__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe48__lane12_strm1_cntl        = 'd0         ;
    std__pe48__lane12_strm1_data        = 'h1234_5678 ;
    std__pe48__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe48__lane13_strm0_cntl        = 'd0         ;
    std__pe48__lane13_strm0_data        = 'h1234_5678 ;
    std__pe48__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe48__lane13_strm1_cntl        = 'd0         ;
    std__pe48__lane13_strm1_data        = 'h1234_5678 ;
    std__pe48__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe48__lane14_strm0_cntl        = 'd0         ;
    std__pe48__lane14_strm0_data        = 'h1234_5678 ;
    std__pe48__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe48__lane14_strm1_cntl        = 'd0         ;
    std__pe48__lane14_strm1_data        = 'h1234_5678 ;
    std__pe48__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe48__lane15_strm0_cntl        = 'd0         ;
    std__pe48__lane15_strm0_data        = 'h1234_5678 ;
    std__pe48__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe48__lane15_strm1_cntl        = 'd0         ;
    std__pe48__lane15_strm1_data        = 'h1234_5678 ;
    std__pe48__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe48__lane16_strm0_cntl        = 'd0         ;
    std__pe48__lane16_strm0_data        = 'h1234_5678 ;
    std__pe48__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe48__lane16_strm1_cntl        = 'd0         ;
    std__pe48__lane16_strm1_data        = 'h1234_5678 ;
    std__pe48__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe48__lane17_strm0_cntl        = 'd0         ;
    std__pe48__lane17_strm0_data        = 'h1234_5678 ;
    std__pe48__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe48__lane17_strm1_cntl        = 'd0         ;
    std__pe48__lane17_strm1_data        = 'h1234_5678 ;
    std__pe48__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe48__lane18_strm0_cntl        = 'd0         ;
    std__pe48__lane18_strm0_data        = 'h1234_5678 ;
    std__pe48__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe48__lane18_strm1_cntl        = 'd0         ;
    std__pe48__lane18_strm1_data        = 'h1234_5678 ;
    std__pe48__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe48__lane19_strm0_cntl        = 'd0         ;
    std__pe48__lane19_strm0_data        = 'h1234_5678 ;
    std__pe48__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe48__lane19_strm1_cntl        = 'd0         ;
    std__pe48__lane19_strm1_data        = 'h1234_5678 ;
    std__pe48__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe48__lane20_strm0_cntl        = 'd0         ;
    std__pe48__lane20_strm0_data        = 'h1234_5678 ;
    std__pe48__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe48__lane20_strm1_cntl        = 'd0         ;
    std__pe48__lane20_strm1_data        = 'h1234_5678 ;
    std__pe48__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe48__lane21_strm0_cntl        = 'd0         ;
    std__pe48__lane21_strm0_data        = 'h1234_5678 ;
    std__pe48__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe48__lane21_strm1_cntl        = 'd0         ;
    std__pe48__lane21_strm1_data        = 'h1234_5678 ;
    std__pe48__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe48__lane22_strm0_cntl        = 'd0         ;
    std__pe48__lane22_strm0_data        = 'h1234_5678 ;
    std__pe48__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe48__lane22_strm1_cntl        = 'd0         ;
    std__pe48__lane22_strm1_data        = 'h1234_5678 ;
    std__pe48__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe48__lane23_strm0_cntl        = 'd0         ;
    std__pe48__lane23_strm0_data        = 'h1234_5678 ;
    std__pe48__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe48__lane23_strm1_cntl        = 'd0         ;
    std__pe48__lane23_strm1_data        = 'h1234_5678 ;
    std__pe48__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe48__lane24_strm0_cntl        = 'd0         ;
    std__pe48__lane24_strm0_data        = 'h1234_5678 ;
    std__pe48__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe48__lane24_strm1_cntl        = 'd0         ;
    std__pe48__lane24_strm1_data        = 'h1234_5678 ;
    std__pe48__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe48__lane25_strm0_cntl        = 'd0         ;
    std__pe48__lane25_strm0_data        = 'h1234_5678 ;
    std__pe48__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe48__lane25_strm1_cntl        = 'd0         ;
    std__pe48__lane25_strm1_data        = 'h1234_5678 ;
    std__pe48__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe48__lane26_strm0_cntl        = 'd0         ;
    std__pe48__lane26_strm0_data        = 'h1234_5678 ;
    std__pe48__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe48__lane26_strm1_cntl        = 'd0         ;
    std__pe48__lane26_strm1_data        = 'h1234_5678 ;
    std__pe48__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe48__lane27_strm0_cntl        = 'd0         ;
    std__pe48__lane27_strm0_data        = 'h1234_5678 ;
    std__pe48__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe48__lane27_strm1_cntl        = 'd0         ;
    std__pe48__lane27_strm1_data        = 'h1234_5678 ;
    std__pe48__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe48__lane28_strm0_cntl        = 'd0         ;
    std__pe48__lane28_strm0_data        = 'h1234_5678 ;
    std__pe48__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe48__lane28_strm1_cntl        = 'd0         ;
    std__pe48__lane28_strm1_data        = 'h1234_5678 ;
    std__pe48__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe48__lane29_strm0_cntl        = 'd0         ;
    std__pe48__lane29_strm0_data        = 'h1234_5678 ;
    std__pe48__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe48__lane29_strm1_cntl        = 'd0         ;
    std__pe48__lane29_strm1_data        = 'h1234_5678 ;
    std__pe48__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe48__lane30_strm0_cntl        = 'd0         ;
    std__pe48__lane30_strm0_data        = 'h1234_5678 ;
    std__pe48__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe48__lane30_strm1_cntl        = 'd0         ;
    std__pe48__lane30_strm1_data        = 'h1234_5678 ;
    std__pe48__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe48__lane31_strm0_cntl        = 'd0         ;
    std__pe48__lane31_strm0_data        = 'h1234_5678 ;
    std__pe48__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe48__lane31_strm1_cntl        = 'd0         ;
    std__pe48__lane31_strm1_data        = 'h1234_5678 ;
    std__pe48__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe49__lane0_strm0_cntl        = 'd0         ;
    std__pe49__lane0_strm0_data        = 'h1234_5678 ;
    std__pe49__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe49__lane0_strm1_cntl        = 'd0         ;
    std__pe49__lane0_strm1_data        = 'h1234_5678 ;
    std__pe49__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe49__lane1_strm0_cntl        = 'd0         ;
    std__pe49__lane1_strm0_data        = 'h1234_5678 ;
    std__pe49__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe49__lane1_strm1_cntl        = 'd0         ;
    std__pe49__lane1_strm1_data        = 'h1234_5678 ;
    std__pe49__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe49__lane2_strm0_cntl        = 'd0         ;
    std__pe49__lane2_strm0_data        = 'h1234_5678 ;
    std__pe49__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe49__lane2_strm1_cntl        = 'd0         ;
    std__pe49__lane2_strm1_data        = 'h1234_5678 ;
    std__pe49__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe49__lane3_strm0_cntl        = 'd0         ;
    std__pe49__lane3_strm0_data        = 'h1234_5678 ;
    std__pe49__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe49__lane3_strm1_cntl        = 'd0         ;
    std__pe49__lane3_strm1_data        = 'h1234_5678 ;
    std__pe49__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe49__lane4_strm0_cntl        = 'd0         ;
    std__pe49__lane4_strm0_data        = 'h1234_5678 ;
    std__pe49__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe49__lane4_strm1_cntl        = 'd0         ;
    std__pe49__lane4_strm1_data        = 'h1234_5678 ;
    std__pe49__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe49__lane5_strm0_cntl        = 'd0         ;
    std__pe49__lane5_strm0_data        = 'h1234_5678 ;
    std__pe49__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe49__lane5_strm1_cntl        = 'd0         ;
    std__pe49__lane5_strm1_data        = 'h1234_5678 ;
    std__pe49__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe49__lane6_strm0_cntl        = 'd0         ;
    std__pe49__lane6_strm0_data        = 'h1234_5678 ;
    std__pe49__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe49__lane6_strm1_cntl        = 'd0         ;
    std__pe49__lane6_strm1_data        = 'h1234_5678 ;
    std__pe49__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe49__lane7_strm0_cntl        = 'd0         ;
    std__pe49__lane7_strm0_data        = 'h1234_5678 ;
    std__pe49__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe49__lane7_strm1_cntl        = 'd0         ;
    std__pe49__lane7_strm1_data        = 'h1234_5678 ;
    std__pe49__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe49__lane8_strm0_cntl        = 'd0         ;
    std__pe49__lane8_strm0_data        = 'h1234_5678 ;
    std__pe49__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe49__lane8_strm1_cntl        = 'd0         ;
    std__pe49__lane8_strm1_data        = 'h1234_5678 ;
    std__pe49__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe49__lane9_strm0_cntl        = 'd0         ;
    std__pe49__lane9_strm0_data        = 'h1234_5678 ;
    std__pe49__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe49__lane9_strm1_cntl        = 'd0         ;
    std__pe49__lane9_strm1_data        = 'h1234_5678 ;
    std__pe49__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe49__lane10_strm0_cntl        = 'd0         ;
    std__pe49__lane10_strm0_data        = 'h1234_5678 ;
    std__pe49__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe49__lane10_strm1_cntl        = 'd0         ;
    std__pe49__lane10_strm1_data        = 'h1234_5678 ;
    std__pe49__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe49__lane11_strm0_cntl        = 'd0         ;
    std__pe49__lane11_strm0_data        = 'h1234_5678 ;
    std__pe49__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe49__lane11_strm1_cntl        = 'd0         ;
    std__pe49__lane11_strm1_data        = 'h1234_5678 ;
    std__pe49__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe49__lane12_strm0_cntl        = 'd0         ;
    std__pe49__lane12_strm0_data        = 'h1234_5678 ;
    std__pe49__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe49__lane12_strm1_cntl        = 'd0         ;
    std__pe49__lane12_strm1_data        = 'h1234_5678 ;
    std__pe49__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe49__lane13_strm0_cntl        = 'd0         ;
    std__pe49__lane13_strm0_data        = 'h1234_5678 ;
    std__pe49__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe49__lane13_strm1_cntl        = 'd0         ;
    std__pe49__lane13_strm1_data        = 'h1234_5678 ;
    std__pe49__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe49__lane14_strm0_cntl        = 'd0         ;
    std__pe49__lane14_strm0_data        = 'h1234_5678 ;
    std__pe49__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe49__lane14_strm1_cntl        = 'd0         ;
    std__pe49__lane14_strm1_data        = 'h1234_5678 ;
    std__pe49__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe49__lane15_strm0_cntl        = 'd0         ;
    std__pe49__lane15_strm0_data        = 'h1234_5678 ;
    std__pe49__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe49__lane15_strm1_cntl        = 'd0         ;
    std__pe49__lane15_strm1_data        = 'h1234_5678 ;
    std__pe49__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe49__lane16_strm0_cntl        = 'd0         ;
    std__pe49__lane16_strm0_data        = 'h1234_5678 ;
    std__pe49__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe49__lane16_strm1_cntl        = 'd0         ;
    std__pe49__lane16_strm1_data        = 'h1234_5678 ;
    std__pe49__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe49__lane17_strm0_cntl        = 'd0         ;
    std__pe49__lane17_strm0_data        = 'h1234_5678 ;
    std__pe49__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe49__lane17_strm1_cntl        = 'd0         ;
    std__pe49__lane17_strm1_data        = 'h1234_5678 ;
    std__pe49__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe49__lane18_strm0_cntl        = 'd0         ;
    std__pe49__lane18_strm0_data        = 'h1234_5678 ;
    std__pe49__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe49__lane18_strm1_cntl        = 'd0         ;
    std__pe49__lane18_strm1_data        = 'h1234_5678 ;
    std__pe49__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe49__lane19_strm0_cntl        = 'd0         ;
    std__pe49__lane19_strm0_data        = 'h1234_5678 ;
    std__pe49__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe49__lane19_strm1_cntl        = 'd0         ;
    std__pe49__lane19_strm1_data        = 'h1234_5678 ;
    std__pe49__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe49__lane20_strm0_cntl        = 'd0         ;
    std__pe49__lane20_strm0_data        = 'h1234_5678 ;
    std__pe49__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe49__lane20_strm1_cntl        = 'd0         ;
    std__pe49__lane20_strm1_data        = 'h1234_5678 ;
    std__pe49__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe49__lane21_strm0_cntl        = 'd0         ;
    std__pe49__lane21_strm0_data        = 'h1234_5678 ;
    std__pe49__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe49__lane21_strm1_cntl        = 'd0         ;
    std__pe49__lane21_strm1_data        = 'h1234_5678 ;
    std__pe49__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe49__lane22_strm0_cntl        = 'd0         ;
    std__pe49__lane22_strm0_data        = 'h1234_5678 ;
    std__pe49__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe49__lane22_strm1_cntl        = 'd0         ;
    std__pe49__lane22_strm1_data        = 'h1234_5678 ;
    std__pe49__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe49__lane23_strm0_cntl        = 'd0         ;
    std__pe49__lane23_strm0_data        = 'h1234_5678 ;
    std__pe49__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe49__lane23_strm1_cntl        = 'd0         ;
    std__pe49__lane23_strm1_data        = 'h1234_5678 ;
    std__pe49__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe49__lane24_strm0_cntl        = 'd0         ;
    std__pe49__lane24_strm0_data        = 'h1234_5678 ;
    std__pe49__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe49__lane24_strm1_cntl        = 'd0         ;
    std__pe49__lane24_strm1_data        = 'h1234_5678 ;
    std__pe49__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe49__lane25_strm0_cntl        = 'd0         ;
    std__pe49__lane25_strm0_data        = 'h1234_5678 ;
    std__pe49__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe49__lane25_strm1_cntl        = 'd0         ;
    std__pe49__lane25_strm1_data        = 'h1234_5678 ;
    std__pe49__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe49__lane26_strm0_cntl        = 'd0         ;
    std__pe49__lane26_strm0_data        = 'h1234_5678 ;
    std__pe49__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe49__lane26_strm1_cntl        = 'd0         ;
    std__pe49__lane26_strm1_data        = 'h1234_5678 ;
    std__pe49__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe49__lane27_strm0_cntl        = 'd0         ;
    std__pe49__lane27_strm0_data        = 'h1234_5678 ;
    std__pe49__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe49__lane27_strm1_cntl        = 'd0         ;
    std__pe49__lane27_strm1_data        = 'h1234_5678 ;
    std__pe49__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe49__lane28_strm0_cntl        = 'd0         ;
    std__pe49__lane28_strm0_data        = 'h1234_5678 ;
    std__pe49__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe49__lane28_strm1_cntl        = 'd0         ;
    std__pe49__lane28_strm1_data        = 'h1234_5678 ;
    std__pe49__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe49__lane29_strm0_cntl        = 'd0         ;
    std__pe49__lane29_strm0_data        = 'h1234_5678 ;
    std__pe49__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe49__lane29_strm1_cntl        = 'd0         ;
    std__pe49__lane29_strm1_data        = 'h1234_5678 ;
    std__pe49__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe49__lane30_strm0_cntl        = 'd0         ;
    std__pe49__lane30_strm0_data        = 'h1234_5678 ;
    std__pe49__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe49__lane30_strm1_cntl        = 'd0         ;
    std__pe49__lane30_strm1_data        = 'h1234_5678 ;
    std__pe49__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe49__lane31_strm0_cntl        = 'd0         ;
    std__pe49__lane31_strm0_data        = 'h1234_5678 ;
    std__pe49__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe49__lane31_strm1_cntl        = 'd0         ;
    std__pe49__lane31_strm1_data        = 'h1234_5678 ;
    std__pe49__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe50__lane0_strm0_cntl        = 'd0         ;
    std__pe50__lane0_strm0_data        = 'h1234_5678 ;
    std__pe50__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe50__lane0_strm1_cntl        = 'd0         ;
    std__pe50__lane0_strm1_data        = 'h1234_5678 ;
    std__pe50__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe50__lane1_strm0_cntl        = 'd0         ;
    std__pe50__lane1_strm0_data        = 'h1234_5678 ;
    std__pe50__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe50__lane1_strm1_cntl        = 'd0         ;
    std__pe50__lane1_strm1_data        = 'h1234_5678 ;
    std__pe50__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe50__lane2_strm0_cntl        = 'd0         ;
    std__pe50__lane2_strm0_data        = 'h1234_5678 ;
    std__pe50__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe50__lane2_strm1_cntl        = 'd0         ;
    std__pe50__lane2_strm1_data        = 'h1234_5678 ;
    std__pe50__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe50__lane3_strm0_cntl        = 'd0         ;
    std__pe50__lane3_strm0_data        = 'h1234_5678 ;
    std__pe50__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe50__lane3_strm1_cntl        = 'd0         ;
    std__pe50__lane3_strm1_data        = 'h1234_5678 ;
    std__pe50__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe50__lane4_strm0_cntl        = 'd0         ;
    std__pe50__lane4_strm0_data        = 'h1234_5678 ;
    std__pe50__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe50__lane4_strm1_cntl        = 'd0         ;
    std__pe50__lane4_strm1_data        = 'h1234_5678 ;
    std__pe50__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe50__lane5_strm0_cntl        = 'd0         ;
    std__pe50__lane5_strm0_data        = 'h1234_5678 ;
    std__pe50__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe50__lane5_strm1_cntl        = 'd0         ;
    std__pe50__lane5_strm1_data        = 'h1234_5678 ;
    std__pe50__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe50__lane6_strm0_cntl        = 'd0         ;
    std__pe50__lane6_strm0_data        = 'h1234_5678 ;
    std__pe50__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe50__lane6_strm1_cntl        = 'd0         ;
    std__pe50__lane6_strm1_data        = 'h1234_5678 ;
    std__pe50__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe50__lane7_strm0_cntl        = 'd0         ;
    std__pe50__lane7_strm0_data        = 'h1234_5678 ;
    std__pe50__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe50__lane7_strm1_cntl        = 'd0         ;
    std__pe50__lane7_strm1_data        = 'h1234_5678 ;
    std__pe50__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe50__lane8_strm0_cntl        = 'd0         ;
    std__pe50__lane8_strm0_data        = 'h1234_5678 ;
    std__pe50__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe50__lane8_strm1_cntl        = 'd0         ;
    std__pe50__lane8_strm1_data        = 'h1234_5678 ;
    std__pe50__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe50__lane9_strm0_cntl        = 'd0         ;
    std__pe50__lane9_strm0_data        = 'h1234_5678 ;
    std__pe50__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe50__lane9_strm1_cntl        = 'd0         ;
    std__pe50__lane9_strm1_data        = 'h1234_5678 ;
    std__pe50__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe50__lane10_strm0_cntl        = 'd0         ;
    std__pe50__lane10_strm0_data        = 'h1234_5678 ;
    std__pe50__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe50__lane10_strm1_cntl        = 'd0         ;
    std__pe50__lane10_strm1_data        = 'h1234_5678 ;
    std__pe50__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe50__lane11_strm0_cntl        = 'd0         ;
    std__pe50__lane11_strm0_data        = 'h1234_5678 ;
    std__pe50__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe50__lane11_strm1_cntl        = 'd0         ;
    std__pe50__lane11_strm1_data        = 'h1234_5678 ;
    std__pe50__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe50__lane12_strm0_cntl        = 'd0         ;
    std__pe50__lane12_strm0_data        = 'h1234_5678 ;
    std__pe50__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe50__lane12_strm1_cntl        = 'd0         ;
    std__pe50__lane12_strm1_data        = 'h1234_5678 ;
    std__pe50__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe50__lane13_strm0_cntl        = 'd0         ;
    std__pe50__lane13_strm0_data        = 'h1234_5678 ;
    std__pe50__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe50__lane13_strm1_cntl        = 'd0         ;
    std__pe50__lane13_strm1_data        = 'h1234_5678 ;
    std__pe50__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe50__lane14_strm0_cntl        = 'd0         ;
    std__pe50__lane14_strm0_data        = 'h1234_5678 ;
    std__pe50__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe50__lane14_strm1_cntl        = 'd0         ;
    std__pe50__lane14_strm1_data        = 'h1234_5678 ;
    std__pe50__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe50__lane15_strm0_cntl        = 'd0         ;
    std__pe50__lane15_strm0_data        = 'h1234_5678 ;
    std__pe50__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe50__lane15_strm1_cntl        = 'd0         ;
    std__pe50__lane15_strm1_data        = 'h1234_5678 ;
    std__pe50__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe50__lane16_strm0_cntl        = 'd0         ;
    std__pe50__lane16_strm0_data        = 'h1234_5678 ;
    std__pe50__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe50__lane16_strm1_cntl        = 'd0         ;
    std__pe50__lane16_strm1_data        = 'h1234_5678 ;
    std__pe50__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe50__lane17_strm0_cntl        = 'd0         ;
    std__pe50__lane17_strm0_data        = 'h1234_5678 ;
    std__pe50__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe50__lane17_strm1_cntl        = 'd0         ;
    std__pe50__lane17_strm1_data        = 'h1234_5678 ;
    std__pe50__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe50__lane18_strm0_cntl        = 'd0         ;
    std__pe50__lane18_strm0_data        = 'h1234_5678 ;
    std__pe50__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe50__lane18_strm1_cntl        = 'd0         ;
    std__pe50__lane18_strm1_data        = 'h1234_5678 ;
    std__pe50__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe50__lane19_strm0_cntl        = 'd0         ;
    std__pe50__lane19_strm0_data        = 'h1234_5678 ;
    std__pe50__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe50__lane19_strm1_cntl        = 'd0         ;
    std__pe50__lane19_strm1_data        = 'h1234_5678 ;
    std__pe50__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe50__lane20_strm0_cntl        = 'd0         ;
    std__pe50__lane20_strm0_data        = 'h1234_5678 ;
    std__pe50__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe50__lane20_strm1_cntl        = 'd0         ;
    std__pe50__lane20_strm1_data        = 'h1234_5678 ;
    std__pe50__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe50__lane21_strm0_cntl        = 'd0         ;
    std__pe50__lane21_strm0_data        = 'h1234_5678 ;
    std__pe50__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe50__lane21_strm1_cntl        = 'd0         ;
    std__pe50__lane21_strm1_data        = 'h1234_5678 ;
    std__pe50__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe50__lane22_strm0_cntl        = 'd0         ;
    std__pe50__lane22_strm0_data        = 'h1234_5678 ;
    std__pe50__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe50__lane22_strm1_cntl        = 'd0         ;
    std__pe50__lane22_strm1_data        = 'h1234_5678 ;
    std__pe50__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe50__lane23_strm0_cntl        = 'd0         ;
    std__pe50__lane23_strm0_data        = 'h1234_5678 ;
    std__pe50__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe50__lane23_strm1_cntl        = 'd0         ;
    std__pe50__lane23_strm1_data        = 'h1234_5678 ;
    std__pe50__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe50__lane24_strm0_cntl        = 'd0         ;
    std__pe50__lane24_strm0_data        = 'h1234_5678 ;
    std__pe50__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe50__lane24_strm1_cntl        = 'd0         ;
    std__pe50__lane24_strm1_data        = 'h1234_5678 ;
    std__pe50__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe50__lane25_strm0_cntl        = 'd0         ;
    std__pe50__lane25_strm0_data        = 'h1234_5678 ;
    std__pe50__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe50__lane25_strm1_cntl        = 'd0         ;
    std__pe50__lane25_strm1_data        = 'h1234_5678 ;
    std__pe50__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe50__lane26_strm0_cntl        = 'd0         ;
    std__pe50__lane26_strm0_data        = 'h1234_5678 ;
    std__pe50__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe50__lane26_strm1_cntl        = 'd0         ;
    std__pe50__lane26_strm1_data        = 'h1234_5678 ;
    std__pe50__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe50__lane27_strm0_cntl        = 'd0         ;
    std__pe50__lane27_strm0_data        = 'h1234_5678 ;
    std__pe50__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe50__lane27_strm1_cntl        = 'd0         ;
    std__pe50__lane27_strm1_data        = 'h1234_5678 ;
    std__pe50__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe50__lane28_strm0_cntl        = 'd0         ;
    std__pe50__lane28_strm0_data        = 'h1234_5678 ;
    std__pe50__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe50__lane28_strm1_cntl        = 'd0         ;
    std__pe50__lane28_strm1_data        = 'h1234_5678 ;
    std__pe50__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe50__lane29_strm0_cntl        = 'd0         ;
    std__pe50__lane29_strm0_data        = 'h1234_5678 ;
    std__pe50__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe50__lane29_strm1_cntl        = 'd0         ;
    std__pe50__lane29_strm1_data        = 'h1234_5678 ;
    std__pe50__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe50__lane30_strm0_cntl        = 'd0         ;
    std__pe50__lane30_strm0_data        = 'h1234_5678 ;
    std__pe50__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe50__lane30_strm1_cntl        = 'd0         ;
    std__pe50__lane30_strm1_data        = 'h1234_5678 ;
    std__pe50__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe50__lane31_strm0_cntl        = 'd0         ;
    std__pe50__lane31_strm0_data        = 'h1234_5678 ;
    std__pe50__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe50__lane31_strm1_cntl        = 'd0         ;
    std__pe50__lane31_strm1_data        = 'h1234_5678 ;
    std__pe50__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe51__lane0_strm0_cntl        = 'd0         ;
    std__pe51__lane0_strm0_data        = 'h1234_5678 ;
    std__pe51__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe51__lane0_strm1_cntl        = 'd0         ;
    std__pe51__lane0_strm1_data        = 'h1234_5678 ;
    std__pe51__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe51__lane1_strm0_cntl        = 'd0         ;
    std__pe51__lane1_strm0_data        = 'h1234_5678 ;
    std__pe51__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe51__lane1_strm1_cntl        = 'd0         ;
    std__pe51__lane1_strm1_data        = 'h1234_5678 ;
    std__pe51__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe51__lane2_strm0_cntl        = 'd0         ;
    std__pe51__lane2_strm0_data        = 'h1234_5678 ;
    std__pe51__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe51__lane2_strm1_cntl        = 'd0         ;
    std__pe51__lane2_strm1_data        = 'h1234_5678 ;
    std__pe51__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe51__lane3_strm0_cntl        = 'd0         ;
    std__pe51__lane3_strm0_data        = 'h1234_5678 ;
    std__pe51__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe51__lane3_strm1_cntl        = 'd0         ;
    std__pe51__lane3_strm1_data        = 'h1234_5678 ;
    std__pe51__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe51__lane4_strm0_cntl        = 'd0         ;
    std__pe51__lane4_strm0_data        = 'h1234_5678 ;
    std__pe51__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe51__lane4_strm1_cntl        = 'd0         ;
    std__pe51__lane4_strm1_data        = 'h1234_5678 ;
    std__pe51__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe51__lane5_strm0_cntl        = 'd0         ;
    std__pe51__lane5_strm0_data        = 'h1234_5678 ;
    std__pe51__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe51__lane5_strm1_cntl        = 'd0         ;
    std__pe51__lane5_strm1_data        = 'h1234_5678 ;
    std__pe51__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe51__lane6_strm0_cntl        = 'd0         ;
    std__pe51__lane6_strm0_data        = 'h1234_5678 ;
    std__pe51__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe51__lane6_strm1_cntl        = 'd0         ;
    std__pe51__lane6_strm1_data        = 'h1234_5678 ;
    std__pe51__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe51__lane7_strm0_cntl        = 'd0         ;
    std__pe51__lane7_strm0_data        = 'h1234_5678 ;
    std__pe51__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe51__lane7_strm1_cntl        = 'd0         ;
    std__pe51__lane7_strm1_data        = 'h1234_5678 ;
    std__pe51__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe51__lane8_strm0_cntl        = 'd0         ;
    std__pe51__lane8_strm0_data        = 'h1234_5678 ;
    std__pe51__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe51__lane8_strm1_cntl        = 'd0         ;
    std__pe51__lane8_strm1_data        = 'h1234_5678 ;
    std__pe51__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe51__lane9_strm0_cntl        = 'd0         ;
    std__pe51__lane9_strm0_data        = 'h1234_5678 ;
    std__pe51__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe51__lane9_strm1_cntl        = 'd0         ;
    std__pe51__lane9_strm1_data        = 'h1234_5678 ;
    std__pe51__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe51__lane10_strm0_cntl        = 'd0         ;
    std__pe51__lane10_strm0_data        = 'h1234_5678 ;
    std__pe51__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe51__lane10_strm1_cntl        = 'd0         ;
    std__pe51__lane10_strm1_data        = 'h1234_5678 ;
    std__pe51__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe51__lane11_strm0_cntl        = 'd0         ;
    std__pe51__lane11_strm0_data        = 'h1234_5678 ;
    std__pe51__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe51__lane11_strm1_cntl        = 'd0         ;
    std__pe51__lane11_strm1_data        = 'h1234_5678 ;
    std__pe51__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe51__lane12_strm0_cntl        = 'd0         ;
    std__pe51__lane12_strm0_data        = 'h1234_5678 ;
    std__pe51__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe51__lane12_strm1_cntl        = 'd0         ;
    std__pe51__lane12_strm1_data        = 'h1234_5678 ;
    std__pe51__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe51__lane13_strm0_cntl        = 'd0         ;
    std__pe51__lane13_strm0_data        = 'h1234_5678 ;
    std__pe51__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe51__lane13_strm1_cntl        = 'd0         ;
    std__pe51__lane13_strm1_data        = 'h1234_5678 ;
    std__pe51__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe51__lane14_strm0_cntl        = 'd0         ;
    std__pe51__lane14_strm0_data        = 'h1234_5678 ;
    std__pe51__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe51__lane14_strm1_cntl        = 'd0         ;
    std__pe51__lane14_strm1_data        = 'h1234_5678 ;
    std__pe51__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe51__lane15_strm0_cntl        = 'd0         ;
    std__pe51__lane15_strm0_data        = 'h1234_5678 ;
    std__pe51__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe51__lane15_strm1_cntl        = 'd0         ;
    std__pe51__lane15_strm1_data        = 'h1234_5678 ;
    std__pe51__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe51__lane16_strm0_cntl        = 'd0         ;
    std__pe51__lane16_strm0_data        = 'h1234_5678 ;
    std__pe51__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe51__lane16_strm1_cntl        = 'd0         ;
    std__pe51__lane16_strm1_data        = 'h1234_5678 ;
    std__pe51__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe51__lane17_strm0_cntl        = 'd0         ;
    std__pe51__lane17_strm0_data        = 'h1234_5678 ;
    std__pe51__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe51__lane17_strm1_cntl        = 'd0         ;
    std__pe51__lane17_strm1_data        = 'h1234_5678 ;
    std__pe51__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe51__lane18_strm0_cntl        = 'd0         ;
    std__pe51__lane18_strm0_data        = 'h1234_5678 ;
    std__pe51__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe51__lane18_strm1_cntl        = 'd0         ;
    std__pe51__lane18_strm1_data        = 'h1234_5678 ;
    std__pe51__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe51__lane19_strm0_cntl        = 'd0         ;
    std__pe51__lane19_strm0_data        = 'h1234_5678 ;
    std__pe51__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe51__lane19_strm1_cntl        = 'd0         ;
    std__pe51__lane19_strm1_data        = 'h1234_5678 ;
    std__pe51__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe51__lane20_strm0_cntl        = 'd0         ;
    std__pe51__lane20_strm0_data        = 'h1234_5678 ;
    std__pe51__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe51__lane20_strm1_cntl        = 'd0         ;
    std__pe51__lane20_strm1_data        = 'h1234_5678 ;
    std__pe51__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe51__lane21_strm0_cntl        = 'd0         ;
    std__pe51__lane21_strm0_data        = 'h1234_5678 ;
    std__pe51__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe51__lane21_strm1_cntl        = 'd0         ;
    std__pe51__lane21_strm1_data        = 'h1234_5678 ;
    std__pe51__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe51__lane22_strm0_cntl        = 'd0         ;
    std__pe51__lane22_strm0_data        = 'h1234_5678 ;
    std__pe51__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe51__lane22_strm1_cntl        = 'd0         ;
    std__pe51__lane22_strm1_data        = 'h1234_5678 ;
    std__pe51__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe51__lane23_strm0_cntl        = 'd0         ;
    std__pe51__lane23_strm0_data        = 'h1234_5678 ;
    std__pe51__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe51__lane23_strm1_cntl        = 'd0         ;
    std__pe51__lane23_strm1_data        = 'h1234_5678 ;
    std__pe51__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe51__lane24_strm0_cntl        = 'd0         ;
    std__pe51__lane24_strm0_data        = 'h1234_5678 ;
    std__pe51__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe51__lane24_strm1_cntl        = 'd0         ;
    std__pe51__lane24_strm1_data        = 'h1234_5678 ;
    std__pe51__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe51__lane25_strm0_cntl        = 'd0         ;
    std__pe51__lane25_strm0_data        = 'h1234_5678 ;
    std__pe51__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe51__lane25_strm1_cntl        = 'd0         ;
    std__pe51__lane25_strm1_data        = 'h1234_5678 ;
    std__pe51__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe51__lane26_strm0_cntl        = 'd0         ;
    std__pe51__lane26_strm0_data        = 'h1234_5678 ;
    std__pe51__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe51__lane26_strm1_cntl        = 'd0         ;
    std__pe51__lane26_strm1_data        = 'h1234_5678 ;
    std__pe51__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe51__lane27_strm0_cntl        = 'd0         ;
    std__pe51__lane27_strm0_data        = 'h1234_5678 ;
    std__pe51__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe51__lane27_strm1_cntl        = 'd0         ;
    std__pe51__lane27_strm1_data        = 'h1234_5678 ;
    std__pe51__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe51__lane28_strm0_cntl        = 'd0         ;
    std__pe51__lane28_strm0_data        = 'h1234_5678 ;
    std__pe51__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe51__lane28_strm1_cntl        = 'd0         ;
    std__pe51__lane28_strm1_data        = 'h1234_5678 ;
    std__pe51__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe51__lane29_strm0_cntl        = 'd0         ;
    std__pe51__lane29_strm0_data        = 'h1234_5678 ;
    std__pe51__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe51__lane29_strm1_cntl        = 'd0         ;
    std__pe51__lane29_strm1_data        = 'h1234_5678 ;
    std__pe51__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe51__lane30_strm0_cntl        = 'd0         ;
    std__pe51__lane30_strm0_data        = 'h1234_5678 ;
    std__pe51__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe51__lane30_strm1_cntl        = 'd0         ;
    std__pe51__lane30_strm1_data        = 'h1234_5678 ;
    std__pe51__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe51__lane31_strm0_cntl        = 'd0         ;
    std__pe51__lane31_strm0_data        = 'h1234_5678 ;
    std__pe51__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe51__lane31_strm1_cntl        = 'd0         ;
    std__pe51__lane31_strm1_data        = 'h1234_5678 ;
    std__pe51__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe52__lane0_strm0_cntl        = 'd0         ;
    std__pe52__lane0_strm0_data        = 'h1234_5678 ;
    std__pe52__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe52__lane0_strm1_cntl        = 'd0         ;
    std__pe52__lane0_strm1_data        = 'h1234_5678 ;
    std__pe52__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe52__lane1_strm0_cntl        = 'd0         ;
    std__pe52__lane1_strm0_data        = 'h1234_5678 ;
    std__pe52__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe52__lane1_strm1_cntl        = 'd0         ;
    std__pe52__lane1_strm1_data        = 'h1234_5678 ;
    std__pe52__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe52__lane2_strm0_cntl        = 'd0         ;
    std__pe52__lane2_strm0_data        = 'h1234_5678 ;
    std__pe52__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe52__lane2_strm1_cntl        = 'd0         ;
    std__pe52__lane2_strm1_data        = 'h1234_5678 ;
    std__pe52__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe52__lane3_strm0_cntl        = 'd0         ;
    std__pe52__lane3_strm0_data        = 'h1234_5678 ;
    std__pe52__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe52__lane3_strm1_cntl        = 'd0         ;
    std__pe52__lane3_strm1_data        = 'h1234_5678 ;
    std__pe52__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe52__lane4_strm0_cntl        = 'd0         ;
    std__pe52__lane4_strm0_data        = 'h1234_5678 ;
    std__pe52__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe52__lane4_strm1_cntl        = 'd0         ;
    std__pe52__lane4_strm1_data        = 'h1234_5678 ;
    std__pe52__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe52__lane5_strm0_cntl        = 'd0         ;
    std__pe52__lane5_strm0_data        = 'h1234_5678 ;
    std__pe52__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe52__lane5_strm1_cntl        = 'd0         ;
    std__pe52__lane5_strm1_data        = 'h1234_5678 ;
    std__pe52__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe52__lane6_strm0_cntl        = 'd0         ;
    std__pe52__lane6_strm0_data        = 'h1234_5678 ;
    std__pe52__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe52__lane6_strm1_cntl        = 'd0         ;
    std__pe52__lane6_strm1_data        = 'h1234_5678 ;
    std__pe52__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe52__lane7_strm0_cntl        = 'd0         ;
    std__pe52__lane7_strm0_data        = 'h1234_5678 ;
    std__pe52__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe52__lane7_strm1_cntl        = 'd0         ;
    std__pe52__lane7_strm1_data        = 'h1234_5678 ;
    std__pe52__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe52__lane8_strm0_cntl        = 'd0         ;
    std__pe52__lane8_strm0_data        = 'h1234_5678 ;
    std__pe52__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe52__lane8_strm1_cntl        = 'd0         ;
    std__pe52__lane8_strm1_data        = 'h1234_5678 ;
    std__pe52__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe52__lane9_strm0_cntl        = 'd0         ;
    std__pe52__lane9_strm0_data        = 'h1234_5678 ;
    std__pe52__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe52__lane9_strm1_cntl        = 'd0         ;
    std__pe52__lane9_strm1_data        = 'h1234_5678 ;
    std__pe52__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe52__lane10_strm0_cntl        = 'd0         ;
    std__pe52__lane10_strm0_data        = 'h1234_5678 ;
    std__pe52__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe52__lane10_strm1_cntl        = 'd0         ;
    std__pe52__lane10_strm1_data        = 'h1234_5678 ;
    std__pe52__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe52__lane11_strm0_cntl        = 'd0         ;
    std__pe52__lane11_strm0_data        = 'h1234_5678 ;
    std__pe52__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe52__lane11_strm1_cntl        = 'd0         ;
    std__pe52__lane11_strm1_data        = 'h1234_5678 ;
    std__pe52__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe52__lane12_strm0_cntl        = 'd0         ;
    std__pe52__lane12_strm0_data        = 'h1234_5678 ;
    std__pe52__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe52__lane12_strm1_cntl        = 'd0         ;
    std__pe52__lane12_strm1_data        = 'h1234_5678 ;
    std__pe52__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe52__lane13_strm0_cntl        = 'd0         ;
    std__pe52__lane13_strm0_data        = 'h1234_5678 ;
    std__pe52__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe52__lane13_strm1_cntl        = 'd0         ;
    std__pe52__lane13_strm1_data        = 'h1234_5678 ;
    std__pe52__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe52__lane14_strm0_cntl        = 'd0         ;
    std__pe52__lane14_strm0_data        = 'h1234_5678 ;
    std__pe52__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe52__lane14_strm1_cntl        = 'd0         ;
    std__pe52__lane14_strm1_data        = 'h1234_5678 ;
    std__pe52__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe52__lane15_strm0_cntl        = 'd0         ;
    std__pe52__lane15_strm0_data        = 'h1234_5678 ;
    std__pe52__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe52__lane15_strm1_cntl        = 'd0         ;
    std__pe52__lane15_strm1_data        = 'h1234_5678 ;
    std__pe52__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe52__lane16_strm0_cntl        = 'd0         ;
    std__pe52__lane16_strm0_data        = 'h1234_5678 ;
    std__pe52__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe52__lane16_strm1_cntl        = 'd0         ;
    std__pe52__lane16_strm1_data        = 'h1234_5678 ;
    std__pe52__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe52__lane17_strm0_cntl        = 'd0         ;
    std__pe52__lane17_strm0_data        = 'h1234_5678 ;
    std__pe52__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe52__lane17_strm1_cntl        = 'd0         ;
    std__pe52__lane17_strm1_data        = 'h1234_5678 ;
    std__pe52__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe52__lane18_strm0_cntl        = 'd0         ;
    std__pe52__lane18_strm0_data        = 'h1234_5678 ;
    std__pe52__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe52__lane18_strm1_cntl        = 'd0         ;
    std__pe52__lane18_strm1_data        = 'h1234_5678 ;
    std__pe52__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe52__lane19_strm0_cntl        = 'd0         ;
    std__pe52__lane19_strm0_data        = 'h1234_5678 ;
    std__pe52__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe52__lane19_strm1_cntl        = 'd0         ;
    std__pe52__lane19_strm1_data        = 'h1234_5678 ;
    std__pe52__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe52__lane20_strm0_cntl        = 'd0         ;
    std__pe52__lane20_strm0_data        = 'h1234_5678 ;
    std__pe52__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe52__lane20_strm1_cntl        = 'd0         ;
    std__pe52__lane20_strm1_data        = 'h1234_5678 ;
    std__pe52__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe52__lane21_strm0_cntl        = 'd0         ;
    std__pe52__lane21_strm0_data        = 'h1234_5678 ;
    std__pe52__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe52__lane21_strm1_cntl        = 'd0         ;
    std__pe52__lane21_strm1_data        = 'h1234_5678 ;
    std__pe52__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe52__lane22_strm0_cntl        = 'd0         ;
    std__pe52__lane22_strm0_data        = 'h1234_5678 ;
    std__pe52__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe52__lane22_strm1_cntl        = 'd0         ;
    std__pe52__lane22_strm1_data        = 'h1234_5678 ;
    std__pe52__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe52__lane23_strm0_cntl        = 'd0         ;
    std__pe52__lane23_strm0_data        = 'h1234_5678 ;
    std__pe52__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe52__lane23_strm1_cntl        = 'd0         ;
    std__pe52__lane23_strm1_data        = 'h1234_5678 ;
    std__pe52__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe52__lane24_strm0_cntl        = 'd0         ;
    std__pe52__lane24_strm0_data        = 'h1234_5678 ;
    std__pe52__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe52__lane24_strm1_cntl        = 'd0         ;
    std__pe52__lane24_strm1_data        = 'h1234_5678 ;
    std__pe52__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe52__lane25_strm0_cntl        = 'd0         ;
    std__pe52__lane25_strm0_data        = 'h1234_5678 ;
    std__pe52__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe52__lane25_strm1_cntl        = 'd0         ;
    std__pe52__lane25_strm1_data        = 'h1234_5678 ;
    std__pe52__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe52__lane26_strm0_cntl        = 'd0         ;
    std__pe52__lane26_strm0_data        = 'h1234_5678 ;
    std__pe52__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe52__lane26_strm1_cntl        = 'd0         ;
    std__pe52__lane26_strm1_data        = 'h1234_5678 ;
    std__pe52__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe52__lane27_strm0_cntl        = 'd0         ;
    std__pe52__lane27_strm0_data        = 'h1234_5678 ;
    std__pe52__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe52__lane27_strm1_cntl        = 'd0         ;
    std__pe52__lane27_strm1_data        = 'h1234_5678 ;
    std__pe52__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe52__lane28_strm0_cntl        = 'd0         ;
    std__pe52__lane28_strm0_data        = 'h1234_5678 ;
    std__pe52__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe52__lane28_strm1_cntl        = 'd0         ;
    std__pe52__lane28_strm1_data        = 'h1234_5678 ;
    std__pe52__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe52__lane29_strm0_cntl        = 'd0         ;
    std__pe52__lane29_strm0_data        = 'h1234_5678 ;
    std__pe52__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe52__lane29_strm1_cntl        = 'd0         ;
    std__pe52__lane29_strm1_data        = 'h1234_5678 ;
    std__pe52__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe52__lane30_strm0_cntl        = 'd0         ;
    std__pe52__lane30_strm0_data        = 'h1234_5678 ;
    std__pe52__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe52__lane30_strm1_cntl        = 'd0         ;
    std__pe52__lane30_strm1_data        = 'h1234_5678 ;
    std__pe52__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe52__lane31_strm0_cntl        = 'd0         ;
    std__pe52__lane31_strm0_data        = 'h1234_5678 ;
    std__pe52__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe52__lane31_strm1_cntl        = 'd0         ;
    std__pe52__lane31_strm1_data        = 'h1234_5678 ;
    std__pe52__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe53__lane0_strm0_cntl        = 'd0         ;
    std__pe53__lane0_strm0_data        = 'h1234_5678 ;
    std__pe53__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe53__lane0_strm1_cntl        = 'd0         ;
    std__pe53__lane0_strm1_data        = 'h1234_5678 ;
    std__pe53__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe53__lane1_strm0_cntl        = 'd0         ;
    std__pe53__lane1_strm0_data        = 'h1234_5678 ;
    std__pe53__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe53__lane1_strm1_cntl        = 'd0         ;
    std__pe53__lane1_strm1_data        = 'h1234_5678 ;
    std__pe53__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe53__lane2_strm0_cntl        = 'd0         ;
    std__pe53__lane2_strm0_data        = 'h1234_5678 ;
    std__pe53__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe53__lane2_strm1_cntl        = 'd0         ;
    std__pe53__lane2_strm1_data        = 'h1234_5678 ;
    std__pe53__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe53__lane3_strm0_cntl        = 'd0         ;
    std__pe53__lane3_strm0_data        = 'h1234_5678 ;
    std__pe53__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe53__lane3_strm1_cntl        = 'd0         ;
    std__pe53__lane3_strm1_data        = 'h1234_5678 ;
    std__pe53__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe53__lane4_strm0_cntl        = 'd0         ;
    std__pe53__lane4_strm0_data        = 'h1234_5678 ;
    std__pe53__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe53__lane4_strm1_cntl        = 'd0         ;
    std__pe53__lane4_strm1_data        = 'h1234_5678 ;
    std__pe53__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe53__lane5_strm0_cntl        = 'd0         ;
    std__pe53__lane5_strm0_data        = 'h1234_5678 ;
    std__pe53__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe53__lane5_strm1_cntl        = 'd0         ;
    std__pe53__lane5_strm1_data        = 'h1234_5678 ;
    std__pe53__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe53__lane6_strm0_cntl        = 'd0         ;
    std__pe53__lane6_strm0_data        = 'h1234_5678 ;
    std__pe53__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe53__lane6_strm1_cntl        = 'd0         ;
    std__pe53__lane6_strm1_data        = 'h1234_5678 ;
    std__pe53__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe53__lane7_strm0_cntl        = 'd0         ;
    std__pe53__lane7_strm0_data        = 'h1234_5678 ;
    std__pe53__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe53__lane7_strm1_cntl        = 'd0         ;
    std__pe53__lane7_strm1_data        = 'h1234_5678 ;
    std__pe53__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe53__lane8_strm0_cntl        = 'd0         ;
    std__pe53__lane8_strm0_data        = 'h1234_5678 ;
    std__pe53__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe53__lane8_strm1_cntl        = 'd0         ;
    std__pe53__lane8_strm1_data        = 'h1234_5678 ;
    std__pe53__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe53__lane9_strm0_cntl        = 'd0         ;
    std__pe53__lane9_strm0_data        = 'h1234_5678 ;
    std__pe53__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe53__lane9_strm1_cntl        = 'd0         ;
    std__pe53__lane9_strm1_data        = 'h1234_5678 ;
    std__pe53__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe53__lane10_strm0_cntl        = 'd0         ;
    std__pe53__lane10_strm0_data        = 'h1234_5678 ;
    std__pe53__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe53__lane10_strm1_cntl        = 'd0         ;
    std__pe53__lane10_strm1_data        = 'h1234_5678 ;
    std__pe53__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe53__lane11_strm0_cntl        = 'd0         ;
    std__pe53__lane11_strm0_data        = 'h1234_5678 ;
    std__pe53__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe53__lane11_strm1_cntl        = 'd0         ;
    std__pe53__lane11_strm1_data        = 'h1234_5678 ;
    std__pe53__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe53__lane12_strm0_cntl        = 'd0         ;
    std__pe53__lane12_strm0_data        = 'h1234_5678 ;
    std__pe53__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe53__lane12_strm1_cntl        = 'd0         ;
    std__pe53__lane12_strm1_data        = 'h1234_5678 ;
    std__pe53__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe53__lane13_strm0_cntl        = 'd0         ;
    std__pe53__lane13_strm0_data        = 'h1234_5678 ;
    std__pe53__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe53__lane13_strm1_cntl        = 'd0         ;
    std__pe53__lane13_strm1_data        = 'h1234_5678 ;
    std__pe53__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe53__lane14_strm0_cntl        = 'd0         ;
    std__pe53__lane14_strm0_data        = 'h1234_5678 ;
    std__pe53__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe53__lane14_strm1_cntl        = 'd0         ;
    std__pe53__lane14_strm1_data        = 'h1234_5678 ;
    std__pe53__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe53__lane15_strm0_cntl        = 'd0         ;
    std__pe53__lane15_strm0_data        = 'h1234_5678 ;
    std__pe53__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe53__lane15_strm1_cntl        = 'd0         ;
    std__pe53__lane15_strm1_data        = 'h1234_5678 ;
    std__pe53__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe53__lane16_strm0_cntl        = 'd0         ;
    std__pe53__lane16_strm0_data        = 'h1234_5678 ;
    std__pe53__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe53__lane16_strm1_cntl        = 'd0         ;
    std__pe53__lane16_strm1_data        = 'h1234_5678 ;
    std__pe53__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe53__lane17_strm0_cntl        = 'd0         ;
    std__pe53__lane17_strm0_data        = 'h1234_5678 ;
    std__pe53__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe53__lane17_strm1_cntl        = 'd0         ;
    std__pe53__lane17_strm1_data        = 'h1234_5678 ;
    std__pe53__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe53__lane18_strm0_cntl        = 'd0         ;
    std__pe53__lane18_strm0_data        = 'h1234_5678 ;
    std__pe53__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe53__lane18_strm1_cntl        = 'd0         ;
    std__pe53__lane18_strm1_data        = 'h1234_5678 ;
    std__pe53__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe53__lane19_strm0_cntl        = 'd0         ;
    std__pe53__lane19_strm0_data        = 'h1234_5678 ;
    std__pe53__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe53__lane19_strm1_cntl        = 'd0         ;
    std__pe53__lane19_strm1_data        = 'h1234_5678 ;
    std__pe53__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe53__lane20_strm0_cntl        = 'd0         ;
    std__pe53__lane20_strm0_data        = 'h1234_5678 ;
    std__pe53__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe53__lane20_strm1_cntl        = 'd0         ;
    std__pe53__lane20_strm1_data        = 'h1234_5678 ;
    std__pe53__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe53__lane21_strm0_cntl        = 'd0         ;
    std__pe53__lane21_strm0_data        = 'h1234_5678 ;
    std__pe53__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe53__lane21_strm1_cntl        = 'd0         ;
    std__pe53__lane21_strm1_data        = 'h1234_5678 ;
    std__pe53__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe53__lane22_strm0_cntl        = 'd0         ;
    std__pe53__lane22_strm0_data        = 'h1234_5678 ;
    std__pe53__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe53__lane22_strm1_cntl        = 'd0         ;
    std__pe53__lane22_strm1_data        = 'h1234_5678 ;
    std__pe53__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe53__lane23_strm0_cntl        = 'd0         ;
    std__pe53__lane23_strm0_data        = 'h1234_5678 ;
    std__pe53__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe53__lane23_strm1_cntl        = 'd0         ;
    std__pe53__lane23_strm1_data        = 'h1234_5678 ;
    std__pe53__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe53__lane24_strm0_cntl        = 'd0         ;
    std__pe53__lane24_strm0_data        = 'h1234_5678 ;
    std__pe53__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe53__lane24_strm1_cntl        = 'd0         ;
    std__pe53__lane24_strm1_data        = 'h1234_5678 ;
    std__pe53__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe53__lane25_strm0_cntl        = 'd0         ;
    std__pe53__lane25_strm0_data        = 'h1234_5678 ;
    std__pe53__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe53__lane25_strm1_cntl        = 'd0         ;
    std__pe53__lane25_strm1_data        = 'h1234_5678 ;
    std__pe53__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe53__lane26_strm0_cntl        = 'd0         ;
    std__pe53__lane26_strm0_data        = 'h1234_5678 ;
    std__pe53__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe53__lane26_strm1_cntl        = 'd0         ;
    std__pe53__lane26_strm1_data        = 'h1234_5678 ;
    std__pe53__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe53__lane27_strm0_cntl        = 'd0         ;
    std__pe53__lane27_strm0_data        = 'h1234_5678 ;
    std__pe53__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe53__lane27_strm1_cntl        = 'd0         ;
    std__pe53__lane27_strm1_data        = 'h1234_5678 ;
    std__pe53__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe53__lane28_strm0_cntl        = 'd0         ;
    std__pe53__lane28_strm0_data        = 'h1234_5678 ;
    std__pe53__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe53__lane28_strm1_cntl        = 'd0         ;
    std__pe53__lane28_strm1_data        = 'h1234_5678 ;
    std__pe53__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe53__lane29_strm0_cntl        = 'd0         ;
    std__pe53__lane29_strm0_data        = 'h1234_5678 ;
    std__pe53__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe53__lane29_strm1_cntl        = 'd0         ;
    std__pe53__lane29_strm1_data        = 'h1234_5678 ;
    std__pe53__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe53__lane30_strm0_cntl        = 'd0         ;
    std__pe53__lane30_strm0_data        = 'h1234_5678 ;
    std__pe53__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe53__lane30_strm1_cntl        = 'd0         ;
    std__pe53__lane30_strm1_data        = 'h1234_5678 ;
    std__pe53__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe53__lane31_strm0_cntl        = 'd0         ;
    std__pe53__lane31_strm0_data        = 'h1234_5678 ;
    std__pe53__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe53__lane31_strm1_cntl        = 'd0         ;
    std__pe53__lane31_strm1_data        = 'h1234_5678 ;
    std__pe53__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe54__lane0_strm0_cntl        = 'd0         ;
    std__pe54__lane0_strm0_data        = 'h1234_5678 ;
    std__pe54__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe54__lane0_strm1_cntl        = 'd0         ;
    std__pe54__lane0_strm1_data        = 'h1234_5678 ;
    std__pe54__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe54__lane1_strm0_cntl        = 'd0         ;
    std__pe54__lane1_strm0_data        = 'h1234_5678 ;
    std__pe54__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe54__lane1_strm1_cntl        = 'd0         ;
    std__pe54__lane1_strm1_data        = 'h1234_5678 ;
    std__pe54__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe54__lane2_strm0_cntl        = 'd0         ;
    std__pe54__lane2_strm0_data        = 'h1234_5678 ;
    std__pe54__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe54__lane2_strm1_cntl        = 'd0         ;
    std__pe54__lane2_strm1_data        = 'h1234_5678 ;
    std__pe54__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe54__lane3_strm0_cntl        = 'd0         ;
    std__pe54__lane3_strm0_data        = 'h1234_5678 ;
    std__pe54__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe54__lane3_strm1_cntl        = 'd0         ;
    std__pe54__lane3_strm1_data        = 'h1234_5678 ;
    std__pe54__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe54__lane4_strm0_cntl        = 'd0         ;
    std__pe54__lane4_strm0_data        = 'h1234_5678 ;
    std__pe54__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe54__lane4_strm1_cntl        = 'd0         ;
    std__pe54__lane4_strm1_data        = 'h1234_5678 ;
    std__pe54__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe54__lane5_strm0_cntl        = 'd0         ;
    std__pe54__lane5_strm0_data        = 'h1234_5678 ;
    std__pe54__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe54__lane5_strm1_cntl        = 'd0         ;
    std__pe54__lane5_strm1_data        = 'h1234_5678 ;
    std__pe54__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe54__lane6_strm0_cntl        = 'd0         ;
    std__pe54__lane6_strm0_data        = 'h1234_5678 ;
    std__pe54__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe54__lane6_strm1_cntl        = 'd0         ;
    std__pe54__lane6_strm1_data        = 'h1234_5678 ;
    std__pe54__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe54__lane7_strm0_cntl        = 'd0         ;
    std__pe54__lane7_strm0_data        = 'h1234_5678 ;
    std__pe54__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe54__lane7_strm1_cntl        = 'd0         ;
    std__pe54__lane7_strm1_data        = 'h1234_5678 ;
    std__pe54__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe54__lane8_strm0_cntl        = 'd0         ;
    std__pe54__lane8_strm0_data        = 'h1234_5678 ;
    std__pe54__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe54__lane8_strm1_cntl        = 'd0         ;
    std__pe54__lane8_strm1_data        = 'h1234_5678 ;
    std__pe54__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe54__lane9_strm0_cntl        = 'd0         ;
    std__pe54__lane9_strm0_data        = 'h1234_5678 ;
    std__pe54__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe54__lane9_strm1_cntl        = 'd0         ;
    std__pe54__lane9_strm1_data        = 'h1234_5678 ;
    std__pe54__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe54__lane10_strm0_cntl        = 'd0         ;
    std__pe54__lane10_strm0_data        = 'h1234_5678 ;
    std__pe54__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe54__lane10_strm1_cntl        = 'd0         ;
    std__pe54__lane10_strm1_data        = 'h1234_5678 ;
    std__pe54__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe54__lane11_strm0_cntl        = 'd0         ;
    std__pe54__lane11_strm0_data        = 'h1234_5678 ;
    std__pe54__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe54__lane11_strm1_cntl        = 'd0         ;
    std__pe54__lane11_strm1_data        = 'h1234_5678 ;
    std__pe54__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe54__lane12_strm0_cntl        = 'd0         ;
    std__pe54__lane12_strm0_data        = 'h1234_5678 ;
    std__pe54__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe54__lane12_strm1_cntl        = 'd0         ;
    std__pe54__lane12_strm1_data        = 'h1234_5678 ;
    std__pe54__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe54__lane13_strm0_cntl        = 'd0         ;
    std__pe54__lane13_strm0_data        = 'h1234_5678 ;
    std__pe54__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe54__lane13_strm1_cntl        = 'd0         ;
    std__pe54__lane13_strm1_data        = 'h1234_5678 ;
    std__pe54__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe54__lane14_strm0_cntl        = 'd0         ;
    std__pe54__lane14_strm0_data        = 'h1234_5678 ;
    std__pe54__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe54__lane14_strm1_cntl        = 'd0         ;
    std__pe54__lane14_strm1_data        = 'h1234_5678 ;
    std__pe54__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe54__lane15_strm0_cntl        = 'd0         ;
    std__pe54__lane15_strm0_data        = 'h1234_5678 ;
    std__pe54__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe54__lane15_strm1_cntl        = 'd0         ;
    std__pe54__lane15_strm1_data        = 'h1234_5678 ;
    std__pe54__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe54__lane16_strm0_cntl        = 'd0         ;
    std__pe54__lane16_strm0_data        = 'h1234_5678 ;
    std__pe54__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe54__lane16_strm1_cntl        = 'd0         ;
    std__pe54__lane16_strm1_data        = 'h1234_5678 ;
    std__pe54__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe54__lane17_strm0_cntl        = 'd0         ;
    std__pe54__lane17_strm0_data        = 'h1234_5678 ;
    std__pe54__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe54__lane17_strm1_cntl        = 'd0         ;
    std__pe54__lane17_strm1_data        = 'h1234_5678 ;
    std__pe54__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe54__lane18_strm0_cntl        = 'd0         ;
    std__pe54__lane18_strm0_data        = 'h1234_5678 ;
    std__pe54__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe54__lane18_strm1_cntl        = 'd0         ;
    std__pe54__lane18_strm1_data        = 'h1234_5678 ;
    std__pe54__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe54__lane19_strm0_cntl        = 'd0         ;
    std__pe54__lane19_strm0_data        = 'h1234_5678 ;
    std__pe54__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe54__lane19_strm1_cntl        = 'd0         ;
    std__pe54__lane19_strm1_data        = 'h1234_5678 ;
    std__pe54__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe54__lane20_strm0_cntl        = 'd0         ;
    std__pe54__lane20_strm0_data        = 'h1234_5678 ;
    std__pe54__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe54__lane20_strm1_cntl        = 'd0         ;
    std__pe54__lane20_strm1_data        = 'h1234_5678 ;
    std__pe54__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe54__lane21_strm0_cntl        = 'd0         ;
    std__pe54__lane21_strm0_data        = 'h1234_5678 ;
    std__pe54__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe54__lane21_strm1_cntl        = 'd0         ;
    std__pe54__lane21_strm1_data        = 'h1234_5678 ;
    std__pe54__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe54__lane22_strm0_cntl        = 'd0         ;
    std__pe54__lane22_strm0_data        = 'h1234_5678 ;
    std__pe54__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe54__lane22_strm1_cntl        = 'd0         ;
    std__pe54__lane22_strm1_data        = 'h1234_5678 ;
    std__pe54__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe54__lane23_strm0_cntl        = 'd0         ;
    std__pe54__lane23_strm0_data        = 'h1234_5678 ;
    std__pe54__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe54__lane23_strm1_cntl        = 'd0         ;
    std__pe54__lane23_strm1_data        = 'h1234_5678 ;
    std__pe54__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe54__lane24_strm0_cntl        = 'd0         ;
    std__pe54__lane24_strm0_data        = 'h1234_5678 ;
    std__pe54__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe54__lane24_strm1_cntl        = 'd0         ;
    std__pe54__lane24_strm1_data        = 'h1234_5678 ;
    std__pe54__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe54__lane25_strm0_cntl        = 'd0         ;
    std__pe54__lane25_strm0_data        = 'h1234_5678 ;
    std__pe54__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe54__lane25_strm1_cntl        = 'd0         ;
    std__pe54__lane25_strm1_data        = 'h1234_5678 ;
    std__pe54__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe54__lane26_strm0_cntl        = 'd0         ;
    std__pe54__lane26_strm0_data        = 'h1234_5678 ;
    std__pe54__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe54__lane26_strm1_cntl        = 'd0         ;
    std__pe54__lane26_strm1_data        = 'h1234_5678 ;
    std__pe54__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe54__lane27_strm0_cntl        = 'd0         ;
    std__pe54__lane27_strm0_data        = 'h1234_5678 ;
    std__pe54__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe54__lane27_strm1_cntl        = 'd0         ;
    std__pe54__lane27_strm1_data        = 'h1234_5678 ;
    std__pe54__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe54__lane28_strm0_cntl        = 'd0         ;
    std__pe54__lane28_strm0_data        = 'h1234_5678 ;
    std__pe54__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe54__lane28_strm1_cntl        = 'd0         ;
    std__pe54__lane28_strm1_data        = 'h1234_5678 ;
    std__pe54__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe54__lane29_strm0_cntl        = 'd0         ;
    std__pe54__lane29_strm0_data        = 'h1234_5678 ;
    std__pe54__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe54__lane29_strm1_cntl        = 'd0         ;
    std__pe54__lane29_strm1_data        = 'h1234_5678 ;
    std__pe54__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe54__lane30_strm0_cntl        = 'd0         ;
    std__pe54__lane30_strm0_data        = 'h1234_5678 ;
    std__pe54__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe54__lane30_strm1_cntl        = 'd0         ;
    std__pe54__lane30_strm1_data        = 'h1234_5678 ;
    std__pe54__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe54__lane31_strm0_cntl        = 'd0         ;
    std__pe54__lane31_strm0_data        = 'h1234_5678 ;
    std__pe54__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe54__lane31_strm1_cntl        = 'd0         ;
    std__pe54__lane31_strm1_data        = 'h1234_5678 ;
    std__pe54__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe55__lane0_strm0_cntl        = 'd0         ;
    std__pe55__lane0_strm0_data        = 'h1234_5678 ;
    std__pe55__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe55__lane0_strm1_cntl        = 'd0         ;
    std__pe55__lane0_strm1_data        = 'h1234_5678 ;
    std__pe55__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe55__lane1_strm0_cntl        = 'd0         ;
    std__pe55__lane1_strm0_data        = 'h1234_5678 ;
    std__pe55__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe55__lane1_strm1_cntl        = 'd0         ;
    std__pe55__lane1_strm1_data        = 'h1234_5678 ;
    std__pe55__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe55__lane2_strm0_cntl        = 'd0         ;
    std__pe55__lane2_strm0_data        = 'h1234_5678 ;
    std__pe55__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe55__lane2_strm1_cntl        = 'd0         ;
    std__pe55__lane2_strm1_data        = 'h1234_5678 ;
    std__pe55__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe55__lane3_strm0_cntl        = 'd0         ;
    std__pe55__lane3_strm0_data        = 'h1234_5678 ;
    std__pe55__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe55__lane3_strm1_cntl        = 'd0         ;
    std__pe55__lane3_strm1_data        = 'h1234_5678 ;
    std__pe55__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe55__lane4_strm0_cntl        = 'd0         ;
    std__pe55__lane4_strm0_data        = 'h1234_5678 ;
    std__pe55__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe55__lane4_strm1_cntl        = 'd0         ;
    std__pe55__lane4_strm1_data        = 'h1234_5678 ;
    std__pe55__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe55__lane5_strm0_cntl        = 'd0         ;
    std__pe55__lane5_strm0_data        = 'h1234_5678 ;
    std__pe55__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe55__lane5_strm1_cntl        = 'd0         ;
    std__pe55__lane5_strm1_data        = 'h1234_5678 ;
    std__pe55__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe55__lane6_strm0_cntl        = 'd0         ;
    std__pe55__lane6_strm0_data        = 'h1234_5678 ;
    std__pe55__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe55__lane6_strm1_cntl        = 'd0         ;
    std__pe55__lane6_strm1_data        = 'h1234_5678 ;
    std__pe55__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe55__lane7_strm0_cntl        = 'd0         ;
    std__pe55__lane7_strm0_data        = 'h1234_5678 ;
    std__pe55__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe55__lane7_strm1_cntl        = 'd0         ;
    std__pe55__lane7_strm1_data        = 'h1234_5678 ;
    std__pe55__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe55__lane8_strm0_cntl        = 'd0         ;
    std__pe55__lane8_strm0_data        = 'h1234_5678 ;
    std__pe55__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe55__lane8_strm1_cntl        = 'd0         ;
    std__pe55__lane8_strm1_data        = 'h1234_5678 ;
    std__pe55__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe55__lane9_strm0_cntl        = 'd0         ;
    std__pe55__lane9_strm0_data        = 'h1234_5678 ;
    std__pe55__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe55__lane9_strm1_cntl        = 'd0         ;
    std__pe55__lane9_strm1_data        = 'h1234_5678 ;
    std__pe55__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe55__lane10_strm0_cntl        = 'd0         ;
    std__pe55__lane10_strm0_data        = 'h1234_5678 ;
    std__pe55__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe55__lane10_strm1_cntl        = 'd0         ;
    std__pe55__lane10_strm1_data        = 'h1234_5678 ;
    std__pe55__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe55__lane11_strm0_cntl        = 'd0         ;
    std__pe55__lane11_strm0_data        = 'h1234_5678 ;
    std__pe55__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe55__lane11_strm1_cntl        = 'd0         ;
    std__pe55__lane11_strm1_data        = 'h1234_5678 ;
    std__pe55__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe55__lane12_strm0_cntl        = 'd0         ;
    std__pe55__lane12_strm0_data        = 'h1234_5678 ;
    std__pe55__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe55__lane12_strm1_cntl        = 'd0         ;
    std__pe55__lane12_strm1_data        = 'h1234_5678 ;
    std__pe55__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe55__lane13_strm0_cntl        = 'd0         ;
    std__pe55__lane13_strm0_data        = 'h1234_5678 ;
    std__pe55__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe55__lane13_strm1_cntl        = 'd0         ;
    std__pe55__lane13_strm1_data        = 'h1234_5678 ;
    std__pe55__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe55__lane14_strm0_cntl        = 'd0         ;
    std__pe55__lane14_strm0_data        = 'h1234_5678 ;
    std__pe55__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe55__lane14_strm1_cntl        = 'd0         ;
    std__pe55__lane14_strm1_data        = 'h1234_5678 ;
    std__pe55__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe55__lane15_strm0_cntl        = 'd0         ;
    std__pe55__lane15_strm0_data        = 'h1234_5678 ;
    std__pe55__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe55__lane15_strm1_cntl        = 'd0         ;
    std__pe55__lane15_strm1_data        = 'h1234_5678 ;
    std__pe55__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe55__lane16_strm0_cntl        = 'd0         ;
    std__pe55__lane16_strm0_data        = 'h1234_5678 ;
    std__pe55__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe55__lane16_strm1_cntl        = 'd0         ;
    std__pe55__lane16_strm1_data        = 'h1234_5678 ;
    std__pe55__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe55__lane17_strm0_cntl        = 'd0         ;
    std__pe55__lane17_strm0_data        = 'h1234_5678 ;
    std__pe55__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe55__lane17_strm1_cntl        = 'd0         ;
    std__pe55__lane17_strm1_data        = 'h1234_5678 ;
    std__pe55__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe55__lane18_strm0_cntl        = 'd0         ;
    std__pe55__lane18_strm0_data        = 'h1234_5678 ;
    std__pe55__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe55__lane18_strm1_cntl        = 'd0         ;
    std__pe55__lane18_strm1_data        = 'h1234_5678 ;
    std__pe55__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe55__lane19_strm0_cntl        = 'd0         ;
    std__pe55__lane19_strm0_data        = 'h1234_5678 ;
    std__pe55__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe55__lane19_strm1_cntl        = 'd0         ;
    std__pe55__lane19_strm1_data        = 'h1234_5678 ;
    std__pe55__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe55__lane20_strm0_cntl        = 'd0         ;
    std__pe55__lane20_strm0_data        = 'h1234_5678 ;
    std__pe55__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe55__lane20_strm1_cntl        = 'd0         ;
    std__pe55__lane20_strm1_data        = 'h1234_5678 ;
    std__pe55__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe55__lane21_strm0_cntl        = 'd0         ;
    std__pe55__lane21_strm0_data        = 'h1234_5678 ;
    std__pe55__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe55__lane21_strm1_cntl        = 'd0         ;
    std__pe55__lane21_strm1_data        = 'h1234_5678 ;
    std__pe55__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe55__lane22_strm0_cntl        = 'd0         ;
    std__pe55__lane22_strm0_data        = 'h1234_5678 ;
    std__pe55__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe55__lane22_strm1_cntl        = 'd0         ;
    std__pe55__lane22_strm1_data        = 'h1234_5678 ;
    std__pe55__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe55__lane23_strm0_cntl        = 'd0         ;
    std__pe55__lane23_strm0_data        = 'h1234_5678 ;
    std__pe55__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe55__lane23_strm1_cntl        = 'd0         ;
    std__pe55__lane23_strm1_data        = 'h1234_5678 ;
    std__pe55__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe55__lane24_strm0_cntl        = 'd0         ;
    std__pe55__lane24_strm0_data        = 'h1234_5678 ;
    std__pe55__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe55__lane24_strm1_cntl        = 'd0         ;
    std__pe55__lane24_strm1_data        = 'h1234_5678 ;
    std__pe55__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe55__lane25_strm0_cntl        = 'd0         ;
    std__pe55__lane25_strm0_data        = 'h1234_5678 ;
    std__pe55__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe55__lane25_strm1_cntl        = 'd0         ;
    std__pe55__lane25_strm1_data        = 'h1234_5678 ;
    std__pe55__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe55__lane26_strm0_cntl        = 'd0         ;
    std__pe55__lane26_strm0_data        = 'h1234_5678 ;
    std__pe55__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe55__lane26_strm1_cntl        = 'd0         ;
    std__pe55__lane26_strm1_data        = 'h1234_5678 ;
    std__pe55__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe55__lane27_strm0_cntl        = 'd0         ;
    std__pe55__lane27_strm0_data        = 'h1234_5678 ;
    std__pe55__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe55__lane27_strm1_cntl        = 'd0         ;
    std__pe55__lane27_strm1_data        = 'h1234_5678 ;
    std__pe55__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe55__lane28_strm0_cntl        = 'd0         ;
    std__pe55__lane28_strm0_data        = 'h1234_5678 ;
    std__pe55__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe55__lane28_strm1_cntl        = 'd0         ;
    std__pe55__lane28_strm1_data        = 'h1234_5678 ;
    std__pe55__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe55__lane29_strm0_cntl        = 'd0         ;
    std__pe55__lane29_strm0_data        = 'h1234_5678 ;
    std__pe55__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe55__lane29_strm1_cntl        = 'd0         ;
    std__pe55__lane29_strm1_data        = 'h1234_5678 ;
    std__pe55__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe55__lane30_strm0_cntl        = 'd0         ;
    std__pe55__lane30_strm0_data        = 'h1234_5678 ;
    std__pe55__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe55__lane30_strm1_cntl        = 'd0         ;
    std__pe55__lane30_strm1_data        = 'h1234_5678 ;
    std__pe55__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe55__lane31_strm0_cntl        = 'd0         ;
    std__pe55__lane31_strm0_data        = 'h1234_5678 ;
    std__pe55__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe55__lane31_strm1_cntl        = 'd0         ;
    std__pe55__lane31_strm1_data        = 'h1234_5678 ;
    std__pe55__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe56__lane0_strm0_cntl        = 'd0         ;
    std__pe56__lane0_strm0_data        = 'h1234_5678 ;
    std__pe56__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe56__lane0_strm1_cntl        = 'd0         ;
    std__pe56__lane0_strm1_data        = 'h1234_5678 ;
    std__pe56__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe56__lane1_strm0_cntl        = 'd0         ;
    std__pe56__lane1_strm0_data        = 'h1234_5678 ;
    std__pe56__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe56__lane1_strm1_cntl        = 'd0         ;
    std__pe56__lane1_strm1_data        = 'h1234_5678 ;
    std__pe56__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe56__lane2_strm0_cntl        = 'd0         ;
    std__pe56__lane2_strm0_data        = 'h1234_5678 ;
    std__pe56__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe56__lane2_strm1_cntl        = 'd0         ;
    std__pe56__lane2_strm1_data        = 'h1234_5678 ;
    std__pe56__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe56__lane3_strm0_cntl        = 'd0         ;
    std__pe56__lane3_strm0_data        = 'h1234_5678 ;
    std__pe56__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe56__lane3_strm1_cntl        = 'd0         ;
    std__pe56__lane3_strm1_data        = 'h1234_5678 ;
    std__pe56__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe56__lane4_strm0_cntl        = 'd0         ;
    std__pe56__lane4_strm0_data        = 'h1234_5678 ;
    std__pe56__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe56__lane4_strm1_cntl        = 'd0         ;
    std__pe56__lane4_strm1_data        = 'h1234_5678 ;
    std__pe56__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe56__lane5_strm0_cntl        = 'd0         ;
    std__pe56__lane5_strm0_data        = 'h1234_5678 ;
    std__pe56__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe56__lane5_strm1_cntl        = 'd0         ;
    std__pe56__lane5_strm1_data        = 'h1234_5678 ;
    std__pe56__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe56__lane6_strm0_cntl        = 'd0         ;
    std__pe56__lane6_strm0_data        = 'h1234_5678 ;
    std__pe56__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe56__lane6_strm1_cntl        = 'd0         ;
    std__pe56__lane6_strm1_data        = 'h1234_5678 ;
    std__pe56__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe56__lane7_strm0_cntl        = 'd0         ;
    std__pe56__lane7_strm0_data        = 'h1234_5678 ;
    std__pe56__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe56__lane7_strm1_cntl        = 'd0         ;
    std__pe56__lane7_strm1_data        = 'h1234_5678 ;
    std__pe56__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe56__lane8_strm0_cntl        = 'd0         ;
    std__pe56__lane8_strm0_data        = 'h1234_5678 ;
    std__pe56__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe56__lane8_strm1_cntl        = 'd0         ;
    std__pe56__lane8_strm1_data        = 'h1234_5678 ;
    std__pe56__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe56__lane9_strm0_cntl        = 'd0         ;
    std__pe56__lane9_strm0_data        = 'h1234_5678 ;
    std__pe56__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe56__lane9_strm1_cntl        = 'd0         ;
    std__pe56__lane9_strm1_data        = 'h1234_5678 ;
    std__pe56__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe56__lane10_strm0_cntl        = 'd0         ;
    std__pe56__lane10_strm0_data        = 'h1234_5678 ;
    std__pe56__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe56__lane10_strm1_cntl        = 'd0         ;
    std__pe56__lane10_strm1_data        = 'h1234_5678 ;
    std__pe56__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe56__lane11_strm0_cntl        = 'd0         ;
    std__pe56__lane11_strm0_data        = 'h1234_5678 ;
    std__pe56__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe56__lane11_strm1_cntl        = 'd0         ;
    std__pe56__lane11_strm1_data        = 'h1234_5678 ;
    std__pe56__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe56__lane12_strm0_cntl        = 'd0         ;
    std__pe56__lane12_strm0_data        = 'h1234_5678 ;
    std__pe56__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe56__lane12_strm1_cntl        = 'd0         ;
    std__pe56__lane12_strm1_data        = 'h1234_5678 ;
    std__pe56__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe56__lane13_strm0_cntl        = 'd0         ;
    std__pe56__lane13_strm0_data        = 'h1234_5678 ;
    std__pe56__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe56__lane13_strm1_cntl        = 'd0         ;
    std__pe56__lane13_strm1_data        = 'h1234_5678 ;
    std__pe56__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe56__lane14_strm0_cntl        = 'd0         ;
    std__pe56__lane14_strm0_data        = 'h1234_5678 ;
    std__pe56__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe56__lane14_strm1_cntl        = 'd0         ;
    std__pe56__lane14_strm1_data        = 'h1234_5678 ;
    std__pe56__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe56__lane15_strm0_cntl        = 'd0         ;
    std__pe56__lane15_strm0_data        = 'h1234_5678 ;
    std__pe56__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe56__lane15_strm1_cntl        = 'd0         ;
    std__pe56__lane15_strm1_data        = 'h1234_5678 ;
    std__pe56__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe56__lane16_strm0_cntl        = 'd0         ;
    std__pe56__lane16_strm0_data        = 'h1234_5678 ;
    std__pe56__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe56__lane16_strm1_cntl        = 'd0         ;
    std__pe56__lane16_strm1_data        = 'h1234_5678 ;
    std__pe56__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe56__lane17_strm0_cntl        = 'd0         ;
    std__pe56__lane17_strm0_data        = 'h1234_5678 ;
    std__pe56__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe56__lane17_strm1_cntl        = 'd0         ;
    std__pe56__lane17_strm1_data        = 'h1234_5678 ;
    std__pe56__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe56__lane18_strm0_cntl        = 'd0         ;
    std__pe56__lane18_strm0_data        = 'h1234_5678 ;
    std__pe56__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe56__lane18_strm1_cntl        = 'd0         ;
    std__pe56__lane18_strm1_data        = 'h1234_5678 ;
    std__pe56__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe56__lane19_strm0_cntl        = 'd0         ;
    std__pe56__lane19_strm0_data        = 'h1234_5678 ;
    std__pe56__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe56__lane19_strm1_cntl        = 'd0         ;
    std__pe56__lane19_strm1_data        = 'h1234_5678 ;
    std__pe56__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe56__lane20_strm0_cntl        = 'd0         ;
    std__pe56__lane20_strm0_data        = 'h1234_5678 ;
    std__pe56__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe56__lane20_strm1_cntl        = 'd0         ;
    std__pe56__lane20_strm1_data        = 'h1234_5678 ;
    std__pe56__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe56__lane21_strm0_cntl        = 'd0         ;
    std__pe56__lane21_strm0_data        = 'h1234_5678 ;
    std__pe56__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe56__lane21_strm1_cntl        = 'd0         ;
    std__pe56__lane21_strm1_data        = 'h1234_5678 ;
    std__pe56__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe56__lane22_strm0_cntl        = 'd0         ;
    std__pe56__lane22_strm0_data        = 'h1234_5678 ;
    std__pe56__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe56__lane22_strm1_cntl        = 'd0         ;
    std__pe56__lane22_strm1_data        = 'h1234_5678 ;
    std__pe56__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe56__lane23_strm0_cntl        = 'd0         ;
    std__pe56__lane23_strm0_data        = 'h1234_5678 ;
    std__pe56__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe56__lane23_strm1_cntl        = 'd0         ;
    std__pe56__lane23_strm1_data        = 'h1234_5678 ;
    std__pe56__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe56__lane24_strm0_cntl        = 'd0         ;
    std__pe56__lane24_strm0_data        = 'h1234_5678 ;
    std__pe56__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe56__lane24_strm1_cntl        = 'd0         ;
    std__pe56__lane24_strm1_data        = 'h1234_5678 ;
    std__pe56__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe56__lane25_strm0_cntl        = 'd0         ;
    std__pe56__lane25_strm0_data        = 'h1234_5678 ;
    std__pe56__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe56__lane25_strm1_cntl        = 'd0         ;
    std__pe56__lane25_strm1_data        = 'h1234_5678 ;
    std__pe56__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe56__lane26_strm0_cntl        = 'd0         ;
    std__pe56__lane26_strm0_data        = 'h1234_5678 ;
    std__pe56__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe56__lane26_strm1_cntl        = 'd0         ;
    std__pe56__lane26_strm1_data        = 'h1234_5678 ;
    std__pe56__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe56__lane27_strm0_cntl        = 'd0         ;
    std__pe56__lane27_strm0_data        = 'h1234_5678 ;
    std__pe56__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe56__lane27_strm1_cntl        = 'd0         ;
    std__pe56__lane27_strm1_data        = 'h1234_5678 ;
    std__pe56__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe56__lane28_strm0_cntl        = 'd0         ;
    std__pe56__lane28_strm0_data        = 'h1234_5678 ;
    std__pe56__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe56__lane28_strm1_cntl        = 'd0         ;
    std__pe56__lane28_strm1_data        = 'h1234_5678 ;
    std__pe56__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe56__lane29_strm0_cntl        = 'd0         ;
    std__pe56__lane29_strm0_data        = 'h1234_5678 ;
    std__pe56__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe56__lane29_strm1_cntl        = 'd0         ;
    std__pe56__lane29_strm1_data        = 'h1234_5678 ;
    std__pe56__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe56__lane30_strm0_cntl        = 'd0         ;
    std__pe56__lane30_strm0_data        = 'h1234_5678 ;
    std__pe56__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe56__lane30_strm1_cntl        = 'd0         ;
    std__pe56__lane30_strm1_data        = 'h1234_5678 ;
    std__pe56__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe56__lane31_strm0_cntl        = 'd0         ;
    std__pe56__lane31_strm0_data        = 'h1234_5678 ;
    std__pe56__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe56__lane31_strm1_cntl        = 'd0         ;
    std__pe56__lane31_strm1_data        = 'h1234_5678 ;
    std__pe56__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe57__lane0_strm0_cntl        = 'd0         ;
    std__pe57__lane0_strm0_data        = 'h1234_5678 ;
    std__pe57__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe57__lane0_strm1_cntl        = 'd0         ;
    std__pe57__lane0_strm1_data        = 'h1234_5678 ;
    std__pe57__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe57__lane1_strm0_cntl        = 'd0         ;
    std__pe57__lane1_strm0_data        = 'h1234_5678 ;
    std__pe57__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe57__lane1_strm1_cntl        = 'd0         ;
    std__pe57__lane1_strm1_data        = 'h1234_5678 ;
    std__pe57__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe57__lane2_strm0_cntl        = 'd0         ;
    std__pe57__lane2_strm0_data        = 'h1234_5678 ;
    std__pe57__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe57__lane2_strm1_cntl        = 'd0         ;
    std__pe57__lane2_strm1_data        = 'h1234_5678 ;
    std__pe57__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe57__lane3_strm0_cntl        = 'd0         ;
    std__pe57__lane3_strm0_data        = 'h1234_5678 ;
    std__pe57__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe57__lane3_strm1_cntl        = 'd0         ;
    std__pe57__lane3_strm1_data        = 'h1234_5678 ;
    std__pe57__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe57__lane4_strm0_cntl        = 'd0         ;
    std__pe57__lane4_strm0_data        = 'h1234_5678 ;
    std__pe57__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe57__lane4_strm1_cntl        = 'd0         ;
    std__pe57__lane4_strm1_data        = 'h1234_5678 ;
    std__pe57__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe57__lane5_strm0_cntl        = 'd0         ;
    std__pe57__lane5_strm0_data        = 'h1234_5678 ;
    std__pe57__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe57__lane5_strm1_cntl        = 'd0         ;
    std__pe57__lane5_strm1_data        = 'h1234_5678 ;
    std__pe57__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe57__lane6_strm0_cntl        = 'd0         ;
    std__pe57__lane6_strm0_data        = 'h1234_5678 ;
    std__pe57__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe57__lane6_strm1_cntl        = 'd0         ;
    std__pe57__lane6_strm1_data        = 'h1234_5678 ;
    std__pe57__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe57__lane7_strm0_cntl        = 'd0         ;
    std__pe57__lane7_strm0_data        = 'h1234_5678 ;
    std__pe57__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe57__lane7_strm1_cntl        = 'd0         ;
    std__pe57__lane7_strm1_data        = 'h1234_5678 ;
    std__pe57__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe57__lane8_strm0_cntl        = 'd0         ;
    std__pe57__lane8_strm0_data        = 'h1234_5678 ;
    std__pe57__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe57__lane8_strm1_cntl        = 'd0         ;
    std__pe57__lane8_strm1_data        = 'h1234_5678 ;
    std__pe57__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe57__lane9_strm0_cntl        = 'd0         ;
    std__pe57__lane9_strm0_data        = 'h1234_5678 ;
    std__pe57__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe57__lane9_strm1_cntl        = 'd0         ;
    std__pe57__lane9_strm1_data        = 'h1234_5678 ;
    std__pe57__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe57__lane10_strm0_cntl        = 'd0         ;
    std__pe57__lane10_strm0_data        = 'h1234_5678 ;
    std__pe57__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe57__lane10_strm1_cntl        = 'd0         ;
    std__pe57__lane10_strm1_data        = 'h1234_5678 ;
    std__pe57__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe57__lane11_strm0_cntl        = 'd0         ;
    std__pe57__lane11_strm0_data        = 'h1234_5678 ;
    std__pe57__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe57__lane11_strm1_cntl        = 'd0         ;
    std__pe57__lane11_strm1_data        = 'h1234_5678 ;
    std__pe57__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe57__lane12_strm0_cntl        = 'd0         ;
    std__pe57__lane12_strm0_data        = 'h1234_5678 ;
    std__pe57__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe57__lane12_strm1_cntl        = 'd0         ;
    std__pe57__lane12_strm1_data        = 'h1234_5678 ;
    std__pe57__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe57__lane13_strm0_cntl        = 'd0         ;
    std__pe57__lane13_strm0_data        = 'h1234_5678 ;
    std__pe57__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe57__lane13_strm1_cntl        = 'd0         ;
    std__pe57__lane13_strm1_data        = 'h1234_5678 ;
    std__pe57__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe57__lane14_strm0_cntl        = 'd0         ;
    std__pe57__lane14_strm0_data        = 'h1234_5678 ;
    std__pe57__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe57__lane14_strm1_cntl        = 'd0         ;
    std__pe57__lane14_strm1_data        = 'h1234_5678 ;
    std__pe57__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe57__lane15_strm0_cntl        = 'd0         ;
    std__pe57__lane15_strm0_data        = 'h1234_5678 ;
    std__pe57__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe57__lane15_strm1_cntl        = 'd0         ;
    std__pe57__lane15_strm1_data        = 'h1234_5678 ;
    std__pe57__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe57__lane16_strm0_cntl        = 'd0         ;
    std__pe57__lane16_strm0_data        = 'h1234_5678 ;
    std__pe57__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe57__lane16_strm1_cntl        = 'd0         ;
    std__pe57__lane16_strm1_data        = 'h1234_5678 ;
    std__pe57__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe57__lane17_strm0_cntl        = 'd0         ;
    std__pe57__lane17_strm0_data        = 'h1234_5678 ;
    std__pe57__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe57__lane17_strm1_cntl        = 'd0         ;
    std__pe57__lane17_strm1_data        = 'h1234_5678 ;
    std__pe57__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe57__lane18_strm0_cntl        = 'd0         ;
    std__pe57__lane18_strm0_data        = 'h1234_5678 ;
    std__pe57__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe57__lane18_strm1_cntl        = 'd0         ;
    std__pe57__lane18_strm1_data        = 'h1234_5678 ;
    std__pe57__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe57__lane19_strm0_cntl        = 'd0         ;
    std__pe57__lane19_strm0_data        = 'h1234_5678 ;
    std__pe57__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe57__lane19_strm1_cntl        = 'd0         ;
    std__pe57__lane19_strm1_data        = 'h1234_5678 ;
    std__pe57__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe57__lane20_strm0_cntl        = 'd0         ;
    std__pe57__lane20_strm0_data        = 'h1234_5678 ;
    std__pe57__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe57__lane20_strm1_cntl        = 'd0         ;
    std__pe57__lane20_strm1_data        = 'h1234_5678 ;
    std__pe57__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe57__lane21_strm0_cntl        = 'd0         ;
    std__pe57__lane21_strm0_data        = 'h1234_5678 ;
    std__pe57__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe57__lane21_strm1_cntl        = 'd0         ;
    std__pe57__lane21_strm1_data        = 'h1234_5678 ;
    std__pe57__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe57__lane22_strm0_cntl        = 'd0         ;
    std__pe57__lane22_strm0_data        = 'h1234_5678 ;
    std__pe57__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe57__lane22_strm1_cntl        = 'd0         ;
    std__pe57__lane22_strm1_data        = 'h1234_5678 ;
    std__pe57__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe57__lane23_strm0_cntl        = 'd0         ;
    std__pe57__lane23_strm0_data        = 'h1234_5678 ;
    std__pe57__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe57__lane23_strm1_cntl        = 'd0         ;
    std__pe57__lane23_strm1_data        = 'h1234_5678 ;
    std__pe57__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe57__lane24_strm0_cntl        = 'd0         ;
    std__pe57__lane24_strm0_data        = 'h1234_5678 ;
    std__pe57__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe57__lane24_strm1_cntl        = 'd0         ;
    std__pe57__lane24_strm1_data        = 'h1234_5678 ;
    std__pe57__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe57__lane25_strm0_cntl        = 'd0         ;
    std__pe57__lane25_strm0_data        = 'h1234_5678 ;
    std__pe57__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe57__lane25_strm1_cntl        = 'd0         ;
    std__pe57__lane25_strm1_data        = 'h1234_5678 ;
    std__pe57__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe57__lane26_strm0_cntl        = 'd0         ;
    std__pe57__lane26_strm0_data        = 'h1234_5678 ;
    std__pe57__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe57__lane26_strm1_cntl        = 'd0         ;
    std__pe57__lane26_strm1_data        = 'h1234_5678 ;
    std__pe57__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe57__lane27_strm0_cntl        = 'd0         ;
    std__pe57__lane27_strm0_data        = 'h1234_5678 ;
    std__pe57__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe57__lane27_strm1_cntl        = 'd0         ;
    std__pe57__lane27_strm1_data        = 'h1234_5678 ;
    std__pe57__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe57__lane28_strm0_cntl        = 'd0         ;
    std__pe57__lane28_strm0_data        = 'h1234_5678 ;
    std__pe57__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe57__lane28_strm1_cntl        = 'd0         ;
    std__pe57__lane28_strm1_data        = 'h1234_5678 ;
    std__pe57__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe57__lane29_strm0_cntl        = 'd0         ;
    std__pe57__lane29_strm0_data        = 'h1234_5678 ;
    std__pe57__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe57__lane29_strm1_cntl        = 'd0         ;
    std__pe57__lane29_strm1_data        = 'h1234_5678 ;
    std__pe57__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe57__lane30_strm0_cntl        = 'd0         ;
    std__pe57__lane30_strm0_data        = 'h1234_5678 ;
    std__pe57__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe57__lane30_strm1_cntl        = 'd0         ;
    std__pe57__lane30_strm1_data        = 'h1234_5678 ;
    std__pe57__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe57__lane31_strm0_cntl        = 'd0         ;
    std__pe57__lane31_strm0_data        = 'h1234_5678 ;
    std__pe57__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe57__lane31_strm1_cntl        = 'd0         ;
    std__pe57__lane31_strm1_data        = 'h1234_5678 ;
    std__pe57__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe58__lane0_strm0_cntl        = 'd0         ;
    std__pe58__lane0_strm0_data        = 'h1234_5678 ;
    std__pe58__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe58__lane0_strm1_cntl        = 'd0         ;
    std__pe58__lane0_strm1_data        = 'h1234_5678 ;
    std__pe58__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe58__lane1_strm0_cntl        = 'd0         ;
    std__pe58__lane1_strm0_data        = 'h1234_5678 ;
    std__pe58__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe58__lane1_strm1_cntl        = 'd0         ;
    std__pe58__lane1_strm1_data        = 'h1234_5678 ;
    std__pe58__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe58__lane2_strm0_cntl        = 'd0         ;
    std__pe58__lane2_strm0_data        = 'h1234_5678 ;
    std__pe58__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe58__lane2_strm1_cntl        = 'd0         ;
    std__pe58__lane2_strm1_data        = 'h1234_5678 ;
    std__pe58__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe58__lane3_strm0_cntl        = 'd0         ;
    std__pe58__lane3_strm0_data        = 'h1234_5678 ;
    std__pe58__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe58__lane3_strm1_cntl        = 'd0         ;
    std__pe58__lane3_strm1_data        = 'h1234_5678 ;
    std__pe58__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe58__lane4_strm0_cntl        = 'd0         ;
    std__pe58__lane4_strm0_data        = 'h1234_5678 ;
    std__pe58__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe58__lane4_strm1_cntl        = 'd0         ;
    std__pe58__lane4_strm1_data        = 'h1234_5678 ;
    std__pe58__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe58__lane5_strm0_cntl        = 'd0         ;
    std__pe58__lane5_strm0_data        = 'h1234_5678 ;
    std__pe58__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe58__lane5_strm1_cntl        = 'd0         ;
    std__pe58__lane5_strm1_data        = 'h1234_5678 ;
    std__pe58__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe58__lane6_strm0_cntl        = 'd0         ;
    std__pe58__lane6_strm0_data        = 'h1234_5678 ;
    std__pe58__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe58__lane6_strm1_cntl        = 'd0         ;
    std__pe58__lane6_strm1_data        = 'h1234_5678 ;
    std__pe58__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe58__lane7_strm0_cntl        = 'd0         ;
    std__pe58__lane7_strm0_data        = 'h1234_5678 ;
    std__pe58__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe58__lane7_strm1_cntl        = 'd0         ;
    std__pe58__lane7_strm1_data        = 'h1234_5678 ;
    std__pe58__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe58__lane8_strm0_cntl        = 'd0         ;
    std__pe58__lane8_strm0_data        = 'h1234_5678 ;
    std__pe58__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe58__lane8_strm1_cntl        = 'd0         ;
    std__pe58__lane8_strm1_data        = 'h1234_5678 ;
    std__pe58__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe58__lane9_strm0_cntl        = 'd0         ;
    std__pe58__lane9_strm0_data        = 'h1234_5678 ;
    std__pe58__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe58__lane9_strm1_cntl        = 'd0         ;
    std__pe58__lane9_strm1_data        = 'h1234_5678 ;
    std__pe58__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe58__lane10_strm0_cntl        = 'd0         ;
    std__pe58__lane10_strm0_data        = 'h1234_5678 ;
    std__pe58__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe58__lane10_strm1_cntl        = 'd0         ;
    std__pe58__lane10_strm1_data        = 'h1234_5678 ;
    std__pe58__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe58__lane11_strm0_cntl        = 'd0         ;
    std__pe58__lane11_strm0_data        = 'h1234_5678 ;
    std__pe58__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe58__lane11_strm1_cntl        = 'd0         ;
    std__pe58__lane11_strm1_data        = 'h1234_5678 ;
    std__pe58__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe58__lane12_strm0_cntl        = 'd0         ;
    std__pe58__lane12_strm0_data        = 'h1234_5678 ;
    std__pe58__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe58__lane12_strm1_cntl        = 'd0         ;
    std__pe58__lane12_strm1_data        = 'h1234_5678 ;
    std__pe58__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe58__lane13_strm0_cntl        = 'd0         ;
    std__pe58__lane13_strm0_data        = 'h1234_5678 ;
    std__pe58__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe58__lane13_strm1_cntl        = 'd0         ;
    std__pe58__lane13_strm1_data        = 'h1234_5678 ;
    std__pe58__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe58__lane14_strm0_cntl        = 'd0         ;
    std__pe58__lane14_strm0_data        = 'h1234_5678 ;
    std__pe58__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe58__lane14_strm1_cntl        = 'd0         ;
    std__pe58__lane14_strm1_data        = 'h1234_5678 ;
    std__pe58__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe58__lane15_strm0_cntl        = 'd0         ;
    std__pe58__lane15_strm0_data        = 'h1234_5678 ;
    std__pe58__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe58__lane15_strm1_cntl        = 'd0         ;
    std__pe58__lane15_strm1_data        = 'h1234_5678 ;
    std__pe58__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe58__lane16_strm0_cntl        = 'd0         ;
    std__pe58__lane16_strm0_data        = 'h1234_5678 ;
    std__pe58__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe58__lane16_strm1_cntl        = 'd0         ;
    std__pe58__lane16_strm1_data        = 'h1234_5678 ;
    std__pe58__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe58__lane17_strm0_cntl        = 'd0         ;
    std__pe58__lane17_strm0_data        = 'h1234_5678 ;
    std__pe58__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe58__lane17_strm1_cntl        = 'd0         ;
    std__pe58__lane17_strm1_data        = 'h1234_5678 ;
    std__pe58__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe58__lane18_strm0_cntl        = 'd0         ;
    std__pe58__lane18_strm0_data        = 'h1234_5678 ;
    std__pe58__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe58__lane18_strm1_cntl        = 'd0         ;
    std__pe58__lane18_strm1_data        = 'h1234_5678 ;
    std__pe58__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe58__lane19_strm0_cntl        = 'd0         ;
    std__pe58__lane19_strm0_data        = 'h1234_5678 ;
    std__pe58__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe58__lane19_strm1_cntl        = 'd0         ;
    std__pe58__lane19_strm1_data        = 'h1234_5678 ;
    std__pe58__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe58__lane20_strm0_cntl        = 'd0         ;
    std__pe58__lane20_strm0_data        = 'h1234_5678 ;
    std__pe58__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe58__lane20_strm1_cntl        = 'd0         ;
    std__pe58__lane20_strm1_data        = 'h1234_5678 ;
    std__pe58__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe58__lane21_strm0_cntl        = 'd0         ;
    std__pe58__lane21_strm0_data        = 'h1234_5678 ;
    std__pe58__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe58__lane21_strm1_cntl        = 'd0         ;
    std__pe58__lane21_strm1_data        = 'h1234_5678 ;
    std__pe58__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe58__lane22_strm0_cntl        = 'd0         ;
    std__pe58__lane22_strm0_data        = 'h1234_5678 ;
    std__pe58__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe58__lane22_strm1_cntl        = 'd0         ;
    std__pe58__lane22_strm1_data        = 'h1234_5678 ;
    std__pe58__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe58__lane23_strm0_cntl        = 'd0         ;
    std__pe58__lane23_strm0_data        = 'h1234_5678 ;
    std__pe58__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe58__lane23_strm1_cntl        = 'd0         ;
    std__pe58__lane23_strm1_data        = 'h1234_5678 ;
    std__pe58__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe58__lane24_strm0_cntl        = 'd0         ;
    std__pe58__lane24_strm0_data        = 'h1234_5678 ;
    std__pe58__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe58__lane24_strm1_cntl        = 'd0         ;
    std__pe58__lane24_strm1_data        = 'h1234_5678 ;
    std__pe58__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe58__lane25_strm0_cntl        = 'd0         ;
    std__pe58__lane25_strm0_data        = 'h1234_5678 ;
    std__pe58__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe58__lane25_strm1_cntl        = 'd0         ;
    std__pe58__lane25_strm1_data        = 'h1234_5678 ;
    std__pe58__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe58__lane26_strm0_cntl        = 'd0         ;
    std__pe58__lane26_strm0_data        = 'h1234_5678 ;
    std__pe58__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe58__lane26_strm1_cntl        = 'd0         ;
    std__pe58__lane26_strm1_data        = 'h1234_5678 ;
    std__pe58__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe58__lane27_strm0_cntl        = 'd0         ;
    std__pe58__lane27_strm0_data        = 'h1234_5678 ;
    std__pe58__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe58__lane27_strm1_cntl        = 'd0         ;
    std__pe58__lane27_strm1_data        = 'h1234_5678 ;
    std__pe58__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe58__lane28_strm0_cntl        = 'd0         ;
    std__pe58__lane28_strm0_data        = 'h1234_5678 ;
    std__pe58__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe58__lane28_strm1_cntl        = 'd0         ;
    std__pe58__lane28_strm1_data        = 'h1234_5678 ;
    std__pe58__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe58__lane29_strm0_cntl        = 'd0         ;
    std__pe58__lane29_strm0_data        = 'h1234_5678 ;
    std__pe58__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe58__lane29_strm1_cntl        = 'd0         ;
    std__pe58__lane29_strm1_data        = 'h1234_5678 ;
    std__pe58__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe58__lane30_strm0_cntl        = 'd0         ;
    std__pe58__lane30_strm0_data        = 'h1234_5678 ;
    std__pe58__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe58__lane30_strm1_cntl        = 'd0         ;
    std__pe58__lane30_strm1_data        = 'h1234_5678 ;
    std__pe58__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe58__lane31_strm0_cntl        = 'd0         ;
    std__pe58__lane31_strm0_data        = 'h1234_5678 ;
    std__pe58__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe58__lane31_strm1_cntl        = 'd0         ;
    std__pe58__lane31_strm1_data        = 'h1234_5678 ;
    std__pe58__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe59__lane0_strm0_cntl        = 'd0         ;
    std__pe59__lane0_strm0_data        = 'h1234_5678 ;
    std__pe59__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe59__lane0_strm1_cntl        = 'd0         ;
    std__pe59__lane0_strm1_data        = 'h1234_5678 ;
    std__pe59__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe59__lane1_strm0_cntl        = 'd0         ;
    std__pe59__lane1_strm0_data        = 'h1234_5678 ;
    std__pe59__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe59__lane1_strm1_cntl        = 'd0         ;
    std__pe59__lane1_strm1_data        = 'h1234_5678 ;
    std__pe59__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe59__lane2_strm0_cntl        = 'd0         ;
    std__pe59__lane2_strm0_data        = 'h1234_5678 ;
    std__pe59__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe59__lane2_strm1_cntl        = 'd0         ;
    std__pe59__lane2_strm1_data        = 'h1234_5678 ;
    std__pe59__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe59__lane3_strm0_cntl        = 'd0         ;
    std__pe59__lane3_strm0_data        = 'h1234_5678 ;
    std__pe59__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe59__lane3_strm1_cntl        = 'd0         ;
    std__pe59__lane3_strm1_data        = 'h1234_5678 ;
    std__pe59__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe59__lane4_strm0_cntl        = 'd0         ;
    std__pe59__lane4_strm0_data        = 'h1234_5678 ;
    std__pe59__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe59__lane4_strm1_cntl        = 'd0         ;
    std__pe59__lane4_strm1_data        = 'h1234_5678 ;
    std__pe59__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe59__lane5_strm0_cntl        = 'd0         ;
    std__pe59__lane5_strm0_data        = 'h1234_5678 ;
    std__pe59__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe59__lane5_strm1_cntl        = 'd0         ;
    std__pe59__lane5_strm1_data        = 'h1234_5678 ;
    std__pe59__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe59__lane6_strm0_cntl        = 'd0         ;
    std__pe59__lane6_strm0_data        = 'h1234_5678 ;
    std__pe59__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe59__lane6_strm1_cntl        = 'd0         ;
    std__pe59__lane6_strm1_data        = 'h1234_5678 ;
    std__pe59__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe59__lane7_strm0_cntl        = 'd0         ;
    std__pe59__lane7_strm0_data        = 'h1234_5678 ;
    std__pe59__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe59__lane7_strm1_cntl        = 'd0         ;
    std__pe59__lane7_strm1_data        = 'h1234_5678 ;
    std__pe59__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe59__lane8_strm0_cntl        = 'd0         ;
    std__pe59__lane8_strm0_data        = 'h1234_5678 ;
    std__pe59__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe59__lane8_strm1_cntl        = 'd0         ;
    std__pe59__lane8_strm1_data        = 'h1234_5678 ;
    std__pe59__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe59__lane9_strm0_cntl        = 'd0         ;
    std__pe59__lane9_strm0_data        = 'h1234_5678 ;
    std__pe59__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe59__lane9_strm1_cntl        = 'd0         ;
    std__pe59__lane9_strm1_data        = 'h1234_5678 ;
    std__pe59__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe59__lane10_strm0_cntl        = 'd0         ;
    std__pe59__lane10_strm0_data        = 'h1234_5678 ;
    std__pe59__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe59__lane10_strm1_cntl        = 'd0         ;
    std__pe59__lane10_strm1_data        = 'h1234_5678 ;
    std__pe59__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe59__lane11_strm0_cntl        = 'd0         ;
    std__pe59__lane11_strm0_data        = 'h1234_5678 ;
    std__pe59__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe59__lane11_strm1_cntl        = 'd0         ;
    std__pe59__lane11_strm1_data        = 'h1234_5678 ;
    std__pe59__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe59__lane12_strm0_cntl        = 'd0         ;
    std__pe59__lane12_strm0_data        = 'h1234_5678 ;
    std__pe59__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe59__lane12_strm1_cntl        = 'd0         ;
    std__pe59__lane12_strm1_data        = 'h1234_5678 ;
    std__pe59__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe59__lane13_strm0_cntl        = 'd0         ;
    std__pe59__lane13_strm0_data        = 'h1234_5678 ;
    std__pe59__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe59__lane13_strm1_cntl        = 'd0         ;
    std__pe59__lane13_strm1_data        = 'h1234_5678 ;
    std__pe59__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe59__lane14_strm0_cntl        = 'd0         ;
    std__pe59__lane14_strm0_data        = 'h1234_5678 ;
    std__pe59__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe59__lane14_strm1_cntl        = 'd0         ;
    std__pe59__lane14_strm1_data        = 'h1234_5678 ;
    std__pe59__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe59__lane15_strm0_cntl        = 'd0         ;
    std__pe59__lane15_strm0_data        = 'h1234_5678 ;
    std__pe59__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe59__lane15_strm1_cntl        = 'd0         ;
    std__pe59__lane15_strm1_data        = 'h1234_5678 ;
    std__pe59__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe59__lane16_strm0_cntl        = 'd0         ;
    std__pe59__lane16_strm0_data        = 'h1234_5678 ;
    std__pe59__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe59__lane16_strm1_cntl        = 'd0         ;
    std__pe59__lane16_strm1_data        = 'h1234_5678 ;
    std__pe59__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe59__lane17_strm0_cntl        = 'd0         ;
    std__pe59__lane17_strm0_data        = 'h1234_5678 ;
    std__pe59__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe59__lane17_strm1_cntl        = 'd0         ;
    std__pe59__lane17_strm1_data        = 'h1234_5678 ;
    std__pe59__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe59__lane18_strm0_cntl        = 'd0         ;
    std__pe59__lane18_strm0_data        = 'h1234_5678 ;
    std__pe59__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe59__lane18_strm1_cntl        = 'd0         ;
    std__pe59__lane18_strm1_data        = 'h1234_5678 ;
    std__pe59__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe59__lane19_strm0_cntl        = 'd0         ;
    std__pe59__lane19_strm0_data        = 'h1234_5678 ;
    std__pe59__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe59__lane19_strm1_cntl        = 'd0         ;
    std__pe59__lane19_strm1_data        = 'h1234_5678 ;
    std__pe59__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe59__lane20_strm0_cntl        = 'd0         ;
    std__pe59__lane20_strm0_data        = 'h1234_5678 ;
    std__pe59__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe59__lane20_strm1_cntl        = 'd0         ;
    std__pe59__lane20_strm1_data        = 'h1234_5678 ;
    std__pe59__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe59__lane21_strm0_cntl        = 'd0         ;
    std__pe59__lane21_strm0_data        = 'h1234_5678 ;
    std__pe59__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe59__lane21_strm1_cntl        = 'd0         ;
    std__pe59__lane21_strm1_data        = 'h1234_5678 ;
    std__pe59__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe59__lane22_strm0_cntl        = 'd0         ;
    std__pe59__lane22_strm0_data        = 'h1234_5678 ;
    std__pe59__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe59__lane22_strm1_cntl        = 'd0         ;
    std__pe59__lane22_strm1_data        = 'h1234_5678 ;
    std__pe59__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe59__lane23_strm0_cntl        = 'd0         ;
    std__pe59__lane23_strm0_data        = 'h1234_5678 ;
    std__pe59__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe59__lane23_strm1_cntl        = 'd0         ;
    std__pe59__lane23_strm1_data        = 'h1234_5678 ;
    std__pe59__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe59__lane24_strm0_cntl        = 'd0         ;
    std__pe59__lane24_strm0_data        = 'h1234_5678 ;
    std__pe59__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe59__lane24_strm1_cntl        = 'd0         ;
    std__pe59__lane24_strm1_data        = 'h1234_5678 ;
    std__pe59__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe59__lane25_strm0_cntl        = 'd0         ;
    std__pe59__lane25_strm0_data        = 'h1234_5678 ;
    std__pe59__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe59__lane25_strm1_cntl        = 'd0         ;
    std__pe59__lane25_strm1_data        = 'h1234_5678 ;
    std__pe59__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe59__lane26_strm0_cntl        = 'd0         ;
    std__pe59__lane26_strm0_data        = 'h1234_5678 ;
    std__pe59__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe59__lane26_strm1_cntl        = 'd0         ;
    std__pe59__lane26_strm1_data        = 'h1234_5678 ;
    std__pe59__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe59__lane27_strm0_cntl        = 'd0         ;
    std__pe59__lane27_strm0_data        = 'h1234_5678 ;
    std__pe59__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe59__lane27_strm1_cntl        = 'd0         ;
    std__pe59__lane27_strm1_data        = 'h1234_5678 ;
    std__pe59__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe59__lane28_strm0_cntl        = 'd0         ;
    std__pe59__lane28_strm0_data        = 'h1234_5678 ;
    std__pe59__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe59__lane28_strm1_cntl        = 'd0         ;
    std__pe59__lane28_strm1_data        = 'h1234_5678 ;
    std__pe59__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe59__lane29_strm0_cntl        = 'd0         ;
    std__pe59__lane29_strm0_data        = 'h1234_5678 ;
    std__pe59__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe59__lane29_strm1_cntl        = 'd0         ;
    std__pe59__lane29_strm1_data        = 'h1234_5678 ;
    std__pe59__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe59__lane30_strm0_cntl        = 'd0         ;
    std__pe59__lane30_strm0_data        = 'h1234_5678 ;
    std__pe59__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe59__lane30_strm1_cntl        = 'd0         ;
    std__pe59__lane30_strm1_data        = 'h1234_5678 ;
    std__pe59__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe59__lane31_strm0_cntl        = 'd0         ;
    std__pe59__lane31_strm0_data        = 'h1234_5678 ;
    std__pe59__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe59__lane31_strm1_cntl        = 'd0         ;
    std__pe59__lane31_strm1_data        = 'h1234_5678 ;
    std__pe59__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe60__lane0_strm0_cntl        = 'd0         ;
    std__pe60__lane0_strm0_data        = 'h1234_5678 ;
    std__pe60__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe60__lane0_strm1_cntl        = 'd0         ;
    std__pe60__lane0_strm1_data        = 'h1234_5678 ;
    std__pe60__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe60__lane1_strm0_cntl        = 'd0         ;
    std__pe60__lane1_strm0_data        = 'h1234_5678 ;
    std__pe60__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe60__lane1_strm1_cntl        = 'd0         ;
    std__pe60__lane1_strm1_data        = 'h1234_5678 ;
    std__pe60__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe60__lane2_strm0_cntl        = 'd0         ;
    std__pe60__lane2_strm0_data        = 'h1234_5678 ;
    std__pe60__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe60__lane2_strm1_cntl        = 'd0         ;
    std__pe60__lane2_strm1_data        = 'h1234_5678 ;
    std__pe60__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe60__lane3_strm0_cntl        = 'd0         ;
    std__pe60__lane3_strm0_data        = 'h1234_5678 ;
    std__pe60__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe60__lane3_strm1_cntl        = 'd0         ;
    std__pe60__lane3_strm1_data        = 'h1234_5678 ;
    std__pe60__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe60__lane4_strm0_cntl        = 'd0         ;
    std__pe60__lane4_strm0_data        = 'h1234_5678 ;
    std__pe60__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe60__lane4_strm1_cntl        = 'd0         ;
    std__pe60__lane4_strm1_data        = 'h1234_5678 ;
    std__pe60__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe60__lane5_strm0_cntl        = 'd0         ;
    std__pe60__lane5_strm0_data        = 'h1234_5678 ;
    std__pe60__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe60__lane5_strm1_cntl        = 'd0         ;
    std__pe60__lane5_strm1_data        = 'h1234_5678 ;
    std__pe60__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe60__lane6_strm0_cntl        = 'd0         ;
    std__pe60__lane6_strm0_data        = 'h1234_5678 ;
    std__pe60__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe60__lane6_strm1_cntl        = 'd0         ;
    std__pe60__lane6_strm1_data        = 'h1234_5678 ;
    std__pe60__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe60__lane7_strm0_cntl        = 'd0         ;
    std__pe60__lane7_strm0_data        = 'h1234_5678 ;
    std__pe60__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe60__lane7_strm1_cntl        = 'd0         ;
    std__pe60__lane7_strm1_data        = 'h1234_5678 ;
    std__pe60__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe60__lane8_strm0_cntl        = 'd0         ;
    std__pe60__lane8_strm0_data        = 'h1234_5678 ;
    std__pe60__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe60__lane8_strm1_cntl        = 'd0         ;
    std__pe60__lane8_strm1_data        = 'h1234_5678 ;
    std__pe60__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe60__lane9_strm0_cntl        = 'd0         ;
    std__pe60__lane9_strm0_data        = 'h1234_5678 ;
    std__pe60__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe60__lane9_strm1_cntl        = 'd0         ;
    std__pe60__lane9_strm1_data        = 'h1234_5678 ;
    std__pe60__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe60__lane10_strm0_cntl        = 'd0         ;
    std__pe60__lane10_strm0_data        = 'h1234_5678 ;
    std__pe60__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe60__lane10_strm1_cntl        = 'd0         ;
    std__pe60__lane10_strm1_data        = 'h1234_5678 ;
    std__pe60__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe60__lane11_strm0_cntl        = 'd0         ;
    std__pe60__lane11_strm0_data        = 'h1234_5678 ;
    std__pe60__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe60__lane11_strm1_cntl        = 'd0         ;
    std__pe60__lane11_strm1_data        = 'h1234_5678 ;
    std__pe60__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe60__lane12_strm0_cntl        = 'd0         ;
    std__pe60__lane12_strm0_data        = 'h1234_5678 ;
    std__pe60__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe60__lane12_strm1_cntl        = 'd0         ;
    std__pe60__lane12_strm1_data        = 'h1234_5678 ;
    std__pe60__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe60__lane13_strm0_cntl        = 'd0         ;
    std__pe60__lane13_strm0_data        = 'h1234_5678 ;
    std__pe60__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe60__lane13_strm1_cntl        = 'd0         ;
    std__pe60__lane13_strm1_data        = 'h1234_5678 ;
    std__pe60__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe60__lane14_strm0_cntl        = 'd0         ;
    std__pe60__lane14_strm0_data        = 'h1234_5678 ;
    std__pe60__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe60__lane14_strm1_cntl        = 'd0         ;
    std__pe60__lane14_strm1_data        = 'h1234_5678 ;
    std__pe60__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe60__lane15_strm0_cntl        = 'd0         ;
    std__pe60__lane15_strm0_data        = 'h1234_5678 ;
    std__pe60__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe60__lane15_strm1_cntl        = 'd0         ;
    std__pe60__lane15_strm1_data        = 'h1234_5678 ;
    std__pe60__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe60__lane16_strm0_cntl        = 'd0         ;
    std__pe60__lane16_strm0_data        = 'h1234_5678 ;
    std__pe60__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe60__lane16_strm1_cntl        = 'd0         ;
    std__pe60__lane16_strm1_data        = 'h1234_5678 ;
    std__pe60__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe60__lane17_strm0_cntl        = 'd0         ;
    std__pe60__lane17_strm0_data        = 'h1234_5678 ;
    std__pe60__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe60__lane17_strm1_cntl        = 'd0         ;
    std__pe60__lane17_strm1_data        = 'h1234_5678 ;
    std__pe60__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe60__lane18_strm0_cntl        = 'd0         ;
    std__pe60__lane18_strm0_data        = 'h1234_5678 ;
    std__pe60__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe60__lane18_strm1_cntl        = 'd0         ;
    std__pe60__lane18_strm1_data        = 'h1234_5678 ;
    std__pe60__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe60__lane19_strm0_cntl        = 'd0         ;
    std__pe60__lane19_strm0_data        = 'h1234_5678 ;
    std__pe60__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe60__lane19_strm1_cntl        = 'd0         ;
    std__pe60__lane19_strm1_data        = 'h1234_5678 ;
    std__pe60__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe60__lane20_strm0_cntl        = 'd0         ;
    std__pe60__lane20_strm0_data        = 'h1234_5678 ;
    std__pe60__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe60__lane20_strm1_cntl        = 'd0         ;
    std__pe60__lane20_strm1_data        = 'h1234_5678 ;
    std__pe60__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe60__lane21_strm0_cntl        = 'd0         ;
    std__pe60__lane21_strm0_data        = 'h1234_5678 ;
    std__pe60__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe60__lane21_strm1_cntl        = 'd0         ;
    std__pe60__lane21_strm1_data        = 'h1234_5678 ;
    std__pe60__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe60__lane22_strm0_cntl        = 'd0         ;
    std__pe60__lane22_strm0_data        = 'h1234_5678 ;
    std__pe60__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe60__lane22_strm1_cntl        = 'd0         ;
    std__pe60__lane22_strm1_data        = 'h1234_5678 ;
    std__pe60__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe60__lane23_strm0_cntl        = 'd0         ;
    std__pe60__lane23_strm0_data        = 'h1234_5678 ;
    std__pe60__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe60__lane23_strm1_cntl        = 'd0         ;
    std__pe60__lane23_strm1_data        = 'h1234_5678 ;
    std__pe60__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe60__lane24_strm0_cntl        = 'd0         ;
    std__pe60__lane24_strm0_data        = 'h1234_5678 ;
    std__pe60__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe60__lane24_strm1_cntl        = 'd0         ;
    std__pe60__lane24_strm1_data        = 'h1234_5678 ;
    std__pe60__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe60__lane25_strm0_cntl        = 'd0         ;
    std__pe60__lane25_strm0_data        = 'h1234_5678 ;
    std__pe60__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe60__lane25_strm1_cntl        = 'd0         ;
    std__pe60__lane25_strm1_data        = 'h1234_5678 ;
    std__pe60__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe60__lane26_strm0_cntl        = 'd0         ;
    std__pe60__lane26_strm0_data        = 'h1234_5678 ;
    std__pe60__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe60__lane26_strm1_cntl        = 'd0         ;
    std__pe60__lane26_strm1_data        = 'h1234_5678 ;
    std__pe60__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe60__lane27_strm0_cntl        = 'd0         ;
    std__pe60__lane27_strm0_data        = 'h1234_5678 ;
    std__pe60__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe60__lane27_strm1_cntl        = 'd0         ;
    std__pe60__lane27_strm1_data        = 'h1234_5678 ;
    std__pe60__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe60__lane28_strm0_cntl        = 'd0         ;
    std__pe60__lane28_strm0_data        = 'h1234_5678 ;
    std__pe60__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe60__lane28_strm1_cntl        = 'd0         ;
    std__pe60__lane28_strm1_data        = 'h1234_5678 ;
    std__pe60__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe60__lane29_strm0_cntl        = 'd0         ;
    std__pe60__lane29_strm0_data        = 'h1234_5678 ;
    std__pe60__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe60__lane29_strm1_cntl        = 'd0         ;
    std__pe60__lane29_strm1_data        = 'h1234_5678 ;
    std__pe60__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe60__lane30_strm0_cntl        = 'd0         ;
    std__pe60__lane30_strm0_data        = 'h1234_5678 ;
    std__pe60__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe60__lane30_strm1_cntl        = 'd0         ;
    std__pe60__lane30_strm1_data        = 'h1234_5678 ;
    std__pe60__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe60__lane31_strm0_cntl        = 'd0         ;
    std__pe60__lane31_strm0_data        = 'h1234_5678 ;
    std__pe60__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe60__lane31_strm1_cntl        = 'd0         ;
    std__pe60__lane31_strm1_data        = 'h1234_5678 ;
    std__pe60__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe61__lane0_strm0_cntl        = 'd0         ;
    std__pe61__lane0_strm0_data        = 'h1234_5678 ;
    std__pe61__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe61__lane0_strm1_cntl        = 'd0         ;
    std__pe61__lane0_strm1_data        = 'h1234_5678 ;
    std__pe61__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe61__lane1_strm0_cntl        = 'd0         ;
    std__pe61__lane1_strm0_data        = 'h1234_5678 ;
    std__pe61__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe61__lane1_strm1_cntl        = 'd0         ;
    std__pe61__lane1_strm1_data        = 'h1234_5678 ;
    std__pe61__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe61__lane2_strm0_cntl        = 'd0         ;
    std__pe61__lane2_strm0_data        = 'h1234_5678 ;
    std__pe61__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe61__lane2_strm1_cntl        = 'd0         ;
    std__pe61__lane2_strm1_data        = 'h1234_5678 ;
    std__pe61__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe61__lane3_strm0_cntl        = 'd0         ;
    std__pe61__lane3_strm0_data        = 'h1234_5678 ;
    std__pe61__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe61__lane3_strm1_cntl        = 'd0         ;
    std__pe61__lane3_strm1_data        = 'h1234_5678 ;
    std__pe61__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe61__lane4_strm0_cntl        = 'd0         ;
    std__pe61__lane4_strm0_data        = 'h1234_5678 ;
    std__pe61__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe61__lane4_strm1_cntl        = 'd0         ;
    std__pe61__lane4_strm1_data        = 'h1234_5678 ;
    std__pe61__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe61__lane5_strm0_cntl        = 'd0         ;
    std__pe61__lane5_strm0_data        = 'h1234_5678 ;
    std__pe61__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe61__lane5_strm1_cntl        = 'd0         ;
    std__pe61__lane5_strm1_data        = 'h1234_5678 ;
    std__pe61__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe61__lane6_strm0_cntl        = 'd0         ;
    std__pe61__lane6_strm0_data        = 'h1234_5678 ;
    std__pe61__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe61__lane6_strm1_cntl        = 'd0         ;
    std__pe61__lane6_strm1_data        = 'h1234_5678 ;
    std__pe61__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe61__lane7_strm0_cntl        = 'd0         ;
    std__pe61__lane7_strm0_data        = 'h1234_5678 ;
    std__pe61__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe61__lane7_strm1_cntl        = 'd0         ;
    std__pe61__lane7_strm1_data        = 'h1234_5678 ;
    std__pe61__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe61__lane8_strm0_cntl        = 'd0         ;
    std__pe61__lane8_strm0_data        = 'h1234_5678 ;
    std__pe61__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe61__lane8_strm1_cntl        = 'd0         ;
    std__pe61__lane8_strm1_data        = 'h1234_5678 ;
    std__pe61__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe61__lane9_strm0_cntl        = 'd0         ;
    std__pe61__lane9_strm0_data        = 'h1234_5678 ;
    std__pe61__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe61__lane9_strm1_cntl        = 'd0         ;
    std__pe61__lane9_strm1_data        = 'h1234_5678 ;
    std__pe61__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe61__lane10_strm0_cntl        = 'd0         ;
    std__pe61__lane10_strm0_data        = 'h1234_5678 ;
    std__pe61__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe61__lane10_strm1_cntl        = 'd0         ;
    std__pe61__lane10_strm1_data        = 'h1234_5678 ;
    std__pe61__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe61__lane11_strm0_cntl        = 'd0         ;
    std__pe61__lane11_strm0_data        = 'h1234_5678 ;
    std__pe61__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe61__lane11_strm1_cntl        = 'd0         ;
    std__pe61__lane11_strm1_data        = 'h1234_5678 ;
    std__pe61__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe61__lane12_strm0_cntl        = 'd0         ;
    std__pe61__lane12_strm0_data        = 'h1234_5678 ;
    std__pe61__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe61__lane12_strm1_cntl        = 'd0         ;
    std__pe61__lane12_strm1_data        = 'h1234_5678 ;
    std__pe61__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe61__lane13_strm0_cntl        = 'd0         ;
    std__pe61__lane13_strm0_data        = 'h1234_5678 ;
    std__pe61__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe61__lane13_strm1_cntl        = 'd0         ;
    std__pe61__lane13_strm1_data        = 'h1234_5678 ;
    std__pe61__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe61__lane14_strm0_cntl        = 'd0         ;
    std__pe61__lane14_strm0_data        = 'h1234_5678 ;
    std__pe61__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe61__lane14_strm1_cntl        = 'd0         ;
    std__pe61__lane14_strm1_data        = 'h1234_5678 ;
    std__pe61__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe61__lane15_strm0_cntl        = 'd0         ;
    std__pe61__lane15_strm0_data        = 'h1234_5678 ;
    std__pe61__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe61__lane15_strm1_cntl        = 'd0         ;
    std__pe61__lane15_strm1_data        = 'h1234_5678 ;
    std__pe61__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe61__lane16_strm0_cntl        = 'd0         ;
    std__pe61__lane16_strm0_data        = 'h1234_5678 ;
    std__pe61__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe61__lane16_strm1_cntl        = 'd0         ;
    std__pe61__lane16_strm1_data        = 'h1234_5678 ;
    std__pe61__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe61__lane17_strm0_cntl        = 'd0         ;
    std__pe61__lane17_strm0_data        = 'h1234_5678 ;
    std__pe61__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe61__lane17_strm1_cntl        = 'd0         ;
    std__pe61__lane17_strm1_data        = 'h1234_5678 ;
    std__pe61__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe61__lane18_strm0_cntl        = 'd0         ;
    std__pe61__lane18_strm0_data        = 'h1234_5678 ;
    std__pe61__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe61__lane18_strm1_cntl        = 'd0         ;
    std__pe61__lane18_strm1_data        = 'h1234_5678 ;
    std__pe61__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe61__lane19_strm0_cntl        = 'd0         ;
    std__pe61__lane19_strm0_data        = 'h1234_5678 ;
    std__pe61__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe61__lane19_strm1_cntl        = 'd0         ;
    std__pe61__lane19_strm1_data        = 'h1234_5678 ;
    std__pe61__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe61__lane20_strm0_cntl        = 'd0         ;
    std__pe61__lane20_strm0_data        = 'h1234_5678 ;
    std__pe61__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe61__lane20_strm1_cntl        = 'd0         ;
    std__pe61__lane20_strm1_data        = 'h1234_5678 ;
    std__pe61__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe61__lane21_strm0_cntl        = 'd0         ;
    std__pe61__lane21_strm0_data        = 'h1234_5678 ;
    std__pe61__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe61__lane21_strm1_cntl        = 'd0         ;
    std__pe61__lane21_strm1_data        = 'h1234_5678 ;
    std__pe61__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe61__lane22_strm0_cntl        = 'd0         ;
    std__pe61__lane22_strm0_data        = 'h1234_5678 ;
    std__pe61__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe61__lane22_strm1_cntl        = 'd0         ;
    std__pe61__lane22_strm1_data        = 'h1234_5678 ;
    std__pe61__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe61__lane23_strm0_cntl        = 'd0         ;
    std__pe61__lane23_strm0_data        = 'h1234_5678 ;
    std__pe61__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe61__lane23_strm1_cntl        = 'd0         ;
    std__pe61__lane23_strm1_data        = 'h1234_5678 ;
    std__pe61__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe61__lane24_strm0_cntl        = 'd0         ;
    std__pe61__lane24_strm0_data        = 'h1234_5678 ;
    std__pe61__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe61__lane24_strm1_cntl        = 'd0         ;
    std__pe61__lane24_strm1_data        = 'h1234_5678 ;
    std__pe61__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe61__lane25_strm0_cntl        = 'd0         ;
    std__pe61__lane25_strm0_data        = 'h1234_5678 ;
    std__pe61__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe61__lane25_strm1_cntl        = 'd0         ;
    std__pe61__lane25_strm1_data        = 'h1234_5678 ;
    std__pe61__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe61__lane26_strm0_cntl        = 'd0         ;
    std__pe61__lane26_strm0_data        = 'h1234_5678 ;
    std__pe61__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe61__lane26_strm1_cntl        = 'd0         ;
    std__pe61__lane26_strm1_data        = 'h1234_5678 ;
    std__pe61__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe61__lane27_strm0_cntl        = 'd0         ;
    std__pe61__lane27_strm0_data        = 'h1234_5678 ;
    std__pe61__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe61__lane27_strm1_cntl        = 'd0         ;
    std__pe61__lane27_strm1_data        = 'h1234_5678 ;
    std__pe61__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe61__lane28_strm0_cntl        = 'd0         ;
    std__pe61__lane28_strm0_data        = 'h1234_5678 ;
    std__pe61__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe61__lane28_strm1_cntl        = 'd0         ;
    std__pe61__lane28_strm1_data        = 'h1234_5678 ;
    std__pe61__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe61__lane29_strm0_cntl        = 'd0         ;
    std__pe61__lane29_strm0_data        = 'h1234_5678 ;
    std__pe61__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe61__lane29_strm1_cntl        = 'd0         ;
    std__pe61__lane29_strm1_data        = 'h1234_5678 ;
    std__pe61__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe61__lane30_strm0_cntl        = 'd0         ;
    std__pe61__lane30_strm0_data        = 'h1234_5678 ;
    std__pe61__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe61__lane30_strm1_cntl        = 'd0         ;
    std__pe61__lane30_strm1_data        = 'h1234_5678 ;
    std__pe61__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe61__lane31_strm0_cntl        = 'd0         ;
    std__pe61__lane31_strm0_data        = 'h1234_5678 ;
    std__pe61__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe61__lane31_strm1_cntl        = 'd0         ;
    std__pe61__lane31_strm1_data        = 'h1234_5678 ;
    std__pe61__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe62__lane0_strm0_cntl        = 'd0         ;
    std__pe62__lane0_strm0_data        = 'h1234_5678 ;
    std__pe62__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe62__lane0_strm1_cntl        = 'd0         ;
    std__pe62__lane0_strm1_data        = 'h1234_5678 ;
    std__pe62__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe62__lane1_strm0_cntl        = 'd0         ;
    std__pe62__lane1_strm0_data        = 'h1234_5678 ;
    std__pe62__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe62__lane1_strm1_cntl        = 'd0         ;
    std__pe62__lane1_strm1_data        = 'h1234_5678 ;
    std__pe62__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe62__lane2_strm0_cntl        = 'd0         ;
    std__pe62__lane2_strm0_data        = 'h1234_5678 ;
    std__pe62__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe62__lane2_strm1_cntl        = 'd0         ;
    std__pe62__lane2_strm1_data        = 'h1234_5678 ;
    std__pe62__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe62__lane3_strm0_cntl        = 'd0         ;
    std__pe62__lane3_strm0_data        = 'h1234_5678 ;
    std__pe62__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe62__lane3_strm1_cntl        = 'd0         ;
    std__pe62__lane3_strm1_data        = 'h1234_5678 ;
    std__pe62__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe62__lane4_strm0_cntl        = 'd0         ;
    std__pe62__lane4_strm0_data        = 'h1234_5678 ;
    std__pe62__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe62__lane4_strm1_cntl        = 'd0         ;
    std__pe62__lane4_strm1_data        = 'h1234_5678 ;
    std__pe62__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe62__lane5_strm0_cntl        = 'd0         ;
    std__pe62__lane5_strm0_data        = 'h1234_5678 ;
    std__pe62__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe62__lane5_strm1_cntl        = 'd0         ;
    std__pe62__lane5_strm1_data        = 'h1234_5678 ;
    std__pe62__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe62__lane6_strm0_cntl        = 'd0         ;
    std__pe62__lane6_strm0_data        = 'h1234_5678 ;
    std__pe62__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe62__lane6_strm1_cntl        = 'd0         ;
    std__pe62__lane6_strm1_data        = 'h1234_5678 ;
    std__pe62__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe62__lane7_strm0_cntl        = 'd0         ;
    std__pe62__lane7_strm0_data        = 'h1234_5678 ;
    std__pe62__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe62__lane7_strm1_cntl        = 'd0         ;
    std__pe62__lane7_strm1_data        = 'h1234_5678 ;
    std__pe62__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe62__lane8_strm0_cntl        = 'd0         ;
    std__pe62__lane8_strm0_data        = 'h1234_5678 ;
    std__pe62__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe62__lane8_strm1_cntl        = 'd0         ;
    std__pe62__lane8_strm1_data        = 'h1234_5678 ;
    std__pe62__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe62__lane9_strm0_cntl        = 'd0         ;
    std__pe62__lane9_strm0_data        = 'h1234_5678 ;
    std__pe62__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe62__lane9_strm1_cntl        = 'd0         ;
    std__pe62__lane9_strm1_data        = 'h1234_5678 ;
    std__pe62__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe62__lane10_strm0_cntl        = 'd0         ;
    std__pe62__lane10_strm0_data        = 'h1234_5678 ;
    std__pe62__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe62__lane10_strm1_cntl        = 'd0         ;
    std__pe62__lane10_strm1_data        = 'h1234_5678 ;
    std__pe62__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe62__lane11_strm0_cntl        = 'd0         ;
    std__pe62__lane11_strm0_data        = 'h1234_5678 ;
    std__pe62__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe62__lane11_strm1_cntl        = 'd0         ;
    std__pe62__lane11_strm1_data        = 'h1234_5678 ;
    std__pe62__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe62__lane12_strm0_cntl        = 'd0         ;
    std__pe62__lane12_strm0_data        = 'h1234_5678 ;
    std__pe62__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe62__lane12_strm1_cntl        = 'd0         ;
    std__pe62__lane12_strm1_data        = 'h1234_5678 ;
    std__pe62__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe62__lane13_strm0_cntl        = 'd0         ;
    std__pe62__lane13_strm0_data        = 'h1234_5678 ;
    std__pe62__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe62__lane13_strm1_cntl        = 'd0         ;
    std__pe62__lane13_strm1_data        = 'h1234_5678 ;
    std__pe62__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe62__lane14_strm0_cntl        = 'd0         ;
    std__pe62__lane14_strm0_data        = 'h1234_5678 ;
    std__pe62__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe62__lane14_strm1_cntl        = 'd0         ;
    std__pe62__lane14_strm1_data        = 'h1234_5678 ;
    std__pe62__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe62__lane15_strm0_cntl        = 'd0         ;
    std__pe62__lane15_strm0_data        = 'h1234_5678 ;
    std__pe62__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe62__lane15_strm1_cntl        = 'd0         ;
    std__pe62__lane15_strm1_data        = 'h1234_5678 ;
    std__pe62__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe62__lane16_strm0_cntl        = 'd0         ;
    std__pe62__lane16_strm0_data        = 'h1234_5678 ;
    std__pe62__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe62__lane16_strm1_cntl        = 'd0         ;
    std__pe62__lane16_strm1_data        = 'h1234_5678 ;
    std__pe62__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe62__lane17_strm0_cntl        = 'd0         ;
    std__pe62__lane17_strm0_data        = 'h1234_5678 ;
    std__pe62__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe62__lane17_strm1_cntl        = 'd0         ;
    std__pe62__lane17_strm1_data        = 'h1234_5678 ;
    std__pe62__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe62__lane18_strm0_cntl        = 'd0         ;
    std__pe62__lane18_strm0_data        = 'h1234_5678 ;
    std__pe62__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe62__lane18_strm1_cntl        = 'd0         ;
    std__pe62__lane18_strm1_data        = 'h1234_5678 ;
    std__pe62__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe62__lane19_strm0_cntl        = 'd0         ;
    std__pe62__lane19_strm0_data        = 'h1234_5678 ;
    std__pe62__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe62__lane19_strm1_cntl        = 'd0         ;
    std__pe62__lane19_strm1_data        = 'h1234_5678 ;
    std__pe62__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe62__lane20_strm0_cntl        = 'd0         ;
    std__pe62__lane20_strm0_data        = 'h1234_5678 ;
    std__pe62__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe62__lane20_strm1_cntl        = 'd0         ;
    std__pe62__lane20_strm1_data        = 'h1234_5678 ;
    std__pe62__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe62__lane21_strm0_cntl        = 'd0         ;
    std__pe62__lane21_strm0_data        = 'h1234_5678 ;
    std__pe62__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe62__lane21_strm1_cntl        = 'd0         ;
    std__pe62__lane21_strm1_data        = 'h1234_5678 ;
    std__pe62__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe62__lane22_strm0_cntl        = 'd0         ;
    std__pe62__lane22_strm0_data        = 'h1234_5678 ;
    std__pe62__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe62__lane22_strm1_cntl        = 'd0         ;
    std__pe62__lane22_strm1_data        = 'h1234_5678 ;
    std__pe62__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe62__lane23_strm0_cntl        = 'd0         ;
    std__pe62__lane23_strm0_data        = 'h1234_5678 ;
    std__pe62__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe62__lane23_strm1_cntl        = 'd0         ;
    std__pe62__lane23_strm1_data        = 'h1234_5678 ;
    std__pe62__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe62__lane24_strm0_cntl        = 'd0         ;
    std__pe62__lane24_strm0_data        = 'h1234_5678 ;
    std__pe62__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe62__lane24_strm1_cntl        = 'd0         ;
    std__pe62__lane24_strm1_data        = 'h1234_5678 ;
    std__pe62__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe62__lane25_strm0_cntl        = 'd0         ;
    std__pe62__lane25_strm0_data        = 'h1234_5678 ;
    std__pe62__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe62__lane25_strm1_cntl        = 'd0         ;
    std__pe62__lane25_strm1_data        = 'h1234_5678 ;
    std__pe62__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe62__lane26_strm0_cntl        = 'd0         ;
    std__pe62__lane26_strm0_data        = 'h1234_5678 ;
    std__pe62__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe62__lane26_strm1_cntl        = 'd0         ;
    std__pe62__lane26_strm1_data        = 'h1234_5678 ;
    std__pe62__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe62__lane27_strm0_cntl        = 'd0         ;
    std__pe62__lane27_strm0_data        = 'h1234_5678 ;
    std__pe62__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe62__lane27_strm1_cntl        = 'd0         ;
    std__pe62__lane27_strm1_data        = 'h1234_5678 ;
    std__pe62__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe62__lane28_strm0_cntl        = 'd0         ;
    std__pe62__lane28_strm0_data        = 'h1234_5678 ;
    std__pe62__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe62__lane28_strm1_cntl        = 'd0         ;
    std__pe62__lane28_strm1_data        = 'h1234_5678 ;
    std__pe62__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe62__lane29_strm0_cntl        = 'd0         ;
    std__pe62__lane29_strm0_data        = 'h1234_5678 ;
    std__pe62__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe62__lane29_strm1_cntl        = 'd0         ;
    std__pe62__lane29_strm1_data        = 'h1234_5678 ;
    std__pe62__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe62__lane30_strm0_cntl        = 'd0         ;
    std__pe62__lane30_strm0_data        = 'h1234_5678 ;
    std__pe62__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe62__lane30_strm1_cntl        = 'd0         ;
    std__pe62__lane30_strm1_data        = 'h1234_5678 ;
    std__pe62__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe62__lane31_strm0_cntl        = 'd0         ;
    std__pe62__lane31_strm0_data        = 'h1234_5678 ;
    std__pe62__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe62__lane31_strm1_cntl        = 'd0         ;
    std__pe62__lane31_strm1_data        = 'h1234_5678 ;
    std__pe62__lane31_strm1_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe63__lane0_strm0_cntl        = 'd0         ;
    std__pe63__lane0_strm0_data        = 'h1234_5678 ;
    std__pe63__lane0_strm0_data_valid  = 'd0         ;
    // Lane 0                 
    std__pe63__lane0_strm1_cntl        = 'd0         ;
    std__pe63__lane0_strm1_data        = 'h1234_5678 ;
    std__pe63__lane0_strm1_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe63__lane1_strm0_cntl        = 'd0         ;
    std__pe63__lane1_strm0_data        = 'h1234_5678 ;
    std__pe63__lane1_strm0_data_valid  = 'd0         ;
    // Lane 1                 
    std__pe63__lane1_strm1_cntl        = 'd0         ;
    std__pe63__lane1_strm1_data        = 'h1234_5678 ;
    std__pe63__lane1_strm1_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe63__lane2_strm0_cntl        = 'd0         ;
    std__pe63__lane2_strm0_data        = 'h1234_5678 ;
    std__pe63__lane2_strm0_data_valid  = 'd0         ;
    // Lane 2                 
    std__pe63__lane2_strm1_cntl        = 'd0         ;
    std__pe63__lane2_strm1_data        = 'h1234_5678 ;
    std__pe63__lane2_strm1_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe63__lane3_strm0_cntl        = 'd0         ;
    std__pe63__lane3_strm0_data        = 'h1234_5678 ;
    std__pe63__lane3_strm0_data_valid  = 'd0         ;
    // Lane 3                 
    std__pe63__lane3_strm1_cntl        = 'd0         ;
    std__pe63__lane3_strm1_data        = 'h1234_5678 ;
    std__pe63__lane3_strm1_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe63__lane4_strm0_cntl        = 'd0         ;
    std__pe63__lane4_strm0_data        = 'h1234_5678 ;
    std__pe63__lane4_strm0_data_valid  = 'd0         ;
    // Lane 4                 
    std__pe63__lane4_strm1_cntl        = 'd0         ;
    std__pe63__lane4_strm1_data        = 'h1234_5678 ;
    std__pe63__lane4_strm1_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe63__lane5_strm0_cntl        = 'd0         ;
    std__pe63__lane5_strm0_data        = 'h1234_5678 ;
    std__pe63__lane5_strm0_data_valid  = 'd0         ;
    // Lane 5                 
    std__pe63__lane5_strm1_cntl        = 'd0         ;
    std__pe63__lane5_strm1_data        = 'h1234_5678 ;
    std__pe63__lane5_strm1_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe63__lane6_strm0_cntl        = 'd0         ;
    std__pe63__lane6_strm0_data        = 'h1234_5678 ;
    std__pe63__lane6_strm0_data_valid  = 'd0         ;
    // Lane 6                 
    std__pe63__lane6_strm1_cntl        = 'd0         ;
    std__pe63__lane6_strm1_data        = 'h1234_5678 ;
    std__pe63__lane6_strm1_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe63__lane7_strm0_cntl        = 'd0         ;
    std__pe63__lane7_strm0_data        = 'h1234_5678 ;
    std__pe63__lane7_strm0_data_valid  = 'd0         ;
    // Lane 7                 
    std__pe63__lane7_strm1_cntl        = 'd0         ;
    std__pe63__lane7_strm1_data        = 'h1234_5678 ;
    std__pe63__lane7_strm1_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe63__lane8_strm0_cntl        = 'd0         ;
    std__pe63__lane8_strm0_data        = 'h1234_5678 ;
    std__pe63__lane8_strm0_data_valid  = 'd0         ;
    // Lane 8                 
    std__pe63__lane8_strm1_cntl        = 'd0         ;
    std__pe63__lane8_strm1_data        = 'h1234_5678 ;
    std__pe63__lane8_strm1_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe63__lane9_strm0_cntl        = 'd0         ;
    std__pe63__lane9_strm0_data        = 'h1234_5678 ;
    std__pe63__lane9_strm0_data_valid  = 'd0         ;
    // Lane 9                 
    std__pe63__lane9_strm1_cntl        = 'd0         ;
    std__pe63__lane9_strm1_data        = 'h1234_5678 ;
    std__pe63__lane9_strm1_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe63__lane10_strm0_cntl        = 'd0         ;
    std__pe63__lane10_strm0_data        = 'h1234_5678 ;
    std__pe63__lane10_strm0_data_valid  = 'd0         ;
    // Lane 10                 
    std__pe63__lane10_strm1_cntl        = 'd0         ;
    std__pe63__lane10_strm1_data        = 'h1234_5678 ;
    std__pe63__lane10_strm1_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe63__lane11_strm0_cntl        = 'd0         ;
    std__pe63__lane11_strm0_data        = 'h1234_5678 ;
    std__pe63__lane11_strm0_data_valid  = 'd0         ;
    // Lane 11                 
    std__pe63__lane11_strm1_cntl        = 'd0         ;
    std__pe63__lane11_strm1_data        = 'h1234_5678 ;
    std__pe63__lane11_strm1_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe63__lane12_strm0_cntl        = 'd0         ;
    std__pe63__lane12_strm0_data        = 'h1234_5678 ;
    std__pe63__lane12_strm0_data_valid  = 'd0         ;
    // Lane 12                 
    std__pe63__lane12_strm1_cntl        = 'd0         ;
    std__pe63__lane12_strm1_data        = 'h1234_5678 ;
    std__pe63__lane12_strm1_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe63__lane13_strm0_cntl        = 'd0         ;
    std__pe63__lane13_strm0_data        = 'h1234_5678 ;
    std__pe63__lane13_strm0_data_valid  = 'd0         ;
    // Lane 13                 
    std__pe63__lane13_strm1_cntl        = 'd0         ;
    std__pe63__lane13_strm1_data        = 'h1234_5678 ;
    std__pe63__lane13_strm1_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe63__lane14_strm0_cntl        = 'd0         ;
    std__pe63__lane14_strm0_data        = 'h1234_5678 ;
    std__pe63__lane14_strm0_data_valid  = 'd0         ;
    // Lane 14                 
    std__pe63__lane14_strm1_cntl        = 'd0         ;
    std__pe63__lane14_strm1_data        = 'h1234_5678 ;
    std__pe63__lane14_strm1_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe63__lane15_strm0_cntl        = 'd0         ;
    std__pe63__lane15_strm0_data        = 'h1234_5678 ;
    std__pe63__lane15_strm0_data_valid  = 'd0         ;
    // Lane 15                 
    std__pe63__lane15_strm1_cntl        = 'd0         ;
    std__pe63__lane15_strm1_data        = 'h1234_5678 ;
    std__pe63__lane15_strm1_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe63__lane16_strm0_cntl        = 'd0         ;
    std__pe63__lane16_strm0_data        = 'h1234_5678 ;
    std__pe63__lane16_strm0_data_valid  = 'd0         ;
    // Lane 16                 
    std__pe63__lane16_strm1_cntl        = 'd0         ;
    std__pe63__lane16_strm1_data        = 'h1234_5678 ;
    std__pe63__lane16_strm1_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe63__lane17_strm0_cntl        = 'd0         ;
    std__pe63__lane17_strm0_data        = 'h1234_5678 ;
    std__pe63__lane17_strm0_data_valid  = 'd0         ;
    // Lane 17                 
    std__pe63__lane17_strm1_cntl        = 'd0         ;
    std__pe63__lane17_strm1_data        = 'h1234_5678 ;
    std__pe63__lane17_strm1_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe63__lane18_strm0_cntl        = 'd0         ;
    std__pe63__lane18_strm0_data        = 'h1234_5678 ;
    std__pe63__lane18_strm0_data_valid  = 'd0         ;
    // Lane 18                 
    std__pe63__lane18_strm1_cntl        = 'd0         ;
    std__pe63__lane18_strm1_data        = 'h1234_5678 ;
    std__pe63__lane18_strm1_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe63__lane19_strm0_cntl        = 'd0         ;
    std__pe63__lane19_strm0_data        = 'h1234_5678 ;
    std__pe63__lane19_strm0_data_valid  = 'd0         ;
    // Lane 19                 
    std__pe63__lane19_strm1_cntl        = 'd0         ;
    std__pe63__lane19_strm1_data        = 'h1234_5678 ;
    std__pe63__lane19_strm1_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe63__lane20_strm0_cntl        = 'd0         ;
    std__pe63__lane20_strm0_data        = 'h1234_5678 ;
    std__pe63__lane20_strm0_data_valid  = 'd0         ;
    // Lane 20                 
    std__pe63__lane20_strm1_cntl        = 'd0         ;
    std__pe63__lane20_strm1_data        = 'h1234_5678 ;
    std__pe63__lane20_strm1_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe63__lane21_strm0_cntl        = 'd0         ;
    std__pe63__lane21_strm0_data        = 'h1234_5678 ;
    std__pe63__lane21_strm0_data_valid  = 'd0         ;
    // Lane 21                 
    std__pe63__lane21_strm1_cntl        = 'd0         ;
    std__pe63__lane21_strm1_data        = 'h1234_5678 ;
    std__pe63__lane21_strm1_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe63__lane22_strm0_cntl        = 'd0         ;
    std__pe63__lane22_strm0_data        = 'h1234_5678 ;
    std__pe63__lane22_strm0_data_valid  = 'd0         ;
    // Lane 22                 
    std__pe63__lane22_strm1_cntl        = 'd0         ;
    std__pe63__lane22_strm1_data        = 'h1234_5678 ;
    std__pe63__lane22_strm1_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe63__lane23_strm0_cntl        = 'd0         ;
    std__pe63__lane23_strm0_data        = 'h1234_5678 ;
    std__pe63__lane23_strm0_data_valid  = 'd0         ;
    // Lane 23                 
    std__pe63__lane23_strm1_cntl        = 'd0         ;
    std__pe63__lane23_strm1_data        = 'h1234_5678 ;
    std__pe63__lane23_strm1_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe63__lane24_strm0_cntl        = 'd0         ;
    std__pe63__lane24_strm0_data        = 'h1234_5678 ;
    std__pe63__lane24_strm0_data_valid  = 'd0         ;
    // Lane 24                 
    std__pe63__lane24_strm1_cntl        = 'd0         ;
    std__pe63__lane24_strm1_data        = 'h1234_5678 ;
    std__pe63__lane24_strm1_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe63__lane25_strm0_cntl        = 'd0         ;
    std__pe63__lane25_strm0_data        = 'h1234_5678 ;
    std__pe63__lane25_strm0_data_valid  = 'd0         ;
    // Lane 25                 
    std__pe63__lane25_strm1_cntl        = 'd0         ;
    std__pe63__lane25_strm1_data        = 'h1234_5678 ;
    std__pe63__lane25_strm1_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe63__lane26_strm0_cntl        = 'd0         ;
    std__pe63__lane26_strm0_data        = 'h1234_5678 ;
    std__pe63__lane26_strm0_data_valid  = 'd0         ;
    // Lane 26                 
    std__pe63__lane26_strm1_cntl        = 'd0         ;
    std__pe63__lane26_strm1_data        = 'h1234_5678 ;
    std__pe63__lane26_strm1_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe63__lane27_strm0_cntl        = 'd0         ;
    std__pe63__lane27_strm0_data        = 'h1234_5678 ;
    std__pe63__lane27_strm0_data_valid  = 'd0         ;
    // Lane 27                 
    std__pe63__lane27_strm1_cntl        = 'd0         ;
    std__pe63__lane27_strm1_data        = 'h1234_5678 ;
    std__pe63__lane27_strm1_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe63__lane28_strm0_cntl        = 'd0         ;
    std__pe63__lane28_strm0_data        = 'h1234_5678 ;
    std__pe63__lane28_strm0_data_valid  = 'd0         ;
    // Lane 28                 
    std__pe63__lane28_strm1_cntl        = 'd0         ;
    std__pe63__lane28_strm1_data        = 'h1234_5678 ;
    std__pe63__lane28_strm1_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe63__lane29_strm0_cntl        = 'd0         ;
    std__pe63__lane29_strm0_data        = 'h1234_5678 ;
    std__pe63__lane29_strm0_data_valid  = 'd0         ;
    // Lane 29                 
    std__pe63__lane29_strm1_cntl        = 'd0         ;
    std__pe63__lane29_strm1_data        = 'h1234_5678 ;
    std__pe63__lane29_strm1_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe63__lane30_strm0_cntl        = 'd0         ;
    std__pe63__lane30_strm0_data        = 'h1234_5678 ;
    std__pe63__lane30_strm0_data_valid  = 'd0         ;
    // Lane 30                 
    std__pe63__lane30_strm1_cntl        = 'd0         ;
    std__pe63__lane30_strm1_data        = 'h1234_5678 ;
    std__pe63__lane30_strm1_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe63__lane31_strm0_cntl        = 'd0         ;
    std__pe63__lane31_strm0_data        = 'h1234_5678 ;
    std__pe63__lane31_strm0_data_valid  = 'd0         ;
    // Lane 31                 
    std__pe63__lane31_strm1_cntl        = 'd0         ;
    std__pe63__lane31_strm1_data        = 'h1234_5678 ;
    std__pe63__lane31_strm1_data_valid  = 'd0         ;