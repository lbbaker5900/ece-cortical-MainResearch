
    // PE0, Port0 next hop mask                 
    assign pe_inst[0].sys__pe__port0_destinationMask    = `NOC_CONT_PE0_PORT0_DESTINATION_PE_BITMASK ;
    // PE0, Port1 next hop mask                 
    assign pe_inst[0].sys__pe__port1_destinationMask    = `NOC_CONT_PE0_PORT1_DESTINATION_PE_BITMASK ;
    // PE0, Port2 next hop mask                 
    assign pe_inst[0].sys__pe__port2_destinationMask    = `NOC_CONT_PE0_PORT2_DESTINATION_PE_BITMASK ;
    // PE0, Port3 next hop mask                 
    assign pe_inst[0].sys__pe__port3_destinationMask    = `NOC_CONT_PE0_PORT3_DESTINATION_PE_BITMASK ;
    // PE1, Port0 next hop mask                 
    assign pe_inst[1].sys__pe__port0_destinationMask    = `NOC_CONT_PE1_PORT0_DESTINATION_PE_BITMASK ;
    // PE1, Port1 next hop mask                 
    assign pe_inst[1].sys__pe__port1_destinationMask    = `NOC_CONT_PE1_PORT1_DESTINATION_PE_BITMASK ;
    // PE1, Port2 next hop mask                 
    assign pe_inst[1].sys__pe__port2_destinationMask    = `NOC_CONT_PE1_PORT2_DESTINATION_PE_BITMASK ;
    // PE1, Port3 next hop mask                 
    assign pe_inst[1].sys__pe__port3_destinationMask    = `NOC_CONT_PE1_PORT3_DESTINATION_PE_BITMASK ;
    // PE2, Port0 next hop mask                 
    assign pe_inst[2].sys__pe__port0_destinationMask    = `NOC_CONT_PE2_PORT0_DESTINATION_PE_BITMASK ;
    // PE2, Port1 next hop mask                 
    assign pe_inst[2].sys__pe__port1_destinationMask    = `NOC_CONT_PE2_PORT1_DESTINATION_PE_BITMASK ;
    // PE2, Port2 next hop mask                 
    assign pe_inst[2].sys__pe__port2_destinationMask    = `NOC_CONT_PE2_PORT2_DESTINATION_PE_BITMASK ;
    // PE2, Port3 next hop mask                 
    assign pe_inst[2].sys__pe__port3_destinationMask    = `NOC_CONT_PE2_PORT3_DESTINATION_PE_BITMASK ;
    // PE3, Port0 next hop mask                 
    assign pe_inst[3].sys__pe__port0_destinationMask    = `NOC_CONT_PE3_PORT0_DESTINATION_PE_BITMASK ;
    // PE3, Port1 next hop mask                 
    assign pe_inst[3].sys__pe__port1_destinationMask    = `NOC_CONT_PE3_PORT1_DESTINATION_PE_BITMASK ;
    // PE3, Port2 next hop mask                 
    assign pe_inst[3].sys__pe__port2_destinationMask    = `NOC_CONT_PE3_PORT2_DESTINATION_PE_BITMASK ;
    // PE3, Port3 next hop mask                 
    assign pe_inst[3].sys__pe__port3_destinationMask    = `NOC_CONT_PE3_PORT3_DESTINATION_PE_BITMASK ;
    // PE4, Port0 next hop mask                 
    assign pe_inst[4].sys__pe__port0_destinationMask    = `NOC_CONT_PE4_PORT0_DESTINATION_PE_BITMASK ;
    // PE4, Port1 next hop mask                 
    assign pe_inst[4].sys__pe__port1_destinationMask    = `NOC_CONT_PE4_PORT1_DESTINATION_PE_BITMASK ;
    // PE4, Port2 next hop mask                 
    assign pe_inst[4].sys__pe__port2_destinationMask    = `NOC_CONT_PE4_PORT2_DESTINATION_PE_BITMASK ;
    // PE4, Port3 next hop mask                 
    assign pe_inst[4].sys__pe__port3_destinationMask    = `NOC_CONT_PE4_PORT3_DESTINATION_PE_BITMASK ;
    // PE5, Port0 next hop mask                 
    assign pe_inst[5].sys__pe__port0_destinationMask    = `NOC_CONT_PE5_PORT0_DESTINATION_PE_BITMASK ;
    // PE5, Port1 next hop mask                 
    assign pe_inst[5].sys__pe__port1_destinationMask    = `NOC_CONT_PE5_PORT1_DESTINATION_PE_BITMASK ;
    // PE5, Port2 next hop mask                 
    assign pe_inst[5].sys__pe__port2_destinationMask    = `NOC_CONT_PE5_PORT2_DESTINATION_PE_BITMASK ;
    // PE5, Port3 next hop mask                 
    assign pe_inst[5].sys__pe__port3_destinationMask    = `NOC_CONT_PE5_PORT3_DESTINATION_PE_BITMASK ;
    // PE6, Port0 next hop mask                 
    assign pe_inst[6].sys__pe__port0_destinationMask    = `NOC_CONT_PE6_PORT0_DESTINATION_PE_BITMASK ;
    // PE6, Port1 next hop mask                 
    assign pe_inst[6].sys__pe__port1_destinationMask    = `NOC_CONT_PE6_PORT1_DESTINATION_PE_BITMASK ;
    // PE6, Port2 next hop mask                 
    assign pe_inst[6].sys__pe__port2_destinationMask    = `NOC_CONT_PE6_PORT2_DESTINATION_PE_BITMASK ;
    // PE6, Port3 next hop mask                 
    assign pe_inst[6].sys__pe__port3_destinationMask    = `NOC_CONT_PE6_PORT3_DESTINATION_PE_BITMASK ;
    // PE7, Port0 next hop mask                 
    assign pe_inst[7].sys__pe__port0_destinationMask    = `NOC_CONT_PE7_PORT0_DESTINATION_PE_BITMASK ;
    // PE7, Port1 next hop mask                 
    assign pe_inst[7].sys__pe__port1_destinationMask    = `NOC_CONT_PE7_PORT1_DESTINATION_PE_BITMASK ;
    // PE7, Port2 next hop mask                 
    assign pe_inst[7].sys__pe__port2_destinationMask    = `NOC_CONT_PE7_PORT2_DESTINATION_PE_BITMASK ;
    // PE7, Port3 next hop mask                 
    assign pe_inst[7].sys__pe__port3_destinationMask    = `NOC_CONT_PE7_PORT3_DESTINATION_PE_BITMASK ;
    // PE8, Port0 next hop mask                 
    assign pe_inst[8].sys__pe__port0_destinationMask    = `NOC_CONT_PE8_PORT0_DESTINATION_PE_BITMASK ;
    // PE8, Port1 next hop mask                 
    assign pe_inst[8].sys__pe__port1_destinationMask    = `NOC_CONT_PE8_PORT1_DESTINATION_PE_BITMASK ;
    // PE8, Port2 next hop mask                 
    assign pe_inst[8].sys__pe__port2_destinationMask    = `NOC_CONT_PE8_PORT2_DESTINATION_PE_BITMASK ;
    // PE8, Port3 next hop mask                 
    assign pe_inst[8].sys__pe__port3_destinationMask    = `NOC_CONT_PE8_PORT3_DESTINATION_PE_BITMASK ;
    // PE9, Port0 next hop mask                 
    assign pe_inst[9].sys__pe__port0_destinationMask    = `NOC_CONT_PE9_PORT0_DESTINATION_PE_BITMASK ;
    // PE9, Port1 next hop mask                 
    assign pe_inst[9].sys__pe__port1_destinationMask    = `NOC_CONT_PE9_PORT1_DESTINATION_PE_BITMASK ;
    // PE9, Port2 next hop mask                 
    assign pe_inst[9].sys__pe__port2_destinationMask    = `NOC_CONT_PE9_PORT2_DESTINATION_PE_BITMASK ;
    // PE9, Port3 next hop mask                 
    assign pe_inst[9].sys__pe__port3_destinationMask    = `NOC_CONT_PE9_PORT3_DESTINATION_PE_BITMASK ;
    // PE10, Port0 next hop mask                 
    assign pe_inst[10].sys__pe__port0_destinationMask    = `NOC_CONT_PE10_PORT0_DESTINATION_PE_BITMASK ;
    // PE10, Port1 next hop mask                 
    assign pe_inst[10].sys__pe__port1_destinationMask    = `NOC_CONT_PE10_PORT1_DESTINATION_PE_BITMASK ;
    // PE10, Port2 next hop mask                 
    assign pe_inst[10].sys__pe__port2_destinationMask    = `NOC_CONT_PE10_PORT2_DESTINATION_PE_BITMASK ;
    // PE10, Port3 next hop mask                 
    assign pe_inst[10].sys__pe__port3_destinationMask    = `NOC_CONT_PE10_PORT3_DESTINATION_PE_BITMASK ;
    // PE11, Port0 next hop mask                 
    assign pe_inst[11].sys__pe__port0_destinationMask    = `NOC_CONT_PE11_PORT0_DESTINATION_PE_BITMASK ;
    // PE11, Port1 next hop mask                 
    assign pe_inst[11].sys__pe__port1_destinationMask    = `NOC_CONT_PE11_PORT1_DESTINATION_PE_BITMASK ;
    // PE11, Port2 next hop mask                 
    assign pe_inst[11].sys__pe__port2_destinationMask    = `NOC_CONT_PE11_PORT2_DESTINATION_PE_BITMASK ;
    // PE11, Port3 next hop mask                 
    assign pe_inst[11].sys__pe__port3_destinationMask    = `NOC_CONT_PE11_PORT3_DESTINATION_PE_BITMASK ;
    // PE12, Port0 next hop mask                 
    assign pe_inst[12].sys__pe__port0_destinationMask    = `NOC_CONT_PE12_PORT0_DESTINATION_PE_BITMASK ;
    // PE12, Port1 next hop mask                 
    assign pe_inst[12].sys__pe__port1_destinationMask    = `NOC_CONT_PE12_PORT1_DESTINATION_PE_BITMASK ;
    // PE12, Port2 next hop mask                 
    assign pe_inst[12].sys__pe__port2_destinationMask    = `NOC_CONT_PE12_PORT2_DESTINATION_PE_BITMASK ;
    // PE12, Port3 next hop mask                 
    assign pe_inst[12].sys__pe__port3_destinationMask    = `NOC_CONT_PE12_PORT3_DESTINATION_PE_BITMASK ;
    // PE13, Port0 next hop mask                 
    assign pe_inst[13].sys__pe__port0_destinationMask    = `NOC_CONT_PE13_PORT0_DESTINATION_PE_BITMASK ;
    // PE13, Port1 next hop mask                 
    assign pe_inst[13].sys__pe__port1_destinationMask    = `NOC_CONT_PE13_PORT1_DESTINATION_PE_BITMASK ;
    // PE13, Port2 next hop mask                 
    assign pe_inst[13].sys__pe__port2_destinationMask    = `NOC_CONT_PE13_PORT2_DESTINATION_PE_BITMASK ;
    // PE13, Port3 next hop mask                 
    assign pe_inst[13].sys__pe__port3_destinationMask    = `NOC_CONT_PE13_PORT3_DESTINATION_PE_BITMASK ;
    // PE14, Port0 next hop mask                 
    assign pe_inst[14].sys__pe__port0_destinationMask    = `NOC_CONT_PE14_PORT0_DESTINATION_PE_BITMASK ;
    // PE14, Port1 next hop mask                 
    assign pe_inst[14].sys__pe__port1_destinationMask    = `NOC_CONT_PE14_PORT1_DESTINATION_PE_BITMASK ;
    // PE14, Port2 next hop mask                 
    assign pe_inst[14].sys__pe__port2_destinationMask    = `NOC_CONT_PE14_PORT2_DESTINATION_PE_BITMASK ;
    // PE14, Port3 next hop mask                 
    assign pe_inst[14].sys__pe__port3_destinationMask    = `NOC_CONT_PE14_PORT3_DESTINATION_PE_BITMASK ;
    // PE15, Port0 next hop mask                 
    assign pe_inst[15].sys__pe__port0_destinationMask    = `NOC_CONT_PE15_PORT0_DESTINATION_PE_BITMASK ;
    // PE15, Port1 next hop mask                 
    assign pe_inst[15].sys__pe__port1_destinationMask    = `NOC_CONT_PE15_PORT1_DESTINATION_PE_BITMASK ;
    // PE15, Port2 next hop mask                 
    assign pe_inst[15].sys__pe__port2_destinationMask    = `NOC_CONT_PE15_PORT2_DESTINATION_PE_BITMASK ;
    // PE15, Port3 next hop mask                 
    assign pe_inst[15].sys__pe__port3_destinationMask    = `NOC_CONT_PE15_PORT3_DESTINATION_PE_BITMASK ;
    // PE16, Port0 next hop mask                 
    assign pe_inst[16].sys__pe__port0_destinationMask    = `NOC_CONT_PE16_PORT0_DESTINATION_PE_BITMASK ;
    // PE16, Port1 next hop mask                 
    assign pe_inst[16].sys__pe__port1_destinationMask    = `NOC_CONT_PE16_PORT1_DESTINATION_PE_BITMASK ;
    // PE16, Port2 next hop mask                 
    assign pe_inst[16].sys__pe__port2_destinationMask    = `NOC_CONT_PE16_PORT2_DESTINATION_PE_BITMASK ;
    // PE16, Port3 next hop mask                 
    assign pe_inst[16].sys__pe__port3_destinationMask    = `NOC_CONT_PE16_PORT3_DESTINATION_PE_BITMASK ;
    // PE17, Port0 next hop mask                 
    assign pe_inst[17].sys__pe__port0_destinationMask    = `NOC_CONT_PE17_PORT0_DESTINATION_PE_BITMASK ;
    // PE17, Port1 next hop mask                 
    assign pe_inst[17].sys__pe__port1_destinationMask    = `NOC_CONT_PE17_PORT1_DESTINATION_PE_BITMASK ;
    // PE17, Port2 next hop mask                 
    assign pe_inst[17].sys__pe__port2_destinationMask    = `NOC_CONT_PE17_PORT2_DESTINATION_PE_BITMASK ;
    // PE17, Port3 next hop mask                 
    assign pe_inst[17].sys__pe__port3_destinationMask    = `NOC_CONT_PE17_PORT3_DESTINATION_PE_BITMASK ;
    // PE18, Port0 next hop mask                 
    assign pe_inst[18].sys__pe__port0_destinationMask    = `NOC_CONT_PE18_PORT0_DESTINATION_PE_BITMASK ;
    // PE18, Port1 next hop mask                 
    assign pe_inst[18].sys__pe__port1_destinationMask    = `NOC_CONT_PE18_PORT1_DESTINATION_PE_BITMASK ;
    // PE18, Port2 next hop mask                 
    assign pe_inst[18].sys__pe__port2_destinationMask    = `NOC_CONT_PE18_PORT2_DESTINATION_PE_BITMASK ;
    // PE18, Port3 next hop mask                 
    assign pe_inst[18].sys__pe__port3_destinationMask    = `NOC_CONT_PE18_PORT3_DESTINATION_PE_BITMASK ;
    // PE19, Port0 next hop mask                 
    assign pe_inst[19].sys__pe__port0_destinationMask    = `NOC_CONT_PE19_PORT0_DESTINATION_PE_BITMASK ;
    // PE19, Port1 next hop mask                 
    assign pe_inst[19].sys__pe__port1_destinationMask    = `NOC_CONT_PE19_PORT1_DESTINATION_PE_BITMASK ;
    // PE19, Port2 next hop mask                 
    assign pe_inst[19].sys__pe__port2_destinationMask    = `NOC_CONT_PE19_PORT2_DESTINATION_PE_BITMASK ;
    // PE19, Port3 next hop mask                 
    assign pe_inst[19].sys__pe__port3_destinationMask    = `NOC_CONT_PE19_PORT3_DESTINATION_PE_BITMASK ;
    // PE20, Port0 next hop mask                 
    assign pe_inst[20].sys__pe__port0_destinationMask    = `NOC_CONT_PE20_PORT0_DESTINATION_PE_BITMASK ;
    // PE20, Port1 next hop mask                 
    assign pe_inst[20].sys__pe__port1_destinationMask    = `NOC_CONT_PE20_PORT1_DESTINATION_PE_BITMASK ;
    // PE20, Port2 next hop mask                 
    assign pe_inst[20].sys__pe__port2_destinationMask    = `NOC_CONT_PE20_PORT2_DESTINATION_PE_BITMASK ;
    // PE20, Port3 next hop mask                 
    assign pe_inst[20].sys__pe__port3_destinationMask    = `NOC_CONT_PE20_PORT3_DESTINATION_PE_BITMASK ;
    // PE21, Port0 next hop mask                 
    assign pe_inst[21].sys__pe__port0_destinationMask    = `NOC_CONT_PE21_PORT0_DESTINATION_PE_BITMASK ;
    // PE21, Port1 next hop mask                 
    assign pe_inst[21].sys__pe__port1_destinationMask    = `NOC_CONT_PE21_PORT1_DESTINATION_PE_BITMASK ;
    // PE21, Port2 next hop mask                 
    assign pe_inst[21].sys__pe__port2_destinationMask    = `NOC_CONT_PE21_PORT2_DESTINATION_PE_BITMASK ;
    // PE21, Port3 next hop mask                 
    assign pe_inst[21].sys__pe__port3_destinationMask    = `NOC_CONT_PE21_PORT3_DESTINATION_PE_BITMASK ;
    // PE22, Port0 next hop mask                 
    assign pe_inst[22].sys__pe__port0_destinationMask    = `NOC_CONT_PE22_PORT0_DESTINATION_PE_BITMASK ;
    // PE22, Port1 next hop mask                 
    assign pe_inst[22].sys__pe__port1_destinationMask    = `NOC_CONT_PE22_PORT1_DESTINATION_PE_BITMASK ;
    // PE22, Port2 next hop mask                 
    assign pe_inst[22].sys__pe__port2_destinationMask    = `NOC_CONT_PE22_PORT2_DESTINATION_PE_BITMASK ;
    // PE22, Port3 next hop mask                 
    assign pe_inst[22].sys__pe__port3_destinationMask    = `NOC_CONT_PE22_PORT3_DESTINATION_PE_BITMASK ;
    // PE23, Port0 next hop mask                 
    assign pe_inst[23].sys__pe__port0_destinationMask    = `NOC_CONT_PE23_PORT0_DESTINATION_PE_BITMASK ;
    // PE23, Port1 next hop mask                 
    assign pe_inst[23].sys__pe__port1_destinationMask    = `NOC_CONT_PE23_PORT1_DESTINATION_PE_BITMASK ;
    // PE23, Port2 next hop mask                 
    assign pe_inst[23].sys__pe__port2_destinationMask    = `NOC_CONT_PE23_PORT2_DESTINATION_PE_BITMASK ;
    // PE23, Port3 next hop mask                 
    assign pe_inst[23].sys__pe__port3_destinationMask    = `NOC_CONT_PE23_PORT3_DESTINATION_PE_BITMASK ;
    // PE24, Port0 next hop mask                 
    assign pe_inst[24].sys__pe__port0_destinationMask    = `NOC_CONT_PE24_PORT0_DESTINATION_PE_BITMASK ;
    // PE24, Port1 next hop mask                 
    assign pe_inst[24].sys__pe__port1_destinationMask    = `NOC_CONT_PE24_PORT1_DESTINATION_PE_BITMASK ;
    // PE24, Port2 next hop mask                 
    assign pe_inst[24].sys__pe__port2_destinationMask    = `NOC_CONT_PE24_PORT2_DESTINATION_PE_BITMASK ;
    // PE24, Port3 next hop mask                 
    assign pe_inst[24].sys__pe__port3_destinationMask    = `NOC_CONT_PE24_PORT3_DESTINATION_PE_BITMASK ;
    // PE25, Port0 next hop mask                 
    assign pe_inst[25].sys__pe__port0_destinationMask    = `NOC_CONT_PE25_PORT0_DESTINATION_PE_BITMASK ;
    // PE25, Port1 next hop mask                 
    assign pe_inst[25].sys__pe__port1_destinationMask    = `NOC_CONT_PE25_PORT1_DESTINATION_PE_BITMASK ;
    // PE25, Port2 next hop mask                 
    assign pe_inst[25].sys__pe__port2_destinationMask    = `NOC_CONT_PE25_PORT2_DESTINATION_PE_BITMASK ;
    // PE25, Port3 next hop mask                 
    assign pe_inst[25].sys__pe__port3_destinationMask    = `NOC_CONT_PE25_PORT3_DESTINATION_PE_BITMASK ;
    // PE26, Port0 next hop mask                 
    assign pe_inst[26].sys__pe__port0_destinationMask    = `NOC_CONT_PE26_PORT0_DESTINATION_PE_BITMASK ;
    // PE26, Port1 next hop mask                 
    assign pe_inst[26].sys__pe__port1_destinationMask    = `NOC_CONT_PE26_PORT1_DESTINATION_PE_BITMASK ;
    // PE26, Port2 next hop mask                 
    assign pe_inst[26].sys__pe__port2_destinationMask    = `NOC_CONT_PE26_PORT2_DESTINATION_PE_BITMASK ;
    // PE26, Port3 next hop mask                 
    assign pe_inst[26].sys__pe__port3_destinationMask    = `NOC_CONT_PE26_PORT3_DESTINATION_PE_BITMASK ;
    // PE27, Port0 next hop mask                 
    assign pe_inst[27].sys__pe__port0_destinationMask    = `NOC_CONT_PE27_PORT0_DESTINATION_PE_BITMASK ;
    // PE27, Port1 next hop mask                 
    assign pe_inst[27].sys__pe__port1_destinationMask    = `NOC_CONT_PE27_PORT1_DESTINATION_PE_BITMASK ;
    // PE27, Port2 next hop mask                 
    assign pe_inst[27].sys__pe__port2_destinationMask    = `NOC_CONT_PE27_PORT2_DESTINATION_PE_BITMASK ;
    // PE27, Port3 next hop mask                 
    assign pe_inst[27].sys__pe__port3_destinationMask    = `NOC_CONT_PE27_PORT3_DESTINATION_PE_BITMASK ;
    // PE28, Port0 next hop mask                 
    assign pe_inst[28].sys__pe__port0_destinationMask    = `NOC_CONT_PE28_PORT0_DESTINATION_PE_BITMASK ;
    // PE28, Port1 next hop mask                 
    assign pe_inst[28].sys__pe__port1_destinationMask    = `NOC_CONT_PE28_PORT1_DESTINATION_PE_BITMASK ;
    // PE28, Port2 next hop mask                 
    assign pe_inst[28].sys__pe__port2_destinationMask    = `NOC_CONT_PE28_PORT2_DESTINATION_PE_BITMASK ;
    // PE28, Port3 next hop mask                 
    assign pe_inst[28].sys__pe__port3_destinationMask    = `NOC_CONT_PE28_PORT3_DESTINATION_PE_BITMASK ;
    // PE29, Port0 next hop mask                 
    assign pe_inst[29].sys__pe__port0_destinationMask    = `NOC_CONT_PE29_PORT0_DESTINATION_PE_BITMASK ;
    // PE29, Port1 next hop mask                 
    assign pe_inst[29].sys__pe__port1_destinationMask    = `NOC_CONT_PE29_PORT1_DESTINATION_PE_BITMASK ;
    // PE29, Port2 next hop mask                 
    assign pe_inst[29].sys__pe__port2_destinationMask    = `NOC_CONT_PE29_PORT2_DESTINATION_PE_BITMASK ;
    // PE29, Port3 next hop mask                 
    assign pe_inst[29].sys__pe__port3_destinationMask    = `NOC_CONT_PE29_PORT3_DESTINATION_PE_BITMASK ;
    // PE30, Port0 next hop mask                 
    assign pe_inst[30].sys__pe__port0_destinationMask    = `NOC_CONT_PE30_PORT0_DESTINATION_PE_BITMASK ;
    // PE30, Port1 next hop mask                 
    assign pe_inst[30].sys__pe__port1_destinationMask    = `NOC_CONT_PE30_PORT1_DESTINATION_PE_BITMASK ;
    // PE30, Port2 next hop mask                 
    assign pe_inst[30].sys__pe__port2_destinationMask    = `NOC_CONT_PE30_PORT2_DESTINATION_PE_BITMASK ;
    // PE30, Port3 next hop mask                 
    assign pe_inst[30].sys__pe__port3_destinationMask    = `NOC_CONT_PE30_PORT3_DESTINATION_PE_BITMASK ;
    // PE31, Port0 next hop mask                 
    assign pe_inst[31].sys__pe__port0_destinationMask    = `NOC_CONT_PE31_PORT0_DESTINATION_PE_BITMASK ;
    // PE31, Port1 next hop mask                 
    assign pe_inst[31].sys__pe__port1_destinationMask    = `NOC_CONT_PE31_PORT1_DESTINATION_PE_BITMASK ;
    // PE31, Port2 next hop mask                 
    assign pe_inst[31].sys__pe__port2_destinationMask    = `NOC_CONT_PE31_PORT2_DESTINATION_PE_BITMASK ;
    // PE31, Port3 next hop mask                 
    assign pe_inst[31].sys__pe__port3_destinationMask    = `NOC_CONT_PE31_PORT3_DESTINATION_PE_BITMASK ;
    // PE32, Port0 next hop mask                 
    assign pe_inst[32].sys__pe__port0_destinationMask    = `NOC_CONT_PE32_PORT0_DESTINATION_PE_BITMASK ;
    // PE32, Port1 next hop mask                 
    assign pe_inst[32].sys__pe__port1_destinationMask    = `NOC_CONT_PE32_PORT1_DESTINATION_PE_BITMASK ;
    // PE32, Port2 next hop mask                 
    assign pe_inst[32].sys__pe__port2_destinationMask    = `NOC_CONT_PE32_PORT2_DESTINATION_PE_BITMASK ;
    // PE32, Port3 next hop mask                 
    assign pe_inst[32].sys__pe__port3_destinationMask    = `NOC_CONT_PE32_PORT3_DESTINATION_PE_BITMASK ;
    // PE33, Port0 next hop mask                 
    assign pe_inst[33].sys__pe__port0_destinationMask    = `NOC_CONT_PE33_PORT0_DESTINATION_PE_BITMASK ;
    // PE33, Port1 next hop mask                 
    assign pe_inst[33].sys__pe__port1_destinationMask    = `NOC_CONT_PE33_PORT1_DESTINATION_PE_BITMASK ;
    // PE33, Port2 next hop mask                 
    assign pe_inst[33].sys__pe__port2_destinationMask    = `NOC_CONT_PE33_PORT2_DESTINATION_PE_BITMASK ;
    // PE33, Port3 next hop mask                 
    assign pe_inst[33].sys__pe__port3_destinationMask    = `NOC_CONT_PE33_PORT3_DESTINATION_PE_BITMASK ;
    // PE34, Port0 next hop mask                 
    assign pe_inst[34].sys__pe__port0_destinationMask    = `NOC_CONT_PE34_PORT0_DESTINATION_PE_BITMASK ;
    // PE34, Port1 next hop mask                 
    assign pe_inst[34].sys__pe__port1_destinationMask    = `NOC_CONT_PE34_PORT1_DESTINATION_PE_BITMASK ;
    // PE34, Port2 next hop mask                 
    assign pe_inst[34].sys__pe__port2_destinationMask    = `NOC_CONT_PE34_PORT2_DESTINATION_PE_BITMASK ;
    // PE34, Port3 next hop mask                 
    assign pe_inst[34].sys__pe__port3_destinationMask    = `NOC_CONT_PE34_PORT3_DESTINATION_PE_BITMASK ;
    // PE35, Port0 next hop mask                 
    assign pe_inst[35].sys__pe__port0_destinationMask    = `NOC_CONT_PE35_PORT0_DESTINATION_PE_BITMASK ;
    // PE35, Port1 next hop mask                 
    assign pe_inst[35].sys__pe__port1_destinationMask    = `NOC_CONT_PE35_PORT1_DESTINATION_PE_BITMASK ;
    // PE35, Port2 next hop mask                 
    assign pe_inst[35].sys__pe__port2_destinationMask    = `NOC_CONT_PE35_PORT2_DESTINATION_PE_BITMASK ;
    // PE35, Port3 next hop mask                 
    assign pe_inst[35].sys__pe__port3_destinationMask    = `NOC_CONT_PE35_PORT3_DESTINATION_PE_BITMASK ;
    // PE36, Port0 next hop mask                 
    assign pe_inst[36].sys__pe__port0_destinationMask    = `NOC_CONT_PE36_PORT0_DESTINATION_PE_BITMASK ;
    // PE36, Port1 next hop mask                 
    assign pe_inst[36].sys__pe__port1_destinationMask    = `NOC_CONT_PE36_PORT1_DESTINATION_PE_BITMASK ;
    // PE36, Port2 next hop mask                 
    assign pe_inst[36].sys__pe__port2_destinationMask    = `NOC_CONT_PE36_PORT2_DESTINATION_PE_BITMASK ;
    // PE36, Port3 next hop mask                 
    assign pe_inst[36].sys__pe__port3_destinationMask    = `NOC_CONT_PE36_PORT3_DESTINATION_PE_BITMASK ;
    // PE37, Port0 next hop mask                 
    assign pe_inst[37].sys__pe__port0_destinationMask    = `NOC_CONT_PE37_PORT0_DESTINATION_PE_BITMASK ;
    // PE37, Port1 next hop mask                 
    assign pe_inst[37].sys__pe__port1_destinationMask    = `NOC_CONT_PE37_PORT1_DESTINATION_PE_BITMASK ;
    // PE37, Port2 next hop mask                 
    assign pe_inst[37].sys__pe__port2_destinationMask    = `NOC_CONT_PE37_PORT2_DESTINATION_PE_BITMASK ;
    // PE37, Port3 next hop mask                 
    assign pe_inst[37].sys__pe__port3_destinationMask    = `NOC_CONT_PE37_PORT3_DESTINATION_PE_BITMASK ;
    // PE38, Port0 next hop mask                 
    assign pe_inst[38].sys__pe__port0_destinationMask    = `NOC_CONT_PE38_PORT0_DESTINATION_PE_BITMASK ;
    // PE38, Port1 next hop mask                 
    assign pe_inst[38].sys__pe__port1_destinationMask    = `NOC_CONT_PE38_PORT1_DESTINATION_PE_BITMASK ;
    // PE38, Port2 next hop mask                 
    assign pe_inst[38].sys__pe__port2_destinationMask    = `NOC_CONT_PE38_PORT2_DESTINATION_PE_BITMASK ;
    // PE38, Port3 next hop mask                 
    assign pe_inst[38].sys__pe__port3_destinationMask    = `NOC_CONT_PE38_PORT3_DESTINATION_PE_BITMASK ;
    // PE39, Port0 next hop mask                 
    assign pe_inst[39].sys__pe__port0_destinationMask    = `NOC_CONT_PE39_PORT0_DESTINATION_PE_BITMASK ;
    // PE39, Port1 next hop mask                 
    assign pe_inst[39].sys__pe__port1_destinationMask    = `NOC_CONT_PE39_PORT1_DESTINATION_PE_BITMASK ;
    // PE39, Port2 next hop mask                 
    assign pe_inst[39].sys__pe__port2_destinationMask    = `NOC_CONT_PE39_PORT2_DESTINATION_PE_BITMASK ;
    // PE39, Port3 next hop mask                 
    assign pe_inst[39].sys__pe__port3_destinationMask    = `NOC_CONT_PE39_PORT3_DESTINATION_PE_BITMASK ;
    // PE40, Port0 next hop mask                 
    assign pe_inst[40].sys__pe__port0_destinationMask    = `NOC_CONT_PE40_PORT0_DESTINATION_PE_BITMASK ;
    // PE40, Port1 next hop mask                 
    assign pe_inst[40].sys__pe__port1_destinationMask    = `NOC_CONT_PE40_PORT1_DESTINATION_PE_BITMASK ;
    // PE40, Port2 next hop mask                 
    assign pe_inst[40].sys__pe__port2_destinationMask    = `NOC_CONT_PE40_PORT2_DESTINATION_PE_BITMASK ;
    // PE40, Port3 next hop mask                 
    assign pe_inst[40].sys__pe__port3_destinationMask    = `NOC_CONT_PE40_PORT3_DESTINATION_PE_BITMASK ;
    // PE41, Port0 next hop mask                 
    assign pe_inst[41].sys__pe__port0_destinationMask    = `NOC_CONT_PE41_PORT0_DESTINATION_PE_BITMASK ;
    // PE41, Port1 next hop mask                 
    assign pe_inst[41].sys__pe__port1_destinationMask    = `NOC_CONT_PE41_PORT1_DESTINATION_PE_BITMASK ;
    // PE41, Port2 next hop mask                 
    assign pe_inst[41].sys__pe__port2_destinationMask    = `NOC_CONT_PE41_PORT2_DESTINATION_PE_BITMASK ;
    // PE41, Port3 next hop mask                 
    assign pe_inst[41].sys__pe__port3_destinationMask    = `NOC_CONT_PE41_PORT3_DESTINATION_PE_BITMASK ;
    // PE42, Port0 next hop mask                 
    assign pe_inst[42].sys__pe__port0_destinationMask    = `NOC_CONT_PE42_PORT0_DESTINATION_PE_BITMASK ;
    // PE42, Port1 next hop mask                 
    assign pe_inst[42].sys__pe__port1_destinationMask    = `NOC_CONT_PE42_PORT1_DESTINATION_PE_BITMASK ;
    // PE42, Port2 next hop mask                 
    assign pe_inst[42].sys__pe__port2_destinationMask    = `NOC_CONT_PE42_PORT2_DESTINATION_PE_BITMASK ;
    // PE42, Port3 next hop mask                 
    assign pe_inst[42].sys__pe__port3_destinationMask    = `NOC_CONT_PE42_PORT3_DESTINATION_PE_BITMASK ;
    // PE43, Port0 next hop mask                 
    assign pe_inst[43].sys__pe__port0_destinationMask    = `NOC_CONT_PE43_PORT0_DESTINATION_PE_BITMASK ;
    // PE43, Port1 next hop mask                 
    assign pe_inst[43].sys__pe__port1_destinationMask    = `NOC_CONT_PE43_PORT1_DESTINATION_PE_BITMASK ;
    // PE43, Port2 next hop mask                 
    assign pe_inst[43].sys__pe__port2_destinationMask    = `NOC_CONT_PE43_PORT2_DESTINATION_PE_BITMASK ;
    // PE43, Port3 next hop mask                 
    assign pe_inst[43].sys__pe__port3_destinationMask    = `NOC_CONT_PE43_PORT3_DESTINATION_PE_BITMASK ;
    // PE44, Port0 next hop mask                 
    assign pe_inst[44].sys__pe__port0_destinationMask    = `NOC_CONT_PE44_PORT0_DESTINATION_PE_BITMASK ;
    // PE44, Port1 next hop mask                 
    assign pe_inst[44].sys__pe__port1_destinationMask    = `NOC_CONT_PE44_PORT1_DESTINATION_PE_BITMASK ;
    // PE44, Port2 next hop mask                 
    assign pe_inst[44].sys__pe__port2_destinationMask    = `NOC_CONT_PE44_PORT2_DESTINATION_PE_BITMASK ;
    // PE44, Port3 next hop mask                 
    assign pe_inst[44].sys__pe__port3_destinationMask    = `NOC_CONT_PE44_PORT3_DESTINATION_PE_BITMASK ;
    // PE45, Port0 next hop mask                 
    assign pe_inst[45].sys__pe__port0_destinationMask    = `NOC_CONT_PE45_PORT0_DESTINATION_PE_BITMASK ;
    // PE45, Port1 next hop mask                 
    assign pe_inst[45].sys__pe__port1_destinationMask    = `NOC_CONT_PE45_PORT1_DESTINATION_PE_BITMASK ;
    // PE45, Port2 next hop mask                 
    assign pe_inst[45].sys__pe__port2_destinationMask    = `NOC_CONT_PE45_PORT2_DESTINATION_PE_BITMASK ;
    // PE45, Port3 next hop mask                 
    assign pe_inst[45].sys__pe__port3_destinationMask    = `NOC_CONT_PE45_PORT3_DESTINATION_PE_BITMASK ;
    // PE46, Port0 next hop mask                 
    assign pe_inst[46].sys__pe__port0_destinationMask    = `NOC_CONT_PE46_PORT0_DESTINATION_PE_BITMASK ;
    // PE46, Port1 next hop mask                 
    assign pe_inst[46].sys__pe__port1_destinationMask    = `NOC_CONT_PE46_PORT1_DESTINATION_PE_BITMASK ;
    // PE46, Port2 next hop mask                 
    assign pe_inst[46].sys__pe__port2_destinationMask    = `NOC_CONT_PE46_PORT2_DESTINATION_PE_BITMASK ;
    // PE46, Port3 next hop mask                 
    assign pe_inst[46].sys__pe__port3_destinationMask    = `NOC_CONT_PE46_PORT3_DESTINATION_PE_BITMASK ;
    // PE47, Port0 next hop mask                 
    assign pe_inst[47].sys__pe__port0_destinationMask    = `NOC_CONT_PE47_PORT0_DESTINATION_PE_BITMASK ;
    // PE47, Port1 next hop mask                 
    assign pe_inst[47].sys__pe__port1_destinationMask    = `NOC_CONT_PE47_PORT1_DESTINATION_PE_BITMASK ;
    // PE47, Port2 next hop mask                 
    assign pe_inst[47].sys__pe__port2_destinationMask    = `NOC_CONT_PE47_PORT2_DESTINATION_PE_BITMASK ;
    // PE47, Port3 next hop mask                 
    assign pe_inst[47].sys__pe__port3_destinationMask    = `NOC_CONT_PE47_PORT3_DESTINATION_PE_BITMASK ;
    // PE48, Port0 next hop mask                 
    assign pe_inst[48].sys__pe__port0_destinationMask    = `NOC_CONT_PE48_PORT0_DESTINATION_PE_BITMASK ;
    // PE48, Port1 next hop mask                 
    assign pe_inst[48].sys__pe__port1_destinationMask    = `NOC_CONT_PE48_PORT1_DESTINATION_PE_BITMASK ;
    // PE48, Port2 next hop mask                 
    assign pe_inst[48].sys__pe__port2_destinationMask    = `NOC_CONT_PE48_PORT2_DESTINATION_PE_BITMASK ;
    // PE48, Port3 next hop mask                 
    assign pe_inst[48].sys__pe__port3_destinationMask    = `NOC_CONT_PE48_PORT3_DESTINATION_PE_BITMASK ;
    // PE49, Port0 next hop mask                 
    assign pe_inst[49].sys__pe__port0_destinationMask    = `NOC_CONT_PE49_PORT0_DESTINATION_PE_BITMASK ;
    // PE49, Port1 next hop mask                 
    assign pe_inst[49].sys__pe__port1_destinationMask    = `NOC_CONT_PE49_PORT1_DESTINATION_PE_BITMASK ;
    // PE49, Port2 next hop mask                 
    assign pe_inst[49].sys__pe__port2_destinationMask    = `NOC_CONT_PE49_PORT2_DESTINATION_PE_BITMASK ;
    // PE49, Port3 next hop mask                 
    assign pe_inst[49].sys__pe__port3_destinationMask    = `NOC_CONT_PE49_PORT3_DESTINATION_PE_BITMASK ;
    // PE50, Port0 next hop mask                 
    assign pe_inst[50].sys__pe__port0_destinationMask    = `NOC_CONT_PE50_PORT0_DESTINATION_PE_BITMASK ;
    // PE50, Port1 next hop mask                 
    assign pe_inst[50].sys__pe__port1_destinationMask    = `NOC_CONT_PE50_PORT1_DESTINATION_PE_BITMASK ;
    // PE50, Port2 next hop mask                 
    assign pe_inst[50].sys__pe__port2_destinationMask    = `NOC_CONT_PE50_PORT2_DESTINATION_PE_BITMASK ;
    // PE50, Port3 next hop mask                 
    assign pe_inst[50].sys__pe__port3_destinationMask    = `NOC_CONT_PE50_PORT3_DESTINATION_PE_BITMASK ;
    // PE51, Port0 next hop mask                 
    assign pe_inst[51].sys__pe__port0_destinationMask    = `NOC_CONT_PE51_PORT0_DESTINATION_PE_BITMASK ;
    // PE51, Port1 next hop mask                 
    assign pe_inst[51].sys__pe__port1_destinationMask    = `NOC_CONT_PE51_PORT1_DESTINATION_PE_BITMASK ;
    // PE51, Port2 next hop mask                 
    assign pe_inst[51].sys__pe__port2_destinationMask    = `NOC_CONT_PE51_PORT2_DESTINATION_PE_BITMASK ;
    // PE51, Port3 next hop mask                 
    assign pe_inst[51].sys__pe__port3_destinationMask    = `NOC_CONT_PE51_PORT3_DESTINATION_PE_BITMASK ;
    // PE52, Port0 next hop mask                 
    assign pe_inst[52].sys__pe__port0_destinationMask    = `NOC_CONT_PE52_PORT0_DESTINATION_PE_BITMASK ;
    // PE52, Port1 next hop mask                 
    assign pe_inst[52].sys__pe__port1_destinationMask    = `NOC_CONT_PE52_PORT1_DESTINATION_PE_BITMASK ;
    // PE52, Port2 next hop mask                 
    assign pe_inst[52].sys__pe__port2_destinationMask    = `NOC_CONT_PE52_PORT2_DESTINATION_PE_BITMASK ;
    // PE52, Port3 next hop mask                 
    assign pe_inst[52].sys__pe__port3_destinationMask    = `NOC_CONT_PE52_PORT3_DESTINATION_PE_BITMASK ;
    // PE53, Port0 next hop mask                 
    assign pe_inst[53].sys__pe__port0_destinationMask    = `NOC_CONT_PE53_PORT0_DESTINATION_PE_BITMASK ;
    // PE53, Port1 next hop mask                 
    assign pe_inst[53].sys__pe__port1_destinationMask    = `NOC_CONT_PE53_PORT1_DESTINATION_PE_BITMASK ;
    // PE53, Port2 next hop mask                 
    assign pe_inst[53].sys__pe__port2_destinationMask    = `NOC_CONT_PE53_PORT2_DESTINATION_PE_BITMASK ;
    // PE53, Port3 next hop mask                 
    assign pe_inst[53].sys__pe__port3_destinationMask    = `NOC_CONT_PE53_PORT3_DESTINATION_PE_BITMASK ;
    // PE54, Port0 next hop mask                 
    assign pe_inst[54].sys__pe__port0_destinationMask    = `NOC_CONT_PE54_PORT0_DESTINATION_PE_BITMASK ;
    // PE54, Port1 next hop mask                 
    assign pe_inst[54].sys__pe__port1_destinationMask    = `NOC_CONT_PE54_PORT1_DESTINATION_PE_BITMASK ;
    // PE54, Port2 next hop mask                 
    assign pe_inst[54].sys__pe__port2_destinationMask    = `NOC_CONT_PE54_PORT2_DESTINATION_PE_BITMASK ;
    // PE54, Port3 next hop mask                 
    assign pe_inst[54].sys__pe__port3_destinationMask    = `NOC_CONT_PE54_PORT3_DESTINATION_PE_BITMASK ;
    // PE55, Port0 next hop mask                 
    assign pe_inst[55].sys__pe__port0_destinationMask    = `NOC_CONT_PE55_PORT0_DESTINATION_PE_BITMASK ;
    // PE55, Port1 next hop mask                 
    assign pe_inst[55].sys__pe__port1_destinationMask    = `NOC_CONT_PE55_PORT1_DESTINATION_PE_BITMASK ;
    // PE55, Port2 next hop mask                 
    assign pe_inst[55].sys__pe__port2_destinationMask    = `NOC_CONT_PE55_PORT2_DESTINATION_PE_BITMASK ;
    // PE55, Port3 next hop mask                 
    assign pe_inst[55].sys__pe__port3_destinationMask    = `NOC_CONT_PE55_PORT3_DESTINATION_PE_BITMASK ;
    // PE56, Port0 next hop mask                 
    assign pe_inst[56].sys__pe__port0_destinationMask    = `NOC_CONT_PE56_PORT0_DESTINATION_PE_BITMASK ;
    // PE56, Port1 next hop mask                 
    assign pe_inst[56].sys__pe__port1_destinationMask    = `NOC_CONT_PE56_PORT1_DESTINATION_PE_BITMASK ;
    // PE56, Port2 next hop mask                 
    assign pe_inst[56].sys__pe__port2_destinationMask    = `NOC_CONT_PE56_PORT2_DESTINATION_PE_BITMASK ;
    // PE56, Port3 next hop mask                 
    assign pe_inst[56].sys__pe__port3_destinationMask    = `NOC_CONT_PE56_PORT3_DESTINATION_PE_BITMASK ;
    // PE57, Port0 next hop mask                 
    assign pe_inst[57].sys__pe__port0_destinationMask    = `NOC_CONT_PE57_PORT0_DESTINATION_PE_BITMASK ;
    // PE57, Port1 next hop mask                 
    assign pe_inst[57].sys__pe__port1_destinationMask    = `NOC_CONT_PE57_PORT1_DESTINATION_PE_BITMASK ;
    // PE57, Port2 next hop mask                 
    assign pe_inst[57].sys__pe__port2_destinationMask    = `NOC_CONT_PE57_PORT2_DESTINATION_PE_BITMASK ;
    // PE57, Port3 next hop mask                 
    assign pe_inst[57].sys__pe__port3_destinationMask    = `NOC_CONT_PE57_PORT3_DESTINATION_PE_BITMASK ;
    // PE58, Port0 next hop mask                 
    assign pe_inst[58].sys__pe__port0_destinationMask    = `NOC_CONT_PE58_PORT0_DESTINATION_PE_BITMASK ;
    // PE58, Port1 next hop mask                 
    assign pe_inst[58].sys__pe__port1_destinationMask    = `NOC_CONT_PE58_PORT1_DESTINATION_PE_BITMASK ;
    // PE58, Port2 next hop mask                 
    assign pe_inst[58].sys__pe__port2_destinationMask    = `NOC_CONT_PE58_PORT2_DESTINATION_PE_BITMASK ;
    // PE58, Port3 next hop mask                 
    assign pe_inst[58].sys__pe__port3_destinationMask    = `NOC_CONT_PE58_PORT3_DESTINATION_PE_BITMASK ;
    // PE59, Port0 next hop mask                 
    assign pe_inst[59].sys__pe__port0_destinationMask    = `NOC_CONT_PE59_PORT0_DESTINATION_PE_BITMASK ;
    // PE59, Port1 next hop mask                 
    assign pe_inst[59].sys__pe__port1_destinationMask    = `NOC_CONT_PE59_PORT1_DESTINATION_PE_BITMASK ;
    // PE59, Port2 next hop mask                 
    assign pe_inst[59].sys__pe__port2_destinationMask    = `NOC_CONT_PE59_PORT2_DESTINATION_PE_BITMASK ;
    // PE59, Port3 next hop mask                 
    assign pe_inst[59].sys__pe__port3_destinationMask    = `NOC_CONT_PE59_PORT3_DESTINATION_PE_BITMASK ;
    // PE60, Port0 next hop mask                 
    assign pe_inst[60].sys__pe__port0_destinationMask    = `NOC_CONT_PE60_PORT0_DESTINATION_PE_BITMASK ;
    // PE60, Port1 next hop mask                 
    assign pe_inst[60].sys__pe__port1_destinationMask    = `NOC_CONT_PE60_PORT1_DESTINATION_PE_BITMASK ;
    // PE60, Port2 next hop mask                 
    assign pe_inst[60].sys__pe__port2_destinationMask    = `NOC_CONT_PE60_PORT2_DESTINATION_PE_BITMASK ;
    // PE60, Port3 next hop mask                 
    assign pe_inst[60].sys__pe__port3_destinationMask    = `NOC_CONT_PE60_PORT3_DESTINATION_PE_BITMASK ;
    // PE61, Port0 next hop mask                 
    assign pe_inst[61].sys__pe__port0_destinationMask    = `NOC_CONT_PE61_PORT0_DESTINATION_PE_BITMASK ;
    // PE61, Port1 next hop mask                 
    assign pe_inst[61].sys__pe__port1_destinationMask    = `NOC_CONT_PE61_PORT1_DESTINATION_PE_BITMASK ;
    // PE61, Port2 next hop mask                 
    assign pe_inst[61].sys__pe__port2_destinationMask    = `NOC_CONT_PE61_PORT2_DESTINATION_PE_BITMASK ;
    // PE61, Port3 next hop mask                 
    assign pe_inst[61].sys__pe__port3_destinationMask    = `NOC_CONT_PE61_PORT3_DESTINATION_PE_BITMASK ;
    // PE62, Port0 next hop mask                 
    assign pe_inst[62].sys__pe__port0_destinationMask    = `NOC_CONT_PE62_PORT0_DESTINATION_PE_BITMASK ;
    // PE62, Port1 next hop mask                 
    assign pe_inst[62].sys__pe__port1_destinationMask    = `NOC_CONT_PE62_PORT1_DESTINATION_PE_BITMASK ;
    // PE62, Port2 next hop mask                 
    assign pe_inst[62].sys__pe__port2_destinationMask    = `NOC_CONT_PE62_PORT2_DESTINATION_PE_BITMASK ;
    // PE62, Port3 next hop mask                 
    assign pe_inst[62].sys__pe__port3_destinationMask    = `NOC_CONT_PE62_PORT3_DESTINATION_PE_BITMASK ;
    // PE63, Port0 next hop mask                 
    assign pe_inst[63].sys__pe__port0_destinationMask    = `NOC_CONT_PE63_PORT0_DESTINATION_PE_BITMASK ;
    // PE63, Port1 next hop mask                 
    assign pe_inst[63].sys__pe__port1_destinationMask    = `NOC_CONT_PE63_PORT1_DESTINATION_PE_BITMASK ;
    // PE63, Port2 next hop mask                 
    assign pe_inst[63].sys__pe__port2_destinationMask    = `NOC_CONT_PE63_PORT2_DESTINATION_PE_BITMASK ;
    // PE63, Port3 next hop mask                 
    assign pe_inst[63].sys__pe__port3_destinationMask    = `NOC_CONT_PE63_PORT3_DESTINATION_PE_BITMASK ;