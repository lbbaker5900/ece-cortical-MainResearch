
    output                                         pe0__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe0__stu__cntl           ;
    input                                          stu__pe0__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe0__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe0__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe0__stu__oob_data       ;

    output                                         pe1__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe1__stu__cntl           ;
    input                                          stu__pe1__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe1__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe1__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe1__stu__oob_data       ;

    output                                         pe2__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe2__stu__cntl           ;
    input                                          stu__pe2__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe2__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe2__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe2__stu__oob_data       ;

    output                                         pe3__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe3__stu__cntl           ;
    input                                          stu__pe3__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe3__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe3__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe3__stu__oob_data       ;

    output                                         pe4__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe4__stu__cntl           ;
    input                                          stu__pe4__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe4__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe4__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe4__stu__oob_data       ;

    output                                         pe5__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe5__stu__cntl           ;
    input                                          stu__pe5__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe5__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe5__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe5__stu__oob_data       ;

    output                                         pe6__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe6__stu__cntl           ;
    input                                          stu__pe6__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe6__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe6__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe6__stu__oob_data       ;

    output                                         pe7__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe7__stu__cntl           ;
    input                                          stu__pe7__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe7__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe7__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe7__stu__oob_data       ;

    output                                         pe8__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe8__stu__cntl           ;
    input                                          stu__pe8__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe8__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe8__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe8__stu__oob_data       ;

    output                                         pe9__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe9__stu__cntl           ;
    input                                          stu__pe9__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe9__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe9__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe9__stu__oob_data       ;

    output                                         pe10__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe10__stu__cntl           ;
    input                                          stu__pe10__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe10__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe10__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe10__stu__oob_data       ;

    output                                         pe11__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe11__stu__cntl           ;
    input                                          stu__pe11__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe11__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe11__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe11__stu__oob_data       ;

    output                                         pe12__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe12__stu__cntl           ;
    input                                          stu__pe12__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe12__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe12__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe12__stu__oob_data       ;

    output                                         pe13__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe13__stu__cntl           ;
    input                                          stu__pe13__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe13__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe13__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe13__stu__oob_data       ;

    output                                         pe14__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe14__stu__cntl           ;
    input                                          stu__pe14__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe14__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe14__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe14__stu__oob_data       ;

    output                                         pe15__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe15__stu__cntl           ;
    input                                          stu__pe15__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe15__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe15__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe15__stu__oob_data       ;

    output                                         pe16__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe16__stu__cntl           ;
    input                                          stu__pe16__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe16__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe16__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe16__stu__oob_data       ;

    output                                         pe17__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe17__stu__cntl           ;
    input                                          stu__pe17__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe17__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe17__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe17__stu__oob_data       ;

    output                                         pe18__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe18__stu__cntl           ;
    input                                          stu__pe18__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe18__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe18__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe18__stu__oob_data       ;

    output                                         pe19__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe19__stu__cntl           ;
    input                                          stu__pe19__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe19__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe19__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe19__stu__oob_data       ;

    output                                         pe20__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe20__stu__cntl           ;
    input                                          stu__pe20__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe20__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe20__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe20__stu__oob_data       ;

    output                                         pe21__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe21__stu__cntl           ;
    input                                          stu__pe21__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe21__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe21__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe21__stu__oob_data       ;

    output                                         pe22__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe22__stu__cntl           ;
    input                                          stu__pe22__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe22__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe22__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe22__stu__oob_data       ;

    output                                         pe23__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe23__stu__cntl           ;
    input                                          stu__pe23__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe23__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe23__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe23__stu__oob_data       ;

    output                                         pe24__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe24__stu__cntl           ;
    input                                          stu__pe24__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe24__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe24__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe24__stu__oob_data       ;

    output                                         pe25__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe25__stu__cntl           ;
    input                                          stu__pe25__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe25__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe25__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe25__stu__oob_data       ;

    output                                         pe26__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe26__stu__cntl           ;
    input                                          stu__pe26__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe26__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe26__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe26__stu__oob_data       ;

    output                                         pe27__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe27__stu__cntl           ;
    input                                          stu__pe27__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe27__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe27__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe27__stu__oob_data       ;

    output                                         pe28__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe28__stu__cntl           ;
    input                                          stu__pe28__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe28__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe28__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe28__stu__oob_data       ;

    output                                         pe29__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe29__stu__cntl           ;
    input                                          stu__pe29__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe29__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe29__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe29__stu__oob_data       ;

    output                                         pe30__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe30__stu__cntl           ;
    input                                          stu__pe30__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe30__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe30__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe30__stu__oob_data       ;

    output                                         pe31__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe31__stu__cntl           ;
    input                                          stu__pe31__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe31__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe31__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe31__stu__oob_data       ;

    output                                         pe32__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe32__stu__cntl           ;
    input                                          stu__pe32__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe32__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe32__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe32__stu__oob_data       ;

    output                                         pe33__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe33__stu__cntl           ;
    input                                          stu__pe33__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe33__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe33__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe33__stu__oob_data       ;

    output                                         pe34__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe34__stu__cntl           ;
    input                                          stu__pe34__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe34__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe34__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe34__stu__oob_data       ;

    output                                         pe35__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe35__stu__cntl           ;
    input                                          stu__pe35__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe35__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe35__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe35__stu__oob_data       ;

    output                                         pe36__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe36__stu__cntl           ;
    input                                          stu__pe36__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe36__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe36__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe36__stu__oob_data       ;

    output                                         pe37__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe37__stu__cntl           ;
    input                                          stu__pe37__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe37__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe37__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe37__stu__oob_data       ;

    output                                         pe38__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe38__stu__cntl           ;
    input                                          stu__pe38__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe38__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe38__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe38__stu__oob_data       ;

    output                                         pe39__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe39__stu__cntl           ;
    input                                          stu__pe39__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe39__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe39__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe39__stu__oob_data       ;

    output                                         pe40__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe40__stu__cntl           ;
    input                                          stu__pe40__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe40__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe40__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe40__stu__oob_data       ;

    output                                         pe41__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe41__stu__cntl           ;
    input                                          stu__pe41__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe41__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe41__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe41__stu__oob_data       ;

    output                                         pe42__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe42__stu__cntl           ;
    input                                          stu__pe42__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe42__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe42__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe42__stu__oob_data       ;

    output                                         pe43__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe43__stu__cntl           ;
    input                                          stu__pe43__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe43__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe43__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe43__stu__oob_data       ;

    output                                         pe44__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe44__stu__cntl           ;
    input                                          stu__pe44__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe44__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe44__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe44__stu__oob_data       ;

    output                                         pe45__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe45__stu__cntl           ;
    input                                          stu__pe45__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe45__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe45__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe45__stu__oob_data       ;

    output                                         pe46__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe46__stu__cntl           ;
    input                                          stu__pe46__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe46__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe46__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe46__stu__oob_data       ;

    output                                         pe47__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe47__stu__cntl           ;
    input                                          stu__pe47__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe47__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe47__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe47__stu__oob_data       ;

    output                                         pe48__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe48__stu__cntl           ;
    input                                          stu__pe48__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe48__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe48__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe48__stu__oob_data       ;

    output                                         pe49__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe49__stu__cntl           ;
    input                                          stu__pe49__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe49__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe49__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe49__stu__oob_data       ;

    output                                         pe50__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe50__stu__cntl           ;
    input                                          stu__pe50__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe50__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe50__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe50__stu__oob_data       ;

    output                                         pe51__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe51__stu__cntl           ;
    input                                          stu__pe51__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe51__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe51__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe51__stu__oob_data       ;

    output                                         pe52__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe52__stu__cntl           ;
    input                                          stu__pe52__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe52__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe52__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe52__stu__oob_data       ;

    output                                         pe53__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe53__stu__cntl           ;
    input                                          stu__pe53__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe53__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe53__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe53__stu__oob_data       ;

    output                                         pe54__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe54__stu__cntl           ;
    input                                          stu__pe54__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe54__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe54__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe54__stu__oob_data       ;

    output                                         pe55__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe55__stu__cntl           ;
    input                                          stu__pe55__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe55__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe55__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe55__stu__oob_data       ;

    output                                         pe56__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe56__stu__cntl           ;
    input                                          stu__pe56__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe56__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe56__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe56__stu__oob_data       ;

    output                                         pe57__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe57__stu__cntl           ;
    input                                          stu__pe57__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe57__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe57__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe57__stu__oob_data       ;

    output                                         pe58__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe58__stu__cntl           ;
    input                                          stu__pe58__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe58__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe58__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe58__stu__oob_data       ;

    output                                         pe59__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe59__stu__cntl           ;
    input                                          stu__pe59__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe59__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe59__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe59__stu__oob_data       ;

    output                                         pe60__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe60__stu__cntl           ;
    input                                          stu__pe60__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe60__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe60__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe60__stu__oob_data       ;

    output                                         pe61__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe61__stu__cntl           ;
    input                                          stu__pe61__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe61__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe61__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe61__stu__oob_data       ;

    output                                         pe62__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe62__stu__cntl           ;
    input                                          stu__pe62__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe62__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe62__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe62__stu__oob_data       ;

    output                                         pe63__stu__valid          ;
    output  [`COMMON_STD_INTF_CNTL_RANGE   ]       pe63__stu__cntl           ;
    input                                          stu__pe63__ready          ;
    output  [`STACK_UP_INTF_TYPE_RANGE     ]       pe63__stu__type           ;
    output  [`STACK_UP_INTF_DATA_RANGE     ]       pe63__stu__data           ;
    output  [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe63__stu__oob_data       ;

