
  // NoC port 0
  wire                                     mgr__noc__port0_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  mgr__noc__port0_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port0_data  ;
  wire                                     noc__mgr__port0_fc    ;
  wire                                     noc__mgr__port0_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  noc__mgr__port0_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port0_data  ;
  wire                                     mgr__noc__port0_fc    ;

  // NoC port 1
  wire                                     mgr__noc__port1_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  mgr__noc__port1_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port1_data  ;
  wire                                     noc__mgr__port1_fc    ;
  wire                                     noc__mgr__port1_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  noc__mgr__port1_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port1_data  ;
  wire                                     mgr__noc__port1_fc    ;

  // NoC port 2
  wire                                     mgr__noc__port2_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  mgr__noc__port2_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port2_data  ;
  wire                                     noc__mgr__port2_fc    ;
  wire                                     noc__mgr__port2_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  noc__mgr__port2_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port2_data  ;
  wire                                     mgr__noc__port2_fc    ;

  // NoC port 3
  wire                                     mgr__noc__port3_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  mgr__noc__port3_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  mgr__noc__port3_data  ;
  wire                                     noc__mgr__port3_fc    ;
  wire                                     noc__mgr__port3_valid ;
  wire   [`NOC_CONT_NOC_PORT_CNTL_RANGE ]  noc__mgr__port3_cntl  ;
  wire   [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__mgr__port3_data  ;
  wire                                     mgr__noc__port3_fc    ;

