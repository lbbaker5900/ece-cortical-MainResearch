
  // General control and status                                                 
  wire                                        mgr0__sys__allSynchronized     ;
  wire                                        sys__mgr0__thisSynchronized    ;
  wire                                        sys__mgr0__ready               ;
  wire                                        sys__mgr0__complete            ;

  // General control and status                                                 
  wire                                        mgr1__sys__allSynchronized     ;
  wire                                        sys__mgr1__thisSynchronized    ;
  wire                                        sys__mgr1__ready               ;
  wire                                        sys__mgr1__complete            ;

  // General control and status                                                 
  wire                                        mgr2__sys__allSynchronized     ;
  wire                                        sys__mgr2__thisSynchronized    ;
  wire                                        sys__mgr2__ready               ;
  wire                                        sys__mgr2__complete            ;

  // General control and status                                                 
  wire                                        mgr3__sys__allSynchronized     ;
  wire                                        sys__mgr3__thisSynchronized    ;
  wire                                        sys__mgr3__ready               ;
  wire                                        sys__mgr3__complete            ;

  // General control and status                                                 
  wire                                        mgr4__sys__allSynchronized     ;
  wire                                        sys__mgr4__thisSynchronized    ;
  wire                                        sys__mgr4__ready               ;
  wire                                        sys__mgr4__complete            ;

  // General control and status                                                 
  wire                                        mgr5__sys__allSynchronized     ;
  wire                                        sys__mgr5__thisSynchronized    ;
  wire                                        sys__mgr5__ready               ;
  wire                                        sys__mgr5__complete            ;

  // General control and status                                                 
  wire                                        mgr6__sys__allSynchronized     ;
  wire                                        sys__mgr6__thisSynchronized    ;
  wire                                        sys__mgr6__ready               ;
  wire                                        sys__mgr6__complete            ;

  // General control and status                                                 
  wire                                        mgr7__sys__allSynchronized     ;
  wire                                        sys__mgr7__thisSynchronized    ;
  wire                                        sys__mgr7__ready               ;
  wire                                        sys__mgr7__complete            ;

  // General control and status                                                 
  wire                                        mgr8__sys__allSynchronized     ;
  wire                                        sys__mgr8__thisSynchronized    ;
  wire                                        sys__mgr8__ready               ;
  wire                                        sys__mgr8__complete            ;

  // General control and status                                                 
  wire                                        mgr9__sys__allSynchronized     ;
  wire                                        sys__mgr9__thisSynchronized    ;
  wire                                        sys__mgr9__ready               ;
  wire                                        sys__mgr9__complete            ;

  // General control and status                                                 
  wire                                        mgr10__sys__allSynchronized     ;
  wire                                        sys__mgr10__thisSynchronized    ;
  wire                                        sys__mgr10__ready               ;
  wire                                        sys__mgr10__complete            ;

  // General control and status                                                 
  wire                                        mgr11__sys__allSynchronized     ;
  wire                                        sys__mgr11__thisSynchronized    ;
  wire                                        sys__mgr11__ready               ;
  wire                                        sys__mgr11__complete            ;

  // General control and status                                                 
  wire                                        mgr12__sys__allSynchronized     ;
  wire                                        sys__mgr12__thisSynchronized    ;
  wire                                        sys__mgr12__ready               ;
  wire                                        sys__mgr12__complete            ;

  // General control and status                                                 
  wire                                        mgr13__sys__allSynchronized     ;
  wire                                        sys__mgr13__thisSynchronized    ;
  wire                                        sys__mgr13__ready               ;
  wire                                        sys__mgr13__complete            ;

  // General control and status                                                 
  wire                                        mgr14__sys__allSynchronized     ;
  wire                                        sys__mgr14__thisSynchronized    ;
  wire                                        sys__mgr14__ready               ;
  wire                                        sys__mgr14__complete            ;

  // General control and status                                                 
  wire                                        mgr15__sys__allSynchronized     ;
  wire                                        sys__mgr15__thisSynchronized    ;
  wire                                        sys__mgr15__ready               ;
  wire                                        sys__mgr15__complete            ;

  // General control and status                                                 
  wire                                        mgr16__sys__allSynchronized     ;
  wire                                        sys__mgr16__thisSynchronized    ;
  wire                                        sys__mgr16__ready               ;
  wire                                        sys__mgr16__complete            ;

  // General control and status                                                 
  wire                                        mgr17__sys__allSynchronized     ;
  wire                                        sys__mgr17__thisSynchronized    ;
  wire                                        sys__mgr17__ready               ;
  wire                                        sys__mgr17__complete            ;

  // General control and status                                                 
  wire                                        mgr18__sys__allSynchronized     ;
  wire                                        sys__mgr18__thisSynchronized    ;
  wire                                        sys__mgr18__ready               ;
  wire                                        sys__mgr18__complete            ;

  // General control and status                                                 
  wire                                        mgr19__sys__allSynchronized     ;
  wire                                        sys__mgr19__thisSynchronized    ;
  wire                                        sys__mgr19__ready               ;
  wire                                        sys__mgr19__complete            ;

  // General control and status                                                 
  wire                                        mgr20__sys__allSynchronized     ;
  wire                                        sys__mgr20__thisSynchronized    ;
  wire                                        sys__mgr20__ready               ;
  wire                                        sys__mgr20__complete            ;

  // General control and status                                                 
  wire                                        mgr21__sys__allSynchronized     ;
  wire                                        sys__mgr21__thisSynchronized    ;
  wire                                        sys__mgr21__ready               ;
  wire                                        sys__mgr21__complete            ;

  // General control and status                                                 
  wire                                        mgr22__sys__allSynchronized     ;
  wire                                        sys__mgr22__thisSynchronized    ;
  wire                                        sys__mgr22__ready               ;
  wire                                        sys__mgr22__complete            ;

  // General control and status                                                 
  wire                                        mgr23__sys__allSynchronized     ;
  wire                                        sys__mgr23__thisSynchronized    ;
  wire                                        sys__mgr23__ready               ;
  wire                                        sys__mgr23__complete            ;

  // General control and status                                                 
  wire                                        mgr24__sys__allSynchronized     ;
  wire                                        sys__mgr24__thisSynchronized    ;
  wire                                        sys__mgr24__ready               ;
  wire                                        sys__mgr24__complete            ;

  // General control and status                                                 
  wire                                        mgr25__sys__allSynchronized     ;
  wire                                        sys__mgr25__thisSynchronized    ;
  wire                                        sys__mgr25__ready               ;
  wire                                        sys__mgr25__complete            ;

  // General control and status                                                 
  wire                                        mgr26__sys__allSynchronized     ;
  wire                                        sys__mgr26__thisSynchronized    ;
  wire                                        sys__mgr26__ready               ;
  wire                                        sys__mgr26__complete            ;

  // General control and status                                                 
  wire                                        mgr27__sys__allSynchronized     ;
  wire                                        sys__mgr27__thisSynchronized    ;
  wire                                        sys__mgr27__ready               ;
  wire                                        sys__mgr27__complete            ;

  // General control and status                                                 
  wire                                        mgr28__sys__allSynchronized     ;
  wire                                        sys__mgr28__thisSynchronized    ;
  wire                                        sys__mgr28__ready               ;
  wire                                        sys__mgr28__complete            ;

  // General control and status                                                 
  wire                                        mgr29__sys__allSynchronized     ;
  wire                                        sys__mgr29__thisSynchronized    ;
  wire                                        sys__mgr29__ready               ;
  wire                                        sys__mgr29__complete            ;

  // General control and status                                                 
  wire                                        mgr30__sys__allSynchronized     ;
  wire                                        sys__mgr30__thisSynchronized    ;
  wire                                        sys__mgr30__ready               ;
  wire                                        sys__mgr30__complete            ;

  // General control and status                                                 
  wire                                        mgr31__sys__allSynchronized     ;
  wire                                        sys__mgr31__thisSynchronized    ;
  wire                                        sys__mgr31__ready               ;
  wire                                        sys__mgr31__complete            ;

  // General control and status                                                 
  wire                                        mgr32__sys__allSynchronized     ;
  wire                                        sys__mgr32__thisSynchronized    ;
  wire                                        sys__mgr32__ready               ;
  wire                                        sys__mgr32__complete            ;

  // General control and status                                                 
  wire                                        mgr33__sys__allSynchronized     ;
  wire                                        sys__mgr33__thisSynchronized    ;
  wire                                        sys__mgr33__ready               ;
  wire                                        sys__mgr33__complete            ;

  // General control and status                                                 
  wire                                        mgr34__sys__allSynchronized     ;
  wire                                        sys__mgr34__thisSynchronized    ;
  wire                                        sys__mgr34__ready               ;
  wire                                        sys__mgr34__complete            ;

  // General control and status                                                 
  wire                                        mgr35__sys__allSynchronized     ;
  wire                                        sys__mgr35__thisSynchronized    ;
  wire                                        sys__mgr35__ready               ;
  wire                                        sys__mgr35__complete            ;

  // General control and status                                                 
  wire                                        mgr36__sys__allSynchronized     ;
  wire                                        sys__mgr36__thisSynchronized    ;
  wire                                        sys__mgr36__ready               ;
  wire                                        sys__mgr36__complete            ;

  // General control and status                                                 
  wire                                        mgr37__sys__allSynchronized     ;
  wire                                        sys__mgr37__thisSynchronized    ;
  wire                                        sys__mgr37__ready               ;
  wire                                        sys__mgr37__complete            ;

  // General control and status                                                 
  wire                                        mgr38__sys__allSynchronized     ;
  wire                                        sys__mgr38__thisSynchronized    ;
  wire                                        sys__mgr38__ready               ;
  wire                                        sys__mgr38__complete            ;

  // General control and status                                                 
  wire                                        mgr39__sys__allSynchronized     ;
  wire                                        sys__mgr39__thisSynchronized    ;
  wire                                        sys__mgr39__ready               ;
  wire                                        sys__mgr39__complete            ;

  // General control and status                                                 
  wire                                        mgr40__sys__allSynchronized     ;
  wire                                        sys__mgr40__thisSynchronized    ;
  wire                                        sys__mgr40__ready               ;
  wire                                        sys__mgr40__complete            ;

  // General control and status                                                 
  wire                                        mgr41__sys__allSynchronized     ;
  wire                                        sys__mgr41__thisSynchronized    ;
  wire                                        sys__mgr41__ready               ;
  wire                                        sys__mgr41__complete            ;

  // General control and status                                                 
  wire                                        mgr42__sys__allSynchronized     ;
  wire                                        sys__mgr42__thisSynchronized    ;
  wire                                        sys__mgr42__ready               ;
  wire                                        sys__mgr42__complete            ;

  // General control and status                                                 
  wire                                        mgr43__sys__allSynchronized     ;
  wire                                        sys__mgr43__thisSynchronized    ;
  wire                                        sys__mgr43__ready               ;
  wire                                        sys__mgr43__complete            ;

  // General control and status                                                 
  wire                                        mgr44__sys__allSynchronized     ;
  wire                                        sys__mgr44__thisSynchronized    ;
  wire                                        sys__mgr44__ready               ;
  wire                                        sys__mgr44__complete            ;

  // General control and status                                                 
  wire                                        mgr45__sys__allSynchronized     ;
  wire                                        sys__mgr45__thisSynchronized    ;
  wire                                        sys__mgr45__ready               ;
  wire                                        sys__mgr45__complete            ;

  // General control and status                                                 
  wire                                        mgr46__sys__allSynchronized     ;
  wire                                        sys__mgr46__thisSynchronized    ;
  wire                                        sys__mgr46__ready               ;
  wire                                        sys__mgr46__complete            ;

  // General control and status                                                 
  wire                                        mgr47__sys__allSynchronized     ;
  wire                                        sys__mgr47__thisSynchronized    ;
  wire                                        sys__mgr47__ready               ;
  wire                                        sys__mgr47__complete            ;

  // General control and status                                                 
  wire                                        mgr48__sys__allSynchronized     ;
  wire                                        sys__mgr48__thisSynchronized    ;
  wire                                        sys__mgr48__ready               ;
  wire                                        sys__mgr48__complete            ;

  // General control and status                                                 
  wire                                        mgr49__sys__allSynchronized     ;
  wire                                        sys__mgr49__thisSynchronized    ;
  wire                                        sys__mgr49__ready               ;
  wire                                        sys__mgr49__complete            ;

  // General control and status                                                 
  wire                                        mgr50__sys__allSynchronized     ;
  wire                                        sys__mgr50__thisSynchronized    ;
  wire                                        sys__mgr50__ready               ;
  wire                                        sys__mgr50__complete            ;

  // General control and status                                                 
  wire                                        mgr51__sys__allSynchronized     ;
  wire                                        sys__mgr51__thisSynchronized    ;
  wire                                        sys__mgr51__ready               ;
  wire                                        sys__mgr51__complete            ;

  // General control and status                                                 
  wire                                        mgr52__sys__allSynchronized     ;
  wire                                        sys__mgr52__thisSynchronized    ;
  wire                                        sys__mgr52__ready               ;
  wire                                        sys__mgr52__complete            ;

  // General control and status                                                 
  wire                                        mgr53__sys__allSynchronized     ;
  wire                                        sys__mgr53__thisSynchronized    ;
  wire                                        sys__mgr53__ready               ;
  wire                                        sys__mgr53__complete            ;

  // General control and status                                                 
  wire                                        mgr54__sys__allSynchronized     ;
  wire                                        sys__mgr54__thisSynchronized    ;
  wire                                        sys__mgr54__ready               ;
  wire                                        sys__mgr54__complete            ;

  // General control and status                                                 
  wire                                        mgr55__sys__allSynchronized     ;
  wire                                        sys__mgr55__thisSynchronized    ;
  wire                                        sys__mgr55__ready               ;
  wire                                        sys__mgr55__complete            ;

  // General control and status                                                 
  wire                                        mgr56__sys__allSynchronized     ;
  wire                                        sys__mgr56__thisSynchronized    ;
  wire                                        sys__mgr56__ready               ;
  wire                                        sys__mgr56__complete            ;

  // General control and status                                                 
  wire                                        mgr57__sys__allSynchronized     ;
  wire                                        sys__mgr57__thisSynchronized    ;
  wire                                        sys__mgr57__ready               ;
  wire                                        sys__mgr57__complete            ;

  // General control and status                                                 
  wire                                        mgr58__sys__allSynchronized     ;
  wire                                        sys__mgr58__thisSynchronized    ;
  wire                                        sys__mgr58__ready               ;
  wire                                        sys__mgr58__complete            ;

  // General control and status                                                 
  wire                                        mgr59__sys__allSynchronized     ;
  wire                                        sys__mgr59__thisSynchronized    ;
  wire                                        sys__mgr59__ready               ;
  wire                                        sys__mgr59__complete            ;

  // General control and status                                                 
  wire                                        mgr60__sys__allSynchronized     ;
  wire                                        sys__mgr60__thisSynchronized    ;
  wire                                        sys__mgr60__ready               ;
  wire                                        sys__mgr60__complete            ;

  // General control and status                                                 
  wire                                        mgr61__sys__allSynchronized     ;
  wire                                        sys__mgr61__thisSynchronized    ;
  wire                                        sys__mgr61__ready               ;
  wire                                        sys__mgr61__complete            ;

  // General control and status                                                 
  wire                                        mgr62__sys__allSynchronized     ;
  wire                                        sys__mgr62__thisSynchronized    ;
  wire                                        sys__mgr62__ready               ;
  wire                                        sys__mgr62__complete            ;

  // General control and status                                                 
  wire                                        mgr63__sys__allSynchronized     ;
  wire                                        sys__mgr63__thisSynchronized    ;
  wire                                        sys__mgr63__ready               ;
  wire                                        sys__mgr63__complete            ;
