
 assign    stu__mgr0__valid       =    pe0__stu__valid          ;
 assign    stu__mgr0__cntl        =    pe0__stu__cntl           ;
 assign    stu__pe0__ready        =    mgr0__stu__ready         ;
 assign    stu__mgr0__type        =    pe0__stu__type           ;
 assign    stu__mgr0__data        =    pe0__stu__data           ;
 assign    stu__mgr0__oob_data    =    pe0__stu__oob_data       ;

 assign    stu__mgr1__valid       =    pe1__stu__valid          ;
 assign    stu__mgr1__cntl        =    pe1__stu__cntl           ;
 assign    stu__pe1__ready        =    mgr1__stu__ready         ;
 assign    stu__mgr1__type        =    pe1__stu__type           ;
 assign    stu__mgr1__data        =    pe1__stu__data           ;
 assign    stu__mgr1__oob_data    =    pe1__stu__oob_data       ;

 assign    stu__mgr2__valid       =    pe2__stu__valid          ;
 assign    stu__mgr2__cntl        =    pe2__stu__cntl           ;
 assign    stu__pe2__ready        =    mgr2__stu__ready         ;
 assign    stu__mgr2__type        =    pe2__stu__type           ;
 assign    stu__mgr2__data        =    pe2__stu__data           ;
 assign    stu__mgr2__oob_data    =    pe2__stu__oob_data       ;

 assign    stu__mgr3__valid       =    pe3__stu__valid          ;
 assign    stu__mgr3__cntl        =    pe3__stu__cntl           ;
 assign    stu__pe3__ready        =    mgr3__stu__ready         ;
 assign    stu__mgr3__type        =    pe3__stu__type           ;
 assign    stu__mgr3__data        =    pe3__stu__data           ;
 assign    stu__mgr3__oob_data    =    pe3__stu__oob_data       ;

 assign    stu__mgr4__valid       =    pe4__stu__valid          ;
 assign    stu__mgr4__cntl        =    pe4__stu__cntl           ;
 assign    stu__pe4__ready        =    mgr4__stu__ready         ;
 assign    stu__mgr4__type        =    pe4__stu__type           ;
 assign    stu__mgr4__data        =    pe4__stu__data           ;
 assign    stu__mgr4__oob_data    =    pe4__stu__oob_data       ;

 assign    stu__mgr5__valid       =    pe5__stu__valid          ;
 assign    stu__mgr5__cntl        =    pe5__stu__cntl           ;
 assign    stu__pe5__ready        =    mgr5__stu__ready         ;
 assign    stu__mgr5__type        =    pe5__stu__type           ;
 assign    stu__mgr5__data        =    pe5__stu__data           ;
 assign    stu__mgr5__oob_data    =    pe5__stu__oob_data       ;

 assign    stu__mgr6__valid       =    pe6__stu__valid          ;
 assign    stu__mgr6__cntl        =    pe6__stu__cntl           ;
 assign    stu__pe6__ready        =    mgr6__stu__ready         ;
 assign    stu__mgr6__type        =    pe6__stu__type           ;
 assign    stu__mgr6__data        =    pe6__stu__data           ;
 assign    stu__mgr6__oob_data    =    pe6__stu__oob_data       ;

 assign    stu__mgr7__valid       =    pe7__stu__valid          ;
 assign    stu__mgr7__cntl        =    pe7__stu__cntl           ;
 assign    stu__pe7__ready        =    mgr7__stu__ready         ;
 assign    stu__mgr7__type        =    pe7__stu__type           ;
 assign    stu__mgr7__data        =    pe7__stu__data           ;
 assign    stu__mgr7__oob_data    =    pe7__stu__oob_data       ;

 assign    stu__mgr8__valid       =    pe8__stu__valid          ;
 assign    stu__mgr8__cntl        =    pe8__stu__cntl           ;
 assign    stu__pe8__ready        =    mgr8__stu__ready         ;
 assign    stu__mgr8__type        =    pe8__stu__type           ;
 assign    stu__mgr8__data        =    pe8__stu__data           ;
 assign    stu__mgr8__oob_data    =    pe8__stu__oob_data       ;

 assign    stu__mgr9__valid       =    pe9__stu__valid          ;
 assign    stu__mgr9__cntl        =    pe9__stu__cntl           ;
 assign    stu__pe9__ready        =    mgr9__stu__ready         ;
 assign    stu__mgr9__type        =    pe9__stu__type           ;
 assign    stu__mgr9__data        =    pe9__stu__data           ;
 assign    stu__mgr9__oob_data    =    pe9__stu__oob_data       ;

 assign    stu__mgr10__valid       =    pe10__stu__valid          ;
 assign    stu__mgr10__cntl        =    pe10__stu__cntl           ;
 assign    stu__pe10__ready        =    mgr10__stu__ready         ;
 assign    stu__mgr10__type        =    pe10__stu__type           ;
 assign    stu__mgr10__data        =    pe10__stu__data           ;
 assign    stu__mgr10__oob_data    =    pe10__stu__oob_data       ;

 assign    stu__mgr11__valid       =    pe11__stu__valid          ;
 assign    stu__mgr11__cntl        =    pe11__stu__cntl           ;
 assign    stu__pe11__ready        =    mgr11__stu__ready         ;
 assign    stu__mgr11__type        =    pe11__stu__type           ;
 assign    stu__mgr11__data        =    pe11__stu__data           ;
 assign    stu__mgr11__oob_data    =    pe11__stu__oob_data       ;

 assign    stu__mgr12__valid       =    pe12__stu__valid          ;
 assign    stu__mgr12__cntl        =    pe12__stu__cntl           ;
 assign    stu__pe12__ready        =    mgr12__stu__ready         ;
 assign    stu__mgr12__type        =    pe12__stu__type           ;
 assign    stu__mgr12__data        =    pe12__stu__data           ;
 assign    stu__mgr12__oob_data    =    pe12__stu__oob_data       ;

 assign    stu__mgr13__valid       =    pe13__stu__valid          ;
 assign    stu__mgr13__cntl        =    pe13__stu__cntl           ;
 assign    stu__pe13__ready        =    mgr13__stu__ready         ;
 assign    stu__mgr13__type        =    pe13__stu__type           ;
 assign    stu__mgr13__data        =    pe13__stu__data           ;
 assign    stu__mgr13__oob_data    =    pe13__stu__oob_data       ;

 assign    stu__mgr14__valid       =    pe14__stu__valid          ;
 assign    stu__mgr14__cntl        =    pe14__stu__cntl           ;
 assign    stu__pe14__ready        =    mgr14__stu__ready         ;
 assign    stu__mgr14__type        =    pe14__stu__type           ;
 assign    stu__mgr14__data        =    pe14__stu__data           ;
 assign    stu__mgr14__oob_data    =    pe14__stu__oob_data       ;

 assign    stu__mgr15__valid       =    pe15__stu__valid          ;
 assign    stu__mgr15__cntl        =    pe15__stu__cntl           ;
 assign    stu__pe15__ready        =    mgr15__stu__ready         ;
 assign    stu__mgr15__type        =    pe15__stu__type           ;
 assign    stu__mgr15__data        =    pe15__stu__data           ;
 assign    stu__mgr15__oob_data    =    pe15__stu__oob_data       ;

 assign    stu__mgr16__valid       =    pe16__stu__valid          ;
 assign    stu__mgr16__cntl        =    pe16__stu__cntl           ;
 assign    stu__pe16__ready        =    mgr16__stu__ready         ;
 assign    stu__mgr16__type        =    pe16__stu__type           ;
 assign    stu__mgr16__data        =    pe16__stu__data           ;
 assign    stu__mgr16__oob_data    =    pe16__stu__oob_data       ;

 assign    stu__mgr17__valid       =    pe17__stu__valid          ;
 assign    stu__mgr17__cntl        =    pe17__stu__cntl           ;
 assign    stu__pe17__ready        =    mgr17__stu__ready         ;
 assign    stu__mgr17__type        =    pe17__stu__type           ;
 assign    stu__mgr17__data        =    pe17__stu__data           ;
 assign    stu__mgr17__oob_data    =    pe17__stu__oob_data       ;

 assign    stu__mgr18__valid       =    pe18__stu__valid          ;
 assign    stu__mgr18__cntl        =    pe18__stu__cntl           ;
 assign    stu__pe18__ready        =    mgr18__stu__ready         ;
 assign    stu__mgr18__type        =    pe18__stu__type           ;
 assign    stu__mgr18__data        =    pe18__stu__data           ;
 assign    stu__mgr18__oob_data    =    pe18__stu__oob_data       ;

 assign    stu__mgr19__valid       =    pe19__stu__valid          ;
 assign    stu__mgr19__cntl        =    pe19__stu__cntl           ;
 assign    stu__pe19__ready        =    mgr19__stu__ready         ;
 assign    stu__mgr19__type        =    pe19__stu__type           ;
 assign    stu__mgr19__data        =    pe19__stu__data           ;
 assign    stu__mgr19__oob_data    =    pe19__stu__oob_data       ;

 assign    stu__mgr20__valid       =    pe20__stu__valid          ;
 assign    stu__mgr20__cntl        =    pe20__stu__cntl           ;
 assign    stu__pe20__ready        =    mgr20__stu__ready         ;
 assign    stu__mgr20__type        =    pe20__stu__type           ;
 assign    stu__mgr20__data        =    pe20__stu__data           ;
 assign    stu__mgr20__oob_data    =    pe20__stu__oob_data       ;

 assign    stu__mgr21__valid       =    pe21__stu__valid          ;
 assign    stu__mgr21__cntl        =    pe21__stu__cntl           ;
 assign    stu__pe21__ready        =    mgr21__stu__ready         ;
 assign    stu__mgr21__type        =    pe21__stu__type           ;
 assign    stu__mgr21__data        =    pe21__stu__data           ;
 assign    stu__mgr21__oob_data    =    pe21__stu__oob_data       ;

 assign    stu__mgr22__valid       =    pe22__stu__valid          ;
 assign    stu__mgr22__cntl        =    pe22__stu__cntl           ;
 assign    stu__pe22__ready        =    mgr22__stu__ready         ;
 assign    stu__mgr22__type        =    pe22__stu__type           ;
 assign    stu__mgr22__data        =    pe22__stu__data           ;
 assign    stu__mgr22__oob_data    =    pe22__stu__oob_data       ;

 assign    stu__mgr23__valid       =    pe23__stu__valid          ;
 assign    stu__mgr23__cntl        =    pe23__stu__cntl           ;
 assign    stu__pe23__ready        =    mgr23__stu__ready         ;
 assign    stu__mgr23__type        =    pe23__stu__type           ;
 assign    stu__mgr23__data        =    pe23__stu__data           ;
 assign    stu__mgr23__oob_data    =    pe23__stu__oob_data       ;

 assign    stu__mgr24__valid       =    pe24__stu__valid          ;
 assign    stu__mgr24__cntl        =    pe24__stu__cntl           ;
 assign    stu__pe24__ready        =    mgr24__stu__ready         ;
 assign    stu__mgr24__type        =    pe24__stu__type           ;
 assign    stu__mgr24__data        =    pe24__stu__data           ;
 assign    stu__mgr24__oob_data    =    pe24__stu__oob_data       ;

 assign    stu__mgr25__valid       =    pe25__stu__valid          ;
 assign    stu__mgr25__cntl        =    pe25__stu__cntl           ;
 assign    stu__pe25__ready        =    mgr25__stu__ready         ;
 assign    stu__mgr25__type        =    pe25__stu__type           ;
 assign    stu__mgr25__data        =    pe25__stu__data           ;
 assign    stu__mgr25__oob_data    =    pe25__stu__oob_data       ;

 assign    stu__mgr26__valid       =    pe26__stu__valid          ;
 assign    stu__mgr26__cntl        =    pe26__stu__cntl           ;
 assign    stu__pe26__ready        =    mgr26__stu__ready         ;
 assign    stu__mgr26__type        =    pe26__stu__type           ;
 assign    stu__mgr26__data        =    pe26__stu__data           ;
 assign    stu__mgr26__oob_data    =    pe26__stu__oob_data       ;

 assign    stu__mgr27__valid       =    pe27__stu__valid          ;
 assign    stu__mgr27__cntl        =    pe27__stu__cntl           ;
 assign    stu__pe27__ready        =    mgr27__stu__ready         ;
 assign    stu__mgr27__type        =    pe27__stu__type           ;
 assign    stu__mgr27__data        =    pe27__stu__data           ;
 assign    stu__mgr27__oob_data    =    pe27__stu__oob_data       ;

 assign    stu__mgr28__valid       =    pe28__stu__valid          ;
 assign    stu__mgr28__cntl        =    pe28__stu__cntl           ;
 assign    stu__pe28__ready        =    mgr28__stu__ready         ;
 assign    stu__mgr28__type        =    pe28__stu__type           ;
 assign    stu__mgr28__data        =    pe28__stu__data           ;
 assign    stu__mgr28__oob_data    =    pe28__stu__oob_data       ;

 assign    stu__mgr29__valid       =    pe29__stu__valid          ;
 assign    stu__mgr29__cntl        =    pe29__stu__cntl           ;
 assign    stu__pe29__ready        =    mgr29__stu__ready         ;
 assign    stu__mgr29__type        =    pe29__stu__type           ;
 assign    stu__mgr29__data        =    pe29__stu__data           ;
 assign    stu__mgr29__oob_data    =    pe29__stu__oob_data       ;

 assign    stu__mgr30__valid       =    pe30__stu__valid          ;
 assign    stu__mgr30__cntl        =    pe30__stu__cntl           ;
 assign    stu__pe30__ready        =    mgr30__stu__ready         ;
 assign    stu__mgr30__type        =    pe30__stu__type           ;
 assign    stu__mgr30__data        =    pe30__stu__data           ;
 assign    stu__mgr30__oob_data    =    pe30__stu__oob_data       ;

 assign    stu__mgr31__valid       =    pe31__stu__valid          ;
 assign    stu__mgr31__cntl        =    pe31__stu__cntl           ;
 assign    stu__pe31__ready        =    mgr31__stu__ready         ;
 assign    stu__mgr31__type        =    pe31__stu__type           ;
 assign    stu__mgr31__data        =    pe31__stu__data           ;
 assign    stu__mgr31__oob_data    =    pe31__stu__oob_data       ;

 assign    stu__mgr32__valid       =    pe32__stu__valid          ;
 assign    stu__mgr32__cntl        =    pe32__stu__cntl           ;
 assign    stu__pe32__ready        =    mgr32__stu__ready         ;
 assign    stu__mgr32__type        =    pe32__stu__type           ;
 assign    stu__mgr32__data        =    pe32__stu__data           ;
 assign    stu__mgr32__oob_data    =    pe32__stu__oob_data       ;

 assign    stu__mgr33__valid       =    pe33__stu__valid          ;
 assign    stu__mgr33__cntl        =    pe33__stu__cntl           ;
 assign    stu__pe33__ready        =    mgr33__stu__ready         ;
 assign    stu__mgr33__type        =    pe33__stu__type           ;
 assign    stu__mgr33__data        =    pe33__stu__data           ;
 assign    stu__mgr33__oob_data    =    pe33__stu__oob_data       ;

 assign    stu__mgr34__valid       =    pe34__stu__valid          ;
 assign    stu__mgr34__cntl        =    pe34__stu__cntl           ;
 assign    stu__pe34__ready        =    mgr34__stu__ready         ;
 assign    stu__mgr34__type        =    pe34__stu__type           ;
 assign    stu__mgr34__data        =    pe34__stu__data           ;
 assign    stu__mgr34__oob_data    =    pe34__stu__oob_data       ;

 assign    stu__mgr35__valid       =    pe35__stu__valid          ;
 assign    stu__mgr35__cntl        =    pe35__stu__cntl           ;
 assign    stu__pe35__ready        =    mgr35__stu__ready         ;
 assign    stu__mgr35__type        =    pe35__stu__type           ;
 assign    stu__mgr35__data        =    pe35__stu__data           ;
 assign    stu__mgr35__oob_data    =    pe35__stu__oob_data       ;

 assign    stu__mgr36__valid       =    pe36__stu__valid          ;
 assign    stu__mgr36__cntl        =    pe36__stu__cntl           ;
 assign    stu__pe36__ready        =    mgr36__stu__ready         ;
 assign    stu__mgr36__type        =    pe36__stu__type           ;
 assign    stu__mgr36__data        =    pe36__stu__data           ;
 assign    stu__mgr36__oob_data    =    pe36__stu__oob_data       ;

 assign    stu__mgr37__valid       =    pe37__stu__valid          ;
 assign    stu__mgr37__cntl        =    pe37__stu__cntl           ;
 assign    stu__pe37__ready        =    mgr37__stu__ready         ;
 assign    stu__mgr37__type        =    pe37__stu__type           ;
 assign    stu__mgr37__data        =    pe37__stu__data           ;
 assign    stu__mgr37__oob_data    =    pe37__stu__oob_data       ;

 assign    stu__mgr38__valid       =    pe38__stu__valid          ;
 assign    stu__mgr38__cntl        =    pe38__stu__cntl           ;
 assign    stu__pe38__ready        =    mgr38__stu__ready         ;
 assign    stu__mgr38__type        =    pe38__stu__type           ;
 assign    stu__mgr38__data        =    pe38__stu__data           ;
 assign    stu__mgr38__oob_data    =    pe38__stu__oob_data       ;

 assign    stu__mgr39__valid       =    pe39__stu__valid          ;
 assign    stu__mgr39__cntl        =    pe39__stu__cntl           ;
 assign    stu__pe39__ready        =    mgr39__stu__ready         ;
 assign    stu__mgr39__type        =    pe39__stu__type           ;
 assign    stu__mgr39__data        =    pe39__stu__data           ;
 assign    stu__mgr39__oob_data    =    pe39__stu__oob_data       ;

 assign    stu__mgr40__valid       =    pe40__stu__valid          ;
 assign    stu__mgr40__cntl        =    pe40__stu__cntl           ;
 assign    stu__pe40__ready        =    mgr40__stu__ready         ;
 assign    stu__mgr40__type        =    pe40__stu__type           ;
 assign    stu__mgr40__data        =    pe40__stu__data           ;
 assign    stu__mgr40__oob_data    =    pe40__stu__oob_data       ;

 assign    stu__mgr41__valid       =    pe41__stu__valid          ;
 assign    stu__mgr41__cntl        =    pe41__stu__cntl           ;
 assign    stu__pe41__ready        =    mgr41__stu__ready         ;
 assign    stu__mgr41__type        =    pe41__stu__type           ;
 assign    stu__mgr41__data        =    pe41__stu__data           ;
 assign    stu__mgr41__oob_data    =    pe41__stu__oob_data       ;

 assign    stu__mgr42__valid       =    pe42__stu__valid          ;
 assign    stu__mgr42__cntl        =    pe42__stu__cntl           ;
 assign    stu__pe42__ready        =    mgr42__stu__ready         ;
 assign    stu__mgr42__type        =    pe42__stu__type           ;
 assign    stu__mgr42__data        =    pe42__stu__data           ;
 assign    stu__mgr42__oob_data    =    pe42__stu__oob_data       ;

 assign    stu__mgr43__valid       =    pe43__stu__valid          ;
 assign    stu__mgr43__cntl        =    pe43__stu__cntl           ;
 assign    stu__pe43__ready        =    mgr43__stu__ready         ;
 assign    stu__mgr43__type        =    pe43__stu__type           ;
 assign    stu__mgr43__data        =    pe43__stu__data           ;
 assign    stu__mgr43__oob_data    =    pe43__stu__oob_data       ;

 assign    stu__mgr44__valid       =    pe44__stu__valid          ;
 assign    stu__mgr44__cntl        =    pe44__stu__cntl           ;
 assign    stu__pe44__ready        =    mgr44__stu__ready         ;
 assign    stu__mgr44__type        =    pe44__stu__type           ;
 assign    stu__mgr44__data        =    pe44__stu__data           ;
 assign    stu__mgr44__oob_data    =    pe44__stu__oob_data       ;

 assign    stu__mgr45__valid       =    pe45__stu__valid          ;
 assign    stu__mgr45__cntl        =    pe45__stu__cntl           ;
 assign    stu__pe45__ready        =    mgr45__stu__ready         ;
 assign    stu__mgr45__type        =    pe45__stu__type           ;
 assign    stu__mgr45__data        =    pe45__stu__data           ;
 assign    stu__mgr45__oob_data    =    pe45__stu__oob_data       ;

 assign    stu__mgr46__valid       =    pe46__stu__valid          ;
 assign    stu__mgr46__cntl        =    pe46__stu__cntl           ;
 assign    stu__pe46__ready        =    mgr46__stu__ready         ;
 assign    stu__mgr46__type        =    pe46__stu__type           ;
 assign    stu__mgr46__data        =    pe46__stu__data           ;
 assign    stu__mgr46__oob_data    =    pe46__stu__oob_data       ;

 assign    stu__mgr47__valid       =    pe47__stu__valid          ;
 assign    stu__mgr47__cntl        =    pe47__stu__cntl           ;
 assign    stu__pe47__ready        =    mgr47__stu__ready         ;
 assign    stu__mgr47__type        =    pe47__stu__type           ;
 assign    stu__mgr47__data        =    pe47__stu__data           ;
 assign    stu__mgr47__oob_data    =    pe47__stu__oob_data       ;

 assign    stu__mgr48__valid       =    pe48__stu__valid          ;
 assign    stu__mgr48__cntl        =    pe48__stu__cntl           ;
 assign    stu__pe48__ready        =    mgr48__stu__ready         ;
 assign    stu__mgr48__type        =    pe48__stu__type           ;
 assign    stu__mgr48__data        =    pe48__stu__data           ;
 assign    stu__mgr48__oob_data    =    pe48__stu__oob_data       ;

 assign    stu__mgr49__valid       =    pe49__stu__valid          ;
 assign    stu__mgr49__cntl        =    pe49__stu__cntl           ;
 assign    stu__pe49__ready        =    mgr49__stu__ready         ;
 assign    stu__mgr49__type        =    pe49__stu__type           ;
 assign    stu__mgr49__data        =    pe49__stu__data           ;
 assign    stu__mgr49__oob_data    =    pe49__stu__oob_data       ;

 assign    stu__mgr50__valid       =    pe50__stu__valid          ;
 assign    stu__mgr50__cntl        =    pe50__stu__cntl           ;
 assign    stu__pe50__ready        =    mgr50__stu__ready         ;
 assign    stu__mgr50__type        =    pe50__stu__type           ;
 assign    stu__mgr50__data        =    pe50__stu__data           ;
 assign    stu__mgr50__oob_data    =    pe50__stu__oob_data       ;

 assign    stu__mgr51__valid       =    pe51__stu__valid          ;
 assign    stu__mgr51__cntl        =    pe51__stu__cntl           ;
 assign    stu__pe51__ready        =    mgr51__stu__ready         ;
 assign    stu__mgr51__type        =    pe51__stu__type           ;
 assign    stu__mgr51__data        =    pe51__stu__data           ;
 assign    stu__mgr51__oob_data    =    pe51__stu__oob_data       ;

 assign    stu__mgr52__valid       =    pe52__stu__valid          ;
 assign    stu__mgr52__cntl        =    pe52__stu__cntl           ;
 assign    stu__pe52__ready        =    mgr52__stu__ready         ;
 assign    stu__mgr52__type        =    pe52__stu__type           ;
 assign    stu__mgr52__data        =    pe52__stu__data           ;
 assign    stu__mgr52__oob_data    =    pe52__stu__oob_data       ;

 assign    stu__mgr53__valid       =    pe53__stu__valid          ;
 assign    stu__mgr53__cntl        =    pe53__stu__cntl           ;
 assign    stu__pe53__ready        =    mgr53__stu__ready         ;
 assign    stu__mgr53__type        =    pe53__stu__type           ;
 assign    stu__mgr53__data        =    pe53__stu__data           ;
 assign    stu__mgr53__oob_data    =    pe53__stu__oob_data       ;

 assign    stu__mgr54__valid       =    pe54__stu__valid          ;
 assign    stu__mgr54__cntl        =    pe54__stu__cntl           ;
 assign    stu__pe54__ready        =    mgr54__stu__ready         ;
 assign    stu__mgr54__type        =    pe54__stu__type           ;
 assign    stu__mgr54__data        =    pe54__stu__data           ;
 assign    stu__mgr54__oob_data    =    pe54__stu__oob_data       ;

 assign    stu__mgr55__valid       =    pe55__stu__valid          ;
 assign    stu__mgr55__cntl        =    pe55__stu__cntl           ;
 assign    stu__pe55__ready        =    mgr55__stu__ready         ;
 assign    stu__mgr55__type        =    pe55__stu__type           ;
 assign    stu__mgr55__data        =    pe55__stu__data           ;
 assign    stu__mgr55__oob_data    =    pe55__stu__oob_data       ;

 assign    stu__mgr56__valid       =    pe56__stu__valid          ;
 assign    stu__mgr56__cntl        =    pe56__stu__cntl           ;
 assign    stu__pe56__ready        =    mgr56__stu__ready         ;
 assign    stu__mgr56__type        =    pe56__stu__type           ;
 assign    stu__mgr56__data        =    pe56__stu__data           ;
 assign    stu__mgr56__oob_data    =    pe56__stu__oob_data       ;

 assign    stu__mgr57__valid       =    pe57__stu__valid          ;
 assign    stu__mgr57__cntl        =    pe57__stu__cntl           ;
 assign    stu__pe57__ready        =    mgr57__stu__ready         ;
 assign    stu__mgr57__type        =    pe57__stu__type           ;
 assign    stu__mgr57__data        =    pe57__stu__data           ;
 assign    stu__mgr57__oob_data    =    pe57__stu__oob_data       ;

 assign    stu__mgr58__valid       =    pe58__stu__valid          ;
 assign    stu__mgr58__cntl        =    pe58__stu__cntl           ;
 assign    stu__pe58__ready        =    mgr58__stu__ready         ;
 assign    stu__mgr58__type        =    pe58__stu__type           ;
 assign    stu__mgr58__data        =    pe58__stu__data           ;
 assign    stu__mgr58__oob_data    =    pe58__stu__oob_data       ;

 assign    stu__mgr59__valid       =    pe59__stu__valid          ;
 assign    stu__mgr59__cntl        =    pe59__stu__cntl           ;
 assign    stu__pe59__ready        =    mgr59__stu__ready         ;
 assign    stu__mgr59__type        =    pe59__stu__type           ;
 assign    stu__mgr59__data        =    pe59__stu__data           ;
 assign    stu__mgr59__oob_data    =    pe59__stu__oob_data       ;

 assign    stu__mgr60__valid       =    pe60__stu__valid          ;
 assign    stu__mgr60__cntl        =    pe60__stu__cntl           ;
 assign    stu__pe60__ready        =    mgr60__stu__ready         ;
 assign    stu__mgr60__type        =    pe60__stu__type           ;
 assign    stu__mgr60__data        =    pe60__stu__data           ;
 assign    stu__mgr60__oob_data    =    pe60__stu__oob_data       ;

 assign    stu__mgr61__valid       =    pe61__stu__valid          ;
 assign    stu__mgr61__cntl        =    pe61__stu__cntl           ;
 assign    stu__pe61__ready        =    mgr61__stu__ready         ;
 assign    stu__mgr61__type        =    pe61__stu__type           ;
 assign    stu__mgr61__data        =    pe61__stu__data           ;
 assign    stu__mgr61__oob_data    =    pe61__stu__oob_data       ;

 assign    stu__mgr62__valid       =    pe62__stu__valid          ;
 assign    stu__mgr62__cntl        =    pe62__stu__cntl           ;
 assign    stu__pe62__ready        =    mgr62__stu__ready         ;
 assign    stu__mgr62__type        =    pe62__stu__type           ;
 assign    stu__mgr62__data        =    pe62__stu__data           ;
 assign    stu__mgr62__oob_data    =    pe62__stu__oob_data       ;

 assign    stu__mgr63__valid       =    pe63__stu__valid          ;
 assign    stu__mgr63__cntl        =    pe63__stu__cntl           ;
 assign    stu__pe63__ready        =    mgr63__stu__ready         ;
 assign    stu__mgr63__type        =    pe63__stu__type           ;
 assign    stu__mgr63__data        =    pe63__stu__data           ;
 assign    stu__mgr63__oob_data    =    pe63__stu__oob_data       ;

