
  // Send an 'all' synchronized to all PE's 
  // pe__sys__thisSyncnronized basically means all the streams in a PE are complete
  // The PE controller will move to a 'final' state once it receives sys__pe__allSynchronized
  assign  DownstreamStackBusOOB[0].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[1].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[2].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[3].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[4].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[5].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[6].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[7].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[8].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[9].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[10].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[11].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[12].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[13].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[14].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[15].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[16].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[17].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[18].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[19].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[20].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[21].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[22].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[23].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[24].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[25].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[26].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[27].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[28].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[29].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[30].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[31].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[32].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[33].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[34].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[35].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[36].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[37].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[38].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[39].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[40].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[41].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[42].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[43].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[44].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[45].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[46].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[47].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[48].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[49].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[50].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[51].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[52].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[53].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[54].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[55].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[56].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[57].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[58].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[59].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[60].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[61].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[62].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 

  assign  DownstreamStackBusOOB[63].sys__pe__allSynchronized = DownstreamStackBusOOB[0].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[1].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[2].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[3].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[4].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[5].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[6].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[7].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[8].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[9].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[10].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[11].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[12].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[13].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[14].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[15].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[16].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[17].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[18].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[19].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[20].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[21].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[22].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[23].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[24].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[25].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[26].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[27].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[28].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[29].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[30].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[31].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[32].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[33].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[34].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[35].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[36].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[37].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[38].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[39].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[40].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[41].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[42].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[43].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[44].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[45].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[46].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[47].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[48].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[49].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[50].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[51].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[52].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[53].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[54].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[55].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[56].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[57].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[58].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[59].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[60].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[61].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[62].pe__sys__thisSynchronized & 
                                   DownstreamStackBusOOB[63].pe__sys__thisSynchronized ; 
