`ifndef _manager_vh
`define _manager_vh

/*****************************************************************

    File name   : manager.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : Mar 2017
    email       : lbbaker@ncsu.edu

*****************************************************************/


//------------------------------------------------
// System
//------------------------------------------------
`define MGR_MGR_ID_WIDTH             (`CLOG2(`MGR_ARRAY_NUM_OF_MGR))
`define MGR_MGR_ID_MSB               (`MGR_MGR_ID_WIDTH-1)
`define MGR_MGR_ID_LSB               0
`define MGR_MGR_ID_SIZE              (`MGR_MGR_ID_MSB - `MGR_MGR_ID_LSB +1)
`define MGR_MGR_ID_RANGE              `MGR_MGR_ID_MSB : `MGR_MGR_ID_LSB

`define MGR_MGR_ID_BITMASK_WIDTH             `MGR_ARRAY_NUM_OF_MGR
`define MGR_MGR_ID_BITMASK_MSB               (`MGR_MGR_ID_BITMASK_WIDTH-1)
`define MGR_MGR_ID_BITMASK_LSB               0
`define MGR_MGR_ID_BITMASK_SIZE              (`MGR_MGR_ID_BITMASK_MSB - `MGR_MGR_ID_BITMASK_LSB +1)
`define MGR_MGR_ID_BITMASK_RANGE              `MGR_MGR_ID_BITMASK_MSB : `MGR_MGR_ID_BITMASK_LSB
//------------------------------------------------
// Stack Bus stream
//------------------------------------------------

`define MGR_INITIAL_TAG          'h81

// we will carry a tag to track result (to possibly support multiple operations before first result is returned)
`define MGR_STD_OOB_TAG_WIDTH          `PE_STD_OOB_TAG_WIDTH
`define MGR_STD_OOB_TAG_MSB            `MGR_STD_OOB_TAG_WIDTH-1
`define MGR_STD_OOB_TAG_LSB            0
`define MGR_STD_OOB_TAG_RANGE          `MGR_STD_OOB_TAG_MSB : `MGR_STD_OOB_TAG_LSB

`define MGR_STD_LANE_DATA_WIDTH          `STACK_DOWN_INTF_STRM_DATA_WIDTH 
`define MGR_STD_LANE_DATA_MSB            `MGR_STD_LANE_DATA_WIDTH-1
`define MGR_STD_LANE_DATA_LSB            0
`define MGR_STD_LANE_DATA_RANGE          `MGR_STD_LANE_DATA_MSB : `MGR_STD_LANE_DATA_LSB

`define MGR_STU_DATA_WIDTH          `STACK_UP_INTF_DATA_WIDTH 
`define MGR_STU_DATA_MSB            `MGR_STU_DATA_WIDTH-1
`define MGR_STU_DATA_LSB            0
`define MGR_STU_DATA_RANGE          `MGR_STU_DATA_MSB : `MGR_STU_DATA_LSB



//------------------------------------------------
// MGR Stack bus streams
//------------------------------------------------

`define MGR_NUM_OF_STREAMS               `PE_NUM_OF_STREAMS 
`define MGR_NUM_OF_STREAMS_MSB           (`MGR_NUM_OF_STREAMS -1)
`define MGR_NUM_OF_STREAMS_LSB            0
`define MGR_NUM_OF_STREAMS_SIZE           (`MGR_NUM_OF_STREAMS_MSB - `MGR_NUM_OF_STREAMS_LSB +1)
`define MGR_NUM_OF_STREAMS_RANGE           `MGR_NUM_OF_STREAMS_MSB : `MGR_NUM_OF_STREAMS_LSB
`define MGR_NUM_OF_STREAMS_VECTOR        `PE_NUM_OF_STREAMS-1 : 0

`define MGR_STREAM_ADDRESS_WIDTH          (`CLOG2(`MGR_NUM_OF_STREAMS))
`define MGR_STREAM_ADDRESS_MSB           `MGR_STREAM_ADDRESS_WIDTH-1
`define MGR_STREAM_ADDRESS_LSB            0
`define MGR_STREAM_ADDRESS_SIZE           (`MGR_STREAM_ADDRESS_MSB - `MGR_STREAM_ADDRESS_LSB +1)
`define MGR_STREAM_ADDRESS_RANGE           `MGR_STREAM_ADDRESS_MSB : `MGR_STREAM_ADDRESS_LSB
//------------------------------------------------
// MGR Execution Lane 
//------------------------------------------------

`define MGR_NUM_OF_EXEC_LANES               `PE_NUM_OF_EXEC_LANES
`define MGR_NUM_OF_EXEC_LANES_MSB           (`MGR_NUM_OF_EXEC_LANES -1)
`define MGR_NUM_OF_EXEC_LANES_LSB            0
`define MGR_NUM_OF_EXEC_LANES_SIZE           (`MGR_NUM_OF_EXEC_LANES_MSB - `MGR_NUM_OF_EXEC_LANES_LSB +1)
`define MGR_NUM_OF_EXEC_LANES_RANGE           `MGR_NUM_OF_EXEC_LANES_MSB : `MGR_NUM_OF_EXEC_LANES_LSB

`define MGR_EXEC_LANE_WIDTH               `PE_EXEC_LANE_WIDTH
`define MGR_EXEC_LANE_WIDTH_MSB           `MGR_EXEC_LANE_WIDTH-1
`define MGR_EXEC_LANE_WIDTH_LSB            0
`define MGR_EXEC_LANE_WIDTH_SIZE           (`MGR_EXEC_LANE_WIDTH_MSB - `MGR_EXEC_LANE_WIDTH_LSB +1)
`define MGR_EXEC_LANE_WIDTH_RANGE           `MGR_EXEC_LANE_WIDTH_MSB : `MGR_EXEC_LANE_WIDTH_LSB

`define MGR_EXEC_LANE_ID_WIDTH            `PE_EXEC_LANE_ID_WIDTH   
`define MGR_EXEC_LANE_ID_MSB              `PE_EXEC_LANE_ID_MSB     
`define MGR_EXEC_LANE_ID_LSB              `PE_EXEC_LANE_ID_LSB     
`define MGR_EXEC_LANE_ID_RANGE            `PE_EXEC_LANE_ID_RANGE   

//--------------------------------------------------------
// In cases where we set number of active lanes, Number of active lanes is 1..32, so need 6 bits
  
`define MGR_NUM_LANES_WIDTH               (`CLOG2(`PE_NUM_OF_EXEC_LANES))+1
`define MGR_NUM_LANES_MSB           `MGR_NUM_LANES_WIDTH-1
`define MGR_NUM_LANES_LSB            0
`define MGR_NUM_LANES_SIZE           (`MGR_NUM_LANES_MSB - `MGR_NUM_LANES_LSB +1)
`define MGR_NUM_LANES_RANGE           `MGR_NUM_LANES_MSB : `MGR_NUM_LANES_LSB
//---------------------------------------------------------------------------------------------------------------------
// Memory

//---------------------------------------------------------------------------------------------------------------------
// WU Memory

// FIXME
`define MGR_WU_MEMORY_DEPTH                      4096
`define MGR_WU_ADDRESS_WIDTH                       (`CLOG2(`MGR_WU_MEMORY_DEPTH))
`define MGR_WU_ADDRESS_MSB                         `MGR_WU_ADDRESS_WIDTH-1
`define MGR_WU_ADDRESS_LSB                         0
`define MGR_WU_ADDRESS_SIZE                        (`MGR_WU_ADDRESS_MSB - `MGR_WU_ADDRESS_LSB +1)
`define MGR_WU_ADDRESS_RANGE                        `MGR_WU_ADDRESS_MSB : `MGR_WU_ADDRESS_LSB

`define MGR_WU_MEMORY_INIT_ENTRIES               16  // DEBUG: numner of initial instruction memory loads


//---------------------------------------------------------------------------------------------------------------------
// WU Instruction

`define MGR_WU_DESC_PER_INST                       4
`define MGR_WU_DESC_PER_INST_WIDTH                 (`CLOG2(`MGR_WU_DESC_PER_INST ))
`define MGR_WU_DESC_PER_INST_MSB                   `MGR_WU_DESC_PER_INST_WIDTH-1
`define MGR_WU_DESC_PER_INST_LSB                   0
`define MGR_WU_DESC_PER_INST_SIZE                  (`MGR_WU_DESC_PER_INST_MSB - `MGR_WU_DESC_PER_INST_LSB +1)
`define MGR_WU_DESC_PER_INST_RANGE                  `MGR_WU_DESC_PER_INST_MSB : `MGR_WU_DESC_PER_INST_LSB

`define MGR_WU_OPT_PER_INST                       3
`define MGR_WU_OPT_PER_INST_WIDTH                 `MGR_WU_OPT_PER_INST   
`define MGR_WU_OPT_PER_INST_MSB                   `MGR_WU_OPT_PER_INST_WIDTH-1
`define MGR_WU_OPT_PER_INST_LSB                   0
`define MGR_WU_OPT_PER_INST_SIZE                  (`MGR_WU_OPT_PER_INST_MSB - `MGR_WU_OPT_PER_INST_LSB +1)
`define MGR_WU_OPT_PER_INST_RANGE                  `MGR_WU_OPT_PER_INST_MSB : `MGR_WU_OPT_PER_INST_LSB


`define MGR_WU_OPT_TYPE_WIDTH                 8
`define MGR_WU_OPT_TYPE_MSB                   `MGR_WU_OPT_TYPE_WIDTH-1
`define MGR_WU_OPT_TYPE_LSB                   0
`define MGR_WU_OPT_TYPE_SIZE                  (`MGR_WU_OPT_TYPE_MSB - `MGR_WU_OPT_TYPE_LSB +1)
`define MGR_WU_OPT_TYPE_RANGE                  `MGR_WU_OPT_TYPE_MSB : `MGR_WU_OPT_TYPE_LSB


`define MGR_WU_OPT_VALUE_WIDTH                 8
`define MGR_WU_OPT_VALUE_MSB                   `MGR_WU_OPT_VALUE_WIDTH-1
`define MGR_WU_OPT_VALUE_LSB                   0
`define MGR_WU_OPT_VALUE_SIZE                  (`MGR_WU_OPT_VALUE_MSB - `MGR_WU_OPT_VALUE_LSB +1)
`define MGR_WU_OPT_VALUE_RANGE                  `MGR_WU_OPT_VALUE_MSB : `MGR_WU_OPT_VALUE_LSB


`define MGR_WU_EXTD_OPT_VALUE_WIDTH                 `MGR_WU_OPT_VALUE_WIDTH  *3
`define MGR_WU_EXTD_OPT_VALUE_MSB                   `MGR_WU_EXTD_OPT_VALUE_WIDTH-1
`define MGR_WU_EXTD_OPT_VALUE_LSB                   0
`define MGR_WU_EXTD_OPT_VALUE_SIZE                  (`MGR_WU_EXTD_OPT_VALUE_MSB - `MGR_WU_EXTD_OPT_VALUE_LSB +1)
`define MGR_WU_EXTD_OPT_VALUE_RANGE                  `MGR_WU_EXTD_OPT_VALUE_MSB : `MGR_WU_EXTD_OPT_VALUE_LSB

`define MGR_WU_TUPLE_WIDTH                 `MGR_WU_OPT_TYPE_WIDTH+`MGR_WU_OPT_VALUE_WIDTH
`define MGR_WU_TUPLE_MSB                   `MGR_WU_TUPLE_WIDTH-1
`define MGR_WU_TUPLE_LSB                   0
`define MGR_WU_TUPLE_SIZE                  (`MGR_WU_TUPLE_MSB - `MGR_WU_TUPLE_LSB +1)
`define MGR_WU_TUPLE_RANGE                  `MGR_WU_TUPLE_MSB : `MGR_WU_TUPLE_LSB

`define MGR_WU_EXTD_TUPLE_WIDTH            `MGR_WU_OPT_TYPE_WIDTH+`MGR_WU_EXTD_OPT_VALUE_WIDTH
`define MGR_WU_EXTD_TUPLE_MSB              `MGR_WU_EXTD_TUPLE_WIDTH-1
`define MGR_WU_EXTD_TUPLE_LSB              0
`define MGR_WU_EXTD_TUPLE_SIZE             (`MGR_WU_EXTD_TUPLE_MSB - `MGR_WU_EXTD_TUPLE_LSB +1)
`define MGR_WU_EXTD_TUPLE_RANGE             `MGR_WU_EXTD_TUPLE_MSB : `MGR_WU_EXTD_TUPLE_LSB

`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB              `MGR_WU_EXTD_TUPLE_MSB
`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB              `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB-(`MGR_WU_OPT_TYPE_WIDTH-1)                 
`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_SIZE             (`MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB - `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB +1)
`define MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_RANGE             `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_MSB : `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB

`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB              `MGR_WU_EXTD_TUPLE_OPT_TYPE_FIELD_LSB-1
`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_LSB              `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB-(`MGR_WU_EXTD_OPT_VALUE_WIDTH-1)
`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_SIZE             (`MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB - `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_LSB +1)
`define MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_RANGE             `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_MSB : `MGR_WU_EXTD_TUPLE_OPT_VAL_FIELD_LSB

//------------------------------------------------------------------------------------------------------------------------------------------------------
// Extended Tuple Mode Registers
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT      1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE     2
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_FLUSH     3


`define MGR_WU_EXTD_TUPLE_MODE_REG_TXFER_INST_DNLD   0
`define MGR_WU_EXTD_TUPLE_MODE_REG_TXFER_GROUP_DNLD  1
`define MGR_WU_EXTD_TUPLE_MODE_REG_TXFER_MEM_DNLD    2
`define MGR_WU_EXTD_TUPLE_MODE_REG_TXFER_MEM_UPLD    3

`define MGR_WU_CONFIG_MODE_REG_ID_WIDTH    3
`define MGR_WU_CONFIG_MODE_REG_ID_MSB      `MGR_WU_CONFIG_MODE_REG_ID_WIDTH-1
`define MGR_WU_CONFIG_MODE_REG_ID_LSB      0
`define MGR_WU_CONFIG_MODE_REG_ID_SIZE     (`MGR_WU_CONFIG_MODE_REG_ID_MSB - `MGR_WU_CONFIG_MODE_REG_ID_LSB +1)
`define MGR_WU_CONFIG_MODE_REG_ID_RANGE     `MGR_WU_CONFIG_MODE_REG_ID_MSB : `MGR_WU_CONFIG_MODE_REG_ID_LSB

`define MGR_WU_CONFIG_MODE_REG_VAL_WIDTH    21
`define MGR_WU_CONFIG_MODE_REG_VAL_MSB      `MGR_WU_CONFIG_MODE_REG_VAL_WIDTH-1
`define MGR_WU_CONFIG_MODE_REG_VAL_LSB      0
`define MGR_WU_CONFIG_MODE_REG_VAL_SIZE     (`MGR_WU_CONFIG_MODE_REG_VAL_MSB - `MGR_WU_CONFIG_MODE_REG_VAL_LSB +1)
`define MGR_WU_CONFIG_MODE_REG_VAL_RANGE     `MGR_WU_CONFIG_MODE_REG_VAL_MSB : `MGR_WU_CONFIG_MODE_REG_VAL_LSB


`define MGR_WU_EXTD_TUPLE_MODE_REG_VAL_WIDTH    21
`define MGR_WU_EXTD_TUPLE_MODE_REG_VAL_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_VAL_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_VAL_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_VAL_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_VAL_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_VAL_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_VAL_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_VAL_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_VAL_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_ID_WIDTH    3
`define MGR_WU_EXTD_TUPLE_MODE_REG_ID_MSB      ((`MGR_WU_EXTD_TUPLE_MODE_REG_ID_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_ID_WIDTH)-1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_ID_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_VAL_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_ID_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_ID_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_ID_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_ID_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_ID_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_ID_LSB


// INSTRUCTION DNLD
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_WIDTH    1
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_WIDTH      7
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_CONT_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_WIDTH      13
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NA_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_INST_DNLD_NUM_OF_WORDS_LSB


// GROUP DNLD
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_WIDTH    1
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_WIDTH      7
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_CONT_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_WIDTH      8
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NA_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_GRP_DNLD_NUM_OF_GRPS_LSB


// MEMORY DNLD
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_WIDTH    21
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_DNLD_CONT_LSB

// MEMORY UPLD
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_WIDTH    21
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_MEM_UPLD_CONT_LSB



// SEND
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_WIDTH    1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_WIDTH      1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_HOST_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_WIDTH      `MGR_NOC_MCAST_GROUP_PTR_WIDTH
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ALL_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_WIDTH      `MGR_NOC_MCAST_GROUP_PTR_WIDTH
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_GRP_PTR_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_SEND_ENA_LSB

// WAIT
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_WIDTH    1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_WIDTH      1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_HOST_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_WIDTH      `MGR_NOC_MCAST_GROUP_PTR_WIDTH
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ALL_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_WIDTH      `MGR_NOC_MCAST_GROUP_PTR_WIDTH
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_GRP_PTR_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_WAIT_ENA_LSB

// PAUSE
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_WIDTH    1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_MSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_WIDTH-1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_LSB      0
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_WIDTH      8
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_INDEF_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_LSB

`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_WIDTH    12
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_MSB      (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_LSB+`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_WIDTH) -1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_LSB      `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_NA_MSB+1
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_SIZE     (`MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_MSB - `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_LSB +1)
`define MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_RANGE     `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_MSB : `MGR_WU_EXTD_TUPLE_MODE_REG_SYNC_PAUSE_COUNT_LSB



//------------------------------------------------------------------------------------------------------------------------------------------------------



// Instruction fields
`define MGR_INST_TYPE_WIDTH               5
`define MGR_INST_TYPE_MSB                `MGR_INST_TYPE_WIDTH-1
`define MGR_INST_TYPE_LSB                 0
`define MGR_INST_TYPE_SIZE              (`MGR_INST_TYPE_MSB - `MGR_INST_TYPE_LSB +1)
`define MGR_INST_TYPE_RANGE              `MGR_INST_TYPE_MSB : `MGR_INST_TYPE_LSB

//-------------------------------------------------------------
// Operands

`define MGR_OP_MAX_NUM_OF_OPERANDS    16384

`define MGR_OP_MAX_NUM_OF_OPERANDS_WIDTH        (`CLOG2(`MGR_OP_MAX_NUM_OF_OPERANDS ))
`define MGR_OP_MAX_NUM_OF_OPERANDS_MSB          `MGR_OP_MAX_NUM_OF_OPERANDS_WIDTH-1
`define MGR_OP_MAX_NUM_OF_OPERANDS_LSB          0
`define MGR_OP_MAX_NUM_OF_OPERANDS_SIZE         (`MGR_OP_MAX_NUM_OF_OPERANDS_MSB - `MGR_OP_MAX_NUM_OF_OPERANDS_LSB +1)
`define MGR_OP_MAX_NUM_OF_OPERANDS_RANGE         `MGR_OP_MAX_NUM_OF_OPERANDS_MSB : `MGR_OP_MAX_NUM_OF_OPERANDS_LSB

//-------------------------------------------------------------
//-------------------------------------------------------------
//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_desc_type
`define MGR_INST_DESC_TYPE_NOP              0
`define MGR_INST_DESC_TYPE_OP               1
`define MGR_INST_DESC_TYPE_MR               2
`define MGR_INST_DESC_TYPE_MW               3
`define MGR_INST_DESC_TYPE_CFG              4
`define MGR_INST_DESC_TYPE_STATUS           5

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_option_type
`define MGR_INST_OPTION_TYPE_NOP                    0
`define MGR_INST_OPTION_TYPE_SRC                    1
`define MGR_INST_OPTION_TYPE_TGT                    2
`define MGR_INST_OPTION_TYPE_TXFER                  3
`define MGR_INST_OPTION_TYPE_NUM_OF_LANES           4
`define MGR_INST_OPTION_TYPE_STOP                   5
`define MGR_INST_OPTION_TYPE_SIMDOP                 6
`define MGR_INST_OPTION_TYPE_MEMORY                 7
`define MGR_INST_OPTION_TYPE_NUM_OF_ARG0_OPERANDS   8
`define MGR_INST_OPTION_TYPE_NUM_OF_ARG1_OPERANDS   9
`define MGR_INST_OPTION_TYPE_CFG_SYNC              10
`define MGR_INST_OPTION_TYPE_CFG_DATA              11
`define MGR_INST_OPTION_TYPE_STATUS                12

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_simd_type
`define MGR_INST_OPTION_SIMD_TYPE_NOP       0
`define MGR_INST_OPTION_SIMD_TYPE_RELU      1

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_stOp_type
`define MGR_INST_OPTION_STOP_TYPE_NOP                                                  0
`define MGR_INST_OPTION_STOP_TYPE_STREAMING_OP_CNTL_OPERATION_STD_STD_FP_MAC_TO_MEM    1
`define MGR_INST_OPTION_STOP_TYPE_STREAMING_OP_CNTL_OPERATION_STD_NONE_NOP_TO_MEM      2
`define MGR_INST_OPTION_STOP_TYPE_STREAMING_OP_CNTL_OPERATION_MEM_STD_FP_MAC_TO_MEM    3

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_target_type
`define MGR_INST_OPTION_TGT_TYPE_STACK_DN_ARG0   0
`define MGR_INST_OPTION_TGT_TYPE_STACK_DN_ARG1   1
`define MGR_INST_OPTION_TGT_TYPE_STACK_UP        2
`define MGR_INST_OPTION_TGT_TYPE_NOC             3
`define MGR_INST_OPTION_TGT_TYPE_NOP             7


`define MGR_INST_OPTION_TGT_WIDTH        3
`define MGR_INST_OPTION_TGT_MSB          `MGR_INST_OPTION_TGT_WIDTH-1
`define MGR_INST_OPTION_TGT_LSB          0
`define MGR_INST_OPTION_TGT_SIZE         (`MGR_INST_OPTION_TGT_MSB - `MGR_INST_OPTION_TGT_LSB +1)
`define MGR_INST_OPTION_TGT_RANGE         `MGR_INST_OPTION_TGT_MSB : `MGR_INST_OPTION_TGT_LSB

//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_transfer_type
`define MGR_INST_OPTION_TRANSFER_TYPE_BCAST    0  
`define MGR_INST_OPTION_TRANSFER_TYPE_VECTOR   1  
`define MGR_INST_OPTION_TRANSFER_TYPE_NOP      2  

`define MGR_INST_OPTION_TRANSFER_WIDTH        2
`define MGR_INST_OPTION_TRANSFER_MSB          `MGR_INST_OPTION_TRANSFER_WIDTH-1
`define MGR_INST_OPTION_TRANSFER_LSB          0
`define MGR_INST_OPTION_TRANSFER_SIZE         (`MGR_INST_OPTION_TRANSFER_MSB - `MGR_INST_OPTION_TRANSFER_LSB +1)
`define MGR_INST_OPTION_TRANSFER_RANGE         `MGR_INST_OPTION_TRANSFER_MSB : `MGR_INST_OPTION_TRANSFER_LSB
//-------------------------------------------------------------
// - FIXME : Must match python_typedef.vh python_order_type
`define MGR_INST_OPTION_ORDER_TYPE_CWBP    0      
`define MGR_INST_OPTION_ORDER_TYPE_WCBP    1      
`define MGR_INST_OPTION_ORDER_TYPE_NOP     2      

`define MGR_INST_OPTION_ORDER_WIDTH        3
`define MGR_INST_OPTION_ORDER_MSB          `MGR_INST_OPTION_ORDER_WIDTH-1
`define MGR_INST_OPTION_ORDER_LSB          0
`define MGR_INST_OPTION_ORDER_SIZE         (`MGR_INST_OPTION_ORDER_MSB - `MGR_INST_OPTION_ORDER_LSB +1)
`define MGR_INST_OPTION_ORDER_RANGE         `MGR_INST_OPTION_ORDER_MSB : `MGR_INST_OPTION_ORDER_LSB


//---------------------------------------------------------------------------------------------------------------------
// Instruction Memory

// Each instruction takes ~10 reads
// If a network has ~1M neurons
// Each instruction is for a group of up to 32 ANs
// 1M/32 ~32000 operations
// ~500 per manager
// Instruction memory ~5000

`define MGR_INSTRUCTION_MEMORY_DEPTH   `MGR_WU_MEMORY_DEPTH 
`define MGR_INSTRUCTION_MEMORY_MSB     `MGR_INSTRUCTION_MEMORY_DEPTH-1
`define MGR_INSTRUCTION_MEMORY_LSB     0
`define MGR_INSTRUCTION_MEMORY_SIZE    (`MGR_INSTRUCTION_MEMORY_MSB - `MGR_INSTRUCTION_MEMORY_LSB +1)
`define MGR_INSTRUCTION_MEMORY_RANGE    `MGR_INSTRUCTION_MEMORY_MSB : `MGR_INSTRUCTION_MEMORY_LSB


`define MGR_INSTRUCTION_ADDRESS_WIDTH   (`CLOG2(`MGR_INSTRUCTION_MEMORY_DEPTH )) 
`define MGR_INSTRUCTION_ADDRESS_MSB     `MGR_INSTRUCTION_ADDRESS_WIDTH-1
`define MGR_INSTRUCTION_ADDRESS_LSB     0
`define MGR_INSTRUCTION_ADDRESS_SIZE    (`MGR_INSTRUCTION_ADDRESS_MSB - `MGR_INSTRUCTION_ADDRESS_LSB +1)
`define MGR_INSTRUCTION_ADDRESS_RANGE    `MGR_INSTRUCTION_ADDRESS_MSB : `MGR_INSTRUCTION_ADDRESS_LSB


`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_WIDTH    `COMMON_STD_INTF_CNTL_WIDTH 
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_WIDTH)-1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_LSB      0
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_WIDTH    `COMMON_STD_INTF_CNTL_WIDTH 
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_WIDTH)-1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_LSB      ( `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_MSB+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_WIDTH      `MGR_INST_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_WIDTH) -1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB      ( `MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_MSB+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_WIDTH      `MGR_WU_OPT_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_WIDTH) -1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB      ( `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_MSB+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_WIDTH      `MGR_WU_OPT_VALUE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_WIDTH) -1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB      ( `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_MSB+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_WIDTH      `MGR_WU_OPT_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_WIDTH) -1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB      ( `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_MSB+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_WIDTH      `MGR_WU_OPT_VALUE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_WIDTH) -1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB      ( `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_MSB+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_WIDTH      `MGR_WU_OPT_TYPE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB+`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_WIDTH) -1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_MSB)+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_SIZE     ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB) - (`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB) +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_LSB

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_WIDTH      `MGR_WU_OPT_VALUE_WIDTH
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_MSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB)+(`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_WIDTH)) -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB      ((`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_MSB)+1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_SIZE     ( `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_RANGE      `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_LSB


`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_WIDTH      `MGR_INSTRUCTION_MEMORY_AGGREGATE_ICNTL_WIDTH     \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_DCNTL_WIDTH     \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPER_WIDTH      \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE0_WIDTH \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL0_WIDTH  \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE1_WIDTH \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL1_WIDTH  \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_TYPE2_WIDTH \
                                                       +`MGR_INSTRUCTION_MEMORY_AGGREGATE_OPT_VAL2_WIDTH  

`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_MSB            `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_WIDTH -1
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_LSB            0
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_SIZE           (`MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_MSB - `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_LSB +1)
`define MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_RANGE           `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_MSB : `MGR_INSTRUCTION_MEMORY_AGGREGATE_MEM_LSB


//---------------------------------------------------------------------------------------------------------------------
// Storage Descriptor Memory

// FIXME - need to check depth equirements (for sim, keep small)
// This is per manager storage. The pointers will include additional bits for
// the manager ID

`define MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH   2048
`define MGR_LOCAL_STORAGE_DESC_MEMORY_MSB     `MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH-1
`define MGR_LOCAL_STORAGE_DESC_MEMORY_LSB     0
`define MGR_LOCAL_STORAGE_DESC_MEMORY_SIZE    (`MGR_LOCAL_STORAGE_DESC_MEMORY_MSB - `MGR_LOCAL_STORAGE_DESC_MEMORY_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_MEMORY_RANGE    `MGR_LOCAL_STORAGE_DESC_MEMORY_MSB : `MGR_LOCAL_STORAGE_DESC_MEMORY_LSB


`define MGR_LOCAL_STORAGE_DESC_ADDRESS_WIDTH   (`CLOG2(`MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH )) 
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_MSB     `MGR_LOCAL_STORAGE_DESC_ADDRESS_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_LSB     0
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_SIZE    (`MGR_LOCAL_STORAGE_DESC_ADDRESS_MSB - `MGR_LOCAL_STORAGE_DESC_ADDRESS_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_ADDRESS_RANGE    `MGR_LOCAL_STORAGE_DESC_ADDRESS_MSB : `MGR_LOCAL_STORAGE_DESC_ADDRESS_LSB




// Average number of consequtive/jump fields per storage descriptor
//`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_PER_DESC   `MGR_INST_CONS_JUMP_DEPTH / `MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH         
//

// size of consequtive and jump fields - FIXME : TBD
// Set to number of operands but may also need to be longer to accomodate number of lanes with vector 
// FIXME: update cjWidth in createReadmem.py
`define MGR_INST_CONS_JUMP_FIELD_WIDTH        `MGR_OP_MAX_NUM_OF_OPERANDS_WIDTH + (`CLOG2(`MGR_NUM_OF_EXEC_LANES))
`define MGR_INST_CONS_JUMP_FIELD_MSB          `MGR_INST_CONS_JUMP_FIELD_WIDTH-1
`define MGR_INST_CONS_JUMP_FIELD_LSB          0
`define MGR_INST_CONS_JUMP_FIELD_SIZE         (`MGR_INST_CONS_JUMP_FIELD_MSB - `MGR_INST_CONS_JUMP_FIELD_LSB +1)
`define MGR_INST_CONS_JUMP_FIELD_RANGE         `MGR_INST_CONS_JUMP_FIELD_MSB : `MGR_INST_CONS_JUMP_FIELD_LSB

// number of consequtive and jump fields - FIXME : TBD
`define MGR_INST_CONS_JUMP_DEPTH        4096
`define MGR_INST_CONS_JUMP_WIDTH        (`CLOG2(`MGR_INST_CONS_JUMP_DEPTH ))
`define MGR_INST_CONS_JUMP_MSB          `MGR_INST_CONS_JUMP_WIDTH-1
`define MGR_INST_CONS_JUMP_LSB          0
`define MGR_INST_CONS_JUMP_SIZE         (`MGR_INST_CONS_JUMP_MSB - `MGR_INST_CONS_JUMP_LSB +1)
`define MGR_INST_CONS_JUMP_RANGE         `MGR_INST_CONS_JUMP_MSB : `MGR_INST_CONS_JUMP_LSB

// This is an array wide pointer address which has the manager id pre-pended
// Note: The pointers in the instructions are array wide pointer addresses
//
`define MGR_STORAGE_DESC_ADDRESS_WIDTH         `MGR_MGR_ID_WIDTH+`MGR_LOCAL_STORAGE_DESC_ADDRESS_WIDTH               
`define MGR_STORAGE_DESC_ADDRESS_MSB           `MGR_STORAGE_DESC_ADDRESS_WIDTH-1
`define MGR_STORAGE_DESC_ADDRESS_LSB           0
`define MGR_STORAGE_DESC_ADDRESS_SIZE          (`MGR_STORAGE_DESC_ADDRESS_MSB - `MGR_STORAGE_DESC_ADDRESS_LSB +1)
`define MGR_STORAGE_DESC_ADDRESS_RANGE          `MGR_STORAGE_DESC_ADDRESS_MSB : `MGR_STORAGE_DESC_ADDRESS_LSB

`define MGR_STORAGE_DESC_MGR_ID_FIELD_MSB      `MGR_STORAGE_DESC_ADDRESS_MSB 
`define MGR_STORAGE_DESC_MGR_ID_FIELD_LSB      `MGR_STORAGE_DESC_MGR_ID_FIELD_MSB-(`MGR_MGR_ID_WIDTH-1)
`define MGR_STORAGE_DESC_MGR_ID_FIELD_RANGE    `MGR_STORAGE_DESC_MGR_ID_FIELD_MSB : `MGR_STORAGE_DESC_MGR_ID_FIELD_LSB


// Now create aggregate memories
// FIXME: Before we can use this we need to aggregate the .dat files


`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_WIDTH    `MGR_DRAM_ADDRESS_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_LSB      0
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_LSB

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_WIDTH      `MGR_INST_OPTION_ORDER_WIDTH  
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB      (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB+`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_WIDTH) -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB+1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_LSB

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_WIDTH      `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_MSB      (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB+`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_WIDTH) -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_MSB+1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_LSB


`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_WIDTH      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CJ_PTR_WIDTH    \
                                                       +`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ORDER_WIDTH     \
                                                       +`MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_WIDTH    

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_MSB            `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_WIDTH -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_LSB            0
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_SIZE           (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_RANGE           `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_MEM_LSB





//`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_DEPTH   `MGR_LOCAL_STORAGE_DESC_MEMORY_DEPTH*`MGR_LOCAL_STORAGE_DESC_CONSJUMP_PER_DESC*2   // 2 ~jump,consequtive
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_DEPTH   `MGR_INST_CONS_JUMP_DEPTH
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_MSB     `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_DEPTH-1
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_LSB     0
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_SIZE    (`MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_MSB - `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_RANGE    `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_MSB : `MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_LSB


`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_WIDTH   (`CLOG2(`MGR_LOCAL_STORAGE_DESC_CONSJUMP_MEMORY_DEPTH )) 
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_MSB     `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_LSB     0
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_SIZE    (`MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_MSB - `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_RANGE    `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_MSB : `MGR_LOCAL_STORAGE_DESC_CONSJUMP_ADDRESS_LSB


`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_WIDTH    `MGR_INST_CONS_JUMP_FIELD_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_MSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_WIDTH-1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_LSB      0
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_LSB

`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_WIDTH      `COMMON_STD_INTF_CNTL_WIDTH 
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_MSB      (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB+`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_WIDTH) -1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB      `MGR_LOCAL_STORAGE_DESC_AGGREGATE_ADDR_MSB+1
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_SIZE     (`MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_MSB - `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_RANGE     `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_MSB : `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_LSB


`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_WIDTH       `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CNTL_WIDTH     \
                                                                + `MGR_LOCAL_STORAGE_DESC_AGGREGATE_CONSJUMP_WIDTH 
                                                                

`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_MSB            `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_WIDTH -1
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_LSB            0
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_SIZE           (`MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_MSB - `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_LSB +1)
`define MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_RANGE           `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_MSB : `MGR_LOCAL_STORAGE_DESC_CONSJUMP_AGGREGATE_MEM_LSB







//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------
// DRAM Memory

`define MGR_DRAM_NUM_CHANNELS                       2
`define MGR_DRAM_NUM_BANKS                          32
`define MGR_DRAM_NUM_PAGES                          4096
`define MGR_DRAM_PAGE_SIZE                          4096
`define MGR_DRAM_NUM_WORDS_PER_PAGE                 `MGR_DRAM_PAGE_SIZE/32
`define MGR_DRAM_BURST_SIZE                         2

// Define state of signals
// CS, CMD1, CMD0
`define MGR_DRAM_COMMAND_NOP          3'b000
`define MGR_DRAM_COMMAND_PO           3'b011
`define MGR_DRAM_COMMAND_PC           3'b010
`define MGR_DRAM_COMMAND_PR           3'b001
`define MGR_DRAM_COMMAND_CR           3'b010
`define MGR_DRAM_COMMAND_CW           3'b011
`define MGR_DRAM_COMMAND_NUM_OF_OPS   6

// cache line size 
`define MGR_DRAM_NUM_CLINES_PER_PAGE             (`MGR_DRAM_PAGE_SIZE/(`MGR_DRAM_INTF_WIDTH*`MGR_DRAM_BURST_SIZE))    // CLINE is the DRAM burst size
`define MGR_DRAM_CLINE_SIZE                      (`MGR_DRAM_PAGE_SIZE/`MGR_DRAM_NUM_CLINES_PER_PAGE              )
`define MGR_DRAM_NUM_LINES_PER_CLINE             (`MGR_DRAM_CLINE_SIZE/`MGR_MMC_TO_MRC_INTF_WIDTH                )    // Line is the transaction size from the MMC
`define MGR_DRAM_NUM_LINES_PER_REQUEST           (`MGR_DRAM_NUM_LINES_PER_CLINE                                  )    // MMC transactions per memory request
`define MGR_DRAM_NUM_WORDS_PER_CLINE             (`MGR_DRAM_NUM_WORDS_PER_PAGE/`MGR_DRAM_NUM_CLINES_PER_PAGE     )
`define MGR_DRAM_NUM_LINES_PER_PAGE              (`MGR_DRAM_NUM_CLINES_PER_PAGE * `MGR_DRAM_NUM_LINES_PER_CLINE  )
`define MGR_DRAM_NUM_WORDS_PER_LINE              (`MGR_DRAM_NUM_WORDS_PER_PAGE/`MGR_DRAM_NUM_LINES_PER_PAGE      )

//****************************************************************************************************
//****************************************************************************************************
// Manually set based on 

`define MGR_DRAM_REQUEST_CLINE_LT_PAGE
`undef  MGR_DRAM_REQUEST_CLINE_LT_PAGE

`undef  MGR_DRAM_REQUEST_LINE_LT_CACHELINE
`define MGR_DRAM_REQUEST_LINE_LT_CACHELINE

//****************************************************************************************************
//****************************************************************************************************
  

`define MGR_DRAM_PHY_ADDRESS_WIDTH               `MGR_DRAM_PAGE_ADDRESS_WIDTH 
`define MGR_DRAM_PHY_ADDRESS_MSB                 `MGR_DRAM_PHY_ADDRESS_WIDTH-1
`define MGR_DRAM_PHY_ADDRESS_LSB                  0
`define MGR_DRAM_PHY_ADDRESS_SIZE                (`MGR_DRAM_PHY_ADDRESS_MSB - `MGR_DRAM_PHY_ADDRESS_LSB +1)
`define MGR_DRAM_PHY_ADDRESS_RANGE                `MGR_DRAM_PHY_ADDRESS_MSB : `MGR_DRAM_PHY_ADDRESS_LSB

`define MGR_DRAM_INTF_WIDTH                          2048
`define MGR_DRAM_INTF_MSB                         `MGR_DRAM_INTF_WIDTH-1
`define MGR_DRAM_INTF_LSB                         0
`define MGR_DRAM_INTF_SIZE                        (`MGR_DRAM_INTF_MSB - `MGR_DRAM_INTF_LSB +1)
`define MGR_DRAM_INTF_RANGE                        `MGR_DRAM_INTF_MSB : `MGR_DRAM_INTF_LSB

`define MGR_DRAM_INTF_MASK_WIDTH                       `MGR_DRAM_INTF_WIDTH/`MGR_EXEC_LANE_WIDTH               
`define MGR_DRAM_INTF_MASK_MSB                         `MGR_DRAM_INTF_MASK_WIDTH-1
`define MGR_DRAM_INTF_MASK_LSB                         0
`define MGR_DRAM_INTF_MASK_SIZE                        (`MGR_DRAM_INTF_MASK_MSB - `MGR_DRAM_INTF_MASK_LSB +1)
`define MGR_DRAM_INTF_MASK_RANGE                        `MGR_DRAM_INTF_MASK_MSB : `MGR_DRAM_INTF_MASK_LSB

`define MGR_DRAM_INTF_BITS_PER_CLOCK_GROUP          32
`define MGR_DRAM_BUS_NUM_CLK_GROUPS                 `MGR_DRAM_INTF_WIDTH / `MGR_DRAM_INTF_BITS_PER_CLOCK_GROUP
`define MGR_DRAM_CLK_GROUP_WIDTH                    `MGR_DRAM_BUS_NUM_CLK_GROUPS 
`define MGR_DRAM_CLK_GROUP_MSB                      `MGR_DRAM_CLK_GROUP_WIDTH-1
`define MGR_DRAM_CLK_GROUP_LSB                      0
`define MGR_DRAM_CLK_GROUP_SIZE                     (`MGR_DRAM_CLK_GROUP_MSB - `MGR_DRAM_CLK_GROUP_LSB +1)
`define MGR_DRAM_CLK_GROUP_RANGE                    `MGR_DRAM_CLK_GROUP_MSB : `MGR_DRAM_CLK_GROUP_LSB



`define MGR_DRAM_NUM_CHANNELS_VECTOR_WIDTH                       `MGR_DRAM_NUM_CHANNELS
`define MGR_DRAM_NUM_CHANNELS_VECTOR_MSB                         `MGR_DRAM_NUM_CHANNELS_VECTOR_WIDTH-1
`define MGR_DRAM_NUM_CHANNELS_VECTOR_LSB                         0
`define MGR_DRAM_NUM_CHANNELS_VECTOR_SIZE                        (`MGR_DRAM_NUM_CHANNELS_VECTOR_MSB - `MGR_DRAM_NUM_CHANNELS_VECTOR_LSB +1)
`define MGR_DRAM_NUM_CHANNELS_VECTOR_RANGE                        `MGR_DRAM_NUM_CHANNELS_VECTOR_MSB : `MGR_DRAM_NUM_CHANNELS_VECTOR_LSB

`define MGR_DRAM_NUM_BANKS_VECTOR_WIDTH                       `MGR_DRAM_NUM_BANKS
`define MGR_DRAM_NUM_BANKS_VECTOR_MSB                         `MGR_DRAM_NUM_BANKS_VECTOR_WIDTH-1
`define MGR_DRAM_NUM_BANKS_VECTOR_LSB                         0
`define MGR_DRAM_NUM_BANKS_VECTOR_SIZE                        (`MGR_DRAM_NUM_BANKS_VECTOR_MSB - `MGR_DRAM_NUM_BANKS_VECTOR_LSB +1)
`define MGR_DRAM_NUM_BANKS_VECTOR_RANGE                        `MGR_DRAM_NUM_BANKS_VECTOR_MSB : `MGR_DRAM_NUM_BANKS_VECTOR_LSB


`define MGR_DRAM_PHY_BURST_WIDTH                      (`CLOG2(`MGR_DRAM_BURST_SIZE ))
`define MGR_DRAM_PHY_BURST_MSB                         `MGR_DRAM_PHY_BURST_WIDTH-1
`define MGR_DRAM_PHY_BURST_LSB                         0
`define MGR_DRAM_PHY_BURST_SIZE                        (`MGR_DRAM_PHY_BURST_MSB - `MGR_DRAM_PHY_BURST_LSB +1)
`define MGR_DRAM_PHY_BURST_RANGE                        `MGR_DRAM_PHY_BURST_MSB : `MGR_DRAM_PHY_BURST_LSB

//---------------------------------------------------------------------------------------------------------------------
// MMC to MRC

`define MGR_MMC_TO_MRC_INTF_WIDTH                       `MGR_DRAM_INTF_WIDTH
`define MGR_MMC_TO_MRC_INTF_MSB                         `MGR_MMC_TO_MRC_INTF_WIDTH-1
`define MGR_MMC_TO_MRC_INTF_LSB                         0
`define MGR_MMC_TO_MRC_INTF_SIZE                        (`MGR_MMC_TO_MRC_INTF_MSB - `MGR_MMC_TO_MRC_INTF_LSB +1)
`define MGR_MMC_TO_MRC_INTF_RANGE                        `MGR_MMC_TO_MRC_INTF_MSB : `MGR_MMC_TO_MRC_INTF_LSB

`define MGR_MMC_TO_MRC_INTF_NUM_WORDS          `MGR_MMC_TO_MRC_INTF_WIDTH/32

`define MGR_MMC_TO_MRC_INTF_NUM_WORDS_WIDTH                       `MGR_MMC_TO_MRC_INTF_NUM_WORDS          
`define MGR_MMC_TO_MRC_INTF_NUM_WORDS_MSB                         `MGR_MMC_TO_MRC_INTF_NUM_WORDS_WIDTH-1
`define MGR_MMC_TO_MRC_INTF_NUM_WORDS_LSB                         0
`define MGR_MMC_TO_MRC_INTF_NUM_WORDS_SIZE                        (`MGR_MMC_TO_MRC_INTF_NUM_WORDS_MSB - `MGR_MMC_TO_MRC_INTF_NUM_WORDS_LSB +1)
`define MGR_MMC_TO_MRC_INTF_NUM_WORDS_RANGE                        `MGR_MMC_TO_MRC_INTF_NUM_WORDS_MSB : `MGR_MMC_TO_MRC_INTF_NUM_WORDS_LSB

`define MGR_MMC_TO_MRC_WORD_ADDRESS_WIDTH                       (`CLOG2(`MGR_MMC_TO_MRC_INTF_NUM_WORDS ))
`define MGR_MMC_TO_MRC_WORD_ADDRESS_MSB                         `MGR_MMC_TO_MRC_WORD_ADDRESS_WIDTH-1
`define MGR_MMC_TO_MRC_WORD_ADDRESS_LSB                         0
`define MGR_MMC_TO_MRC_WORD_ADDRESS_SIZE                        (`MGR_MMC_TO_MRC_WORD_ADDRESS_MSB - `MGR_MMC_TO_MRC_WORD_ADDRESS_LSB +1)
`define MGR_MMC_TO_MRC_WORD_ADDRESS_RANGE                        `MGR_MMC_TO_MRC_WORD_ADDRESS_MSB : `MGR_MMC_TO_MRC_WORD_ADDRESS_LSB

//------------------------------------------------------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------------------------------------------------------
// HOW MANY BITS TO ADDRESS A 64Gb MEMORY WITH 64 PORTS
//  - use byte address
//  - need to address 8GB
//  pow(2,33) = 8589934592 ~ 8G
//  we need 33 bits to address 8G e.g. 2^32 ~ 4G, + 2^31 ~ 2G + ....... + 2^0 ~ 1  ~= 8G
//  = 1

`define MGR_DRAM_CHANNEL_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_CHANNELS ))
`define MGR_DRAM_CHANNEL_ADDRESS_MSB                         `MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_CHANNEL_ADDRESS_LSB                         0
`define MGR_DRAM_CHANNEL_ADDRESS_SIZE                        (`MGR_DRAM_CHANNEL_ADDRESS_MSB - `MGR_DRAM_CHANNEL_ADDRESS_LSB +1)
`define MGR_DRAM_CHANNEL_ADDRESS_RANGE                        `MGR_DRAM_CHANNEL_ADDRESS_MSB : `MGR_DRAM_CHANNEL_ADDRESS_LSB

`define MGR_DRAM_BANK_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_BANKS ))
`define MGR_DRAM_BANK_ADDRESS_MSB                         `MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_BANK_ADDRESS_LSB                         0
`define MGR_DRAM_BANK_ADDRESS_SIZE                        (`MGR_DRAM_BANK_ADDRESS_MSB - `MGR_DRAM_BANK_ADDRESS_LSB +1)
`define MGR_DRAM_BANK_ADDRESS_RANGE                        `MGR_DRAM_BANK_ADDRESS_MSB : `MGR_DRAM_BANK_ADDRESS_LSB

`define MGR_DRAM_PAGE_ADDRESS_WIDTH                      (`CLOG2(`MGR_DRAM_NUM_PAGES ))
`define MGR_DRAM_PAGE_ADDRESS_MSB                         `MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_PAGE_ADDRESS_LSB                         0
`define MGR_DRAM_PAGE_ADDRESS_SIZE                        (`MGR_DRAM_PAGE_ADDRESS_MSB - `MGR_DRAM_PAGE_ADDRESS_LSB +1)
`define MGR_DRAM_PAGE_ADDRESS_RANGE                        `MGR_DRAM_PAGE_ADDRESS_MSB : `MGR_DRAM_PAGE_ADDRESS_LSB

`define MGR_DRAM_WORD_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_WORDS_PER_PAGE ))
`define MGR_DRAM_WORD_ADDRESS_MSB                         `MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_WORD_ADDRESS_LSB                         0
`define MGR_DRAM_WORD_ADDRESS_SIZE                        (`MGR_DRAM_WORD_ADDRESS_MSB - `MGR_DRAM_WORD_ADDRESS_LSB +1)
`define MGR_DRAM_WORD_ADDRESS_RANGE                        `MGR_DRAM_WORD_ADDRESS_MSB : `MGR_DRAM_WORD_ADDRESS_LSB

// We need to make a distinction between a LINE and a CACHELINE
// A line is a single transaction/cycle of data from the MMC. Currently, in our case the interface is 2048 bits so a line is 32 words
// A cacheline is the amount of data the DRAM provides during a read (or needs during a write). The DRAM interface is 2048 bits with a burst of
// 2, so the DRAM provides 4096 bits per cacheline (which the the baeline DRAM is a page)
//
// If the interface from the MMC were to be 4096 bits, a line and cachline would be the same
// When we parse memory descriptors, we are looking for line transitions, not cacheline transitions.
// However, when we need to remember each request will actually provide two lines
//
// We access a cache line for each read. We need to know which line is being accessed for the given word address in the page
`define MGR_DRAM_LINE_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_LINES_PER_CLINE))
`define MGR_DRAM_LINE_ADDRESS_MSB                         `MGR_DRAM_LINE_ADDRESS_WIDTH-1
`define MGR_DRAM_LINE_ADDRESS_LSB                         0
`define MGR_DRAM_LINE_ADDRESS_SIZE                        (`MGR_DRAM_LINE_ADDRESS_MSB - `MGR_DRAM_LINE_ADDRESS_LSB +1)
`define MGR_DRAM_LINE_ADDRESS_RANGE                        `MGR_DRAM_LINE_ADDRESS_MSB : `MGR_DRAM_LINE_ADDRESS_LSB

`define MGR_DRAM_LINE_IN_WORD_ADDRESS_RANGE                    `MGR_DRAM_WORD_ADDRESS_MSB : (`MGR_DRAM_WORD_ADDRESS_MSB-(`MGR_DRAM_LINE_ADDRESS_WIDTH-1))
`define MGR_DRAM_WORD_WO_LINE_ADDRESS_RANGE                    (`MGR_DRAM_WORD_ADDRESS_MSB-`MGR_DRAM_LINE_ADDRESS_WIDTH):0

`ifdef  MGR_DRAM_REQUEST_CLINE_LT_PAGE
  // We access a cache line for each read. We need to know which line is being accessed for the given word address in the page
  `define MGR_DRAM_CLINE_ADDRESS_WIDTH                       (`CLOG2(`MGR_DRAM_NUM_CLINES_PER_PAGE
  `define MGR_DRAM_CLINE_ADDRESS_MSB                         `MGR_DRAM_CLINE_ADDRESS_WIDTH-1
  `define MGR_DRAM_CLINE_ADDRESS_LSB                         0
  `define MGR_DRAM_CLINE_ADDRESS_SIZE                        (`MGR_DRAM_CLINE_ADDRESS_MSB - `MGR_DRAM_CLINE_ADDRESS_LSB +1)
  `define MGR_DRAM_CLINE_ADDRESS_RANGE                        `MGR_DRAM_CLINE_ADDRESS_MSB : `MGR_DRAM_CLINE_ADDRESS_LSB
  
  `define MGR_DRAM_CLINE_IN_WORD_ADDRESS_RANGE                    `MGR_DRAM_WORD_ADDRESS_MSB : (`MGR_DRAM_WORD_ADDRESS_MSB-(`MGR_DRAM_CLINE_ADDRESS_WIDTH-1))
  `define MGR_DRAM_WORD_WO_CLINE_ADDRESS_RANGE                    (`MGR_DRAM_WORD_ADDRESS_MSB-`MGR_DRAM_CLINE_ADDRESS_WIDTH):0
`endif



// DRAM has 64 interface, 2 channels,  32 banks, 4096 pages and 4096 bits per page
`define MGR_DRAM_ADDRESS_WIDTH             `MGR_MGR_ID_WIDTH+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH+`MGR_DRAM_BANK_ADDRESS_WIDTH+`MGR_DRAM_PAGE_ADDRESS_WIDTH+`MGR_DRAM_WORD_ADDRESS_WIDTH+2  // byte address
`define MGR_DRAM_ADDRESS_MSB               `MGR_DRAM_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_LSB               0
`define MGR_DRAM_ADDRESS_SIZE              (`MGR_DRAM_ADDRESS_MSB - `MGR_DRAM_ADDRESS_LSB +1)
`define MGR_DRAM_ADDRESS_RANGE              `MGR_DRAM_ADDRESS_MSB : `MGR_DRAM_ADDRESS_LSB

// DRAM local address width (doesnt include manager ID
`define MGR_DRAM_LOCAL_ADDRESS_WIDTH             `MGR_DRAM_CHANNEL_ADDRESS_WIDTH+`MGR_DRAM_BANK_ADDRESS_WIDTH+`MGR_DRAM_PAGE_ADDRESS_WIDTH+`MGR_DRAM_WORD_ADDRESS_WIDTH+2  // byte address
`define MGR_DRAM_LOCAL_ADDRESS_MSB               `MGR_DRAM_LOCAL_ADDRESS_WIDTH-1
`define MGR_DRAM_LOCAL_ADDRESS_LSB               0
`define MGR_DRAM_LOCAL_ADDRESS_SIZE              (`MGR_DRAM_LOCAL_ADDRESS_MSB - `MGR_DRAM_LOCAL_ADDRESS_LSB +1)
`define MGR_DRAM_LOCAL_ADDRESS_RANGE              `MGR_DRAM_LOCAL_ADDRESS_MSB : `MGR_DRAM_LOCAL_ADDRESS_LSB

// generate ranges so we can extract the fields from a given address
`define MGR_DRAM_ADDRESS_WORD_FIELD_LSB                         2  // account for byte address
`define MGR_DRAM_ADDRESS_WORD_FIELD_MSB                         `MGR_DRAM_ADDRESS_WORD_FIELD_LSB+`MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_WORD_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_WORD_FIELD_MSB - `MGR_DRAM_ADDRESS_WORD_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_WORD_FIELD_RANGE                        `MGR_DRAM_ADDRESS_WORD_FIELD_MSB : `MGR_DRAM_ADDRESS_WORD_FIELD_LSB

`ifdef MGR_DRAM_REQUEST_CLINE_LT_PAGE
  `define MGR_DRAM_ADDRESS_CLINE_FIELD_MSB                         `MGR_DRAM_ADDRESS_WORD_FIELD_MSB
  `define MGR_DRAM_ADDRESS_CLINE_FIELD_LSB                         (`MGR_DRAM_ADDRESS_CLINE_FIELD_MSB-`MGR_DRAM_CLINE_ADDRESS_WIDTH)+1
  `define MGR_DRAM_ADDRESS_CLINE_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_CLINE_FIELD_MSB - `MGR_DRAM_ADDRESS_CLINE_FIELD_LSB +1)
  `define MGR_DRAM_ADDRESS_CLINE_FIELD_RANGE                        `MGR_DRAM_ADDRESS_CLINE_FIELD_MSB : `MGR_DRAM_ADDRESS_CLINE_FIELD_LSB
`endif

`ifdef  MGR_DRAM_REQUEST_LINE_LT_CACHELINE
  `define MGR_DRAM_ADDRESS_LINE_FIELD_MSB                         `MGR_DRAM_ADDRESS_WORD_FIELD_MSB
  `define MGR_DRAM_ADDRESS_LINE_FIELD_LSB                         (`MGR_DRAM_ADDRESS_LINE_FIELD_MSB-`MGR_DRAM_LINE_ADDRESS_WIDTH)+1
  `define MGR_DRAM_ADDRESS_LINE_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_LINE_FIELD_MSB - `MGR_DRAM_ADDRESS_LINE_FIELD_LSB +1)
  `define MGR_DRAM_ADDRESS_LINE_FIELD_RANGE                        `MGR_DRAM_ADDRESS_LINE_FIELD_MSB : `MGR_DRAM_ADDRESS_LINE_FIELD_LSB
`endif

`define MGR_DRAM_ADDRESS_PAGE_FIELD_LSB                         `MGR_DRAM_ADDRESS_WORD_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_PAGE_FIELD_MSB                         `MGR_DRAM_ADDRESS_PAGE_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_PAGE_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_PAGE_FIELD_MSB - `MGR_DRAM_ADDRESS_PAGE_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_PAGE_FIELD_RANGE                        `MGR_DRAM_ADDRESS_PAGE_FIELD_MSB : `MGR_DRAM_ADDRESS_PAGE_FIELD_LSB

`define MGR_DRAM_ADDRESS_BANK_FIELD_LSB                         `MGR_DRAM_ADDRESS_PAGE_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_BANK_FIELD_MSB                         `MGR_DRAM_ADDRESS_BANK_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_BANK_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_BANK_FIELD_MSB - `MGR_DRAM_ADDRESS_BANK_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_BANK_FIELD_RANGE                        `MGR_DRAM_ADDRESS_BANK_FIELD_MSB : `MGR_DRAM_ADDRESS_BANK_FIELD_LSB

`define MGR_DRAM_ADDRESS_CHAN_FIELD_LSB                         `MGR_DRAM_ADDRESS_BANK_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_CHAN_FIELD_MSB                         `MGR_DRAM_ADDRESS_CHAN_FIELD_LSB+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_ADDRESS_CHAN_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_CHAN_FIELD_MSB - `MGR_DRAM_ADDRESS_CHAN_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_CHAN_FIELD_RANGE                        `MGR_DRAM_ADDRESS_CHAN_FIELD_MSB : `MGR_DRAM_ADDRESS_CHAN_FIELD_LSB

`define MGR_DRAM_ADDRESS_MGR_FIELD_LSB                         `MGR_DRAM_ADDRESS_CHAN_FIELD_MSB+1
`define MGR_DRAM_ADDRESS_MGR_FIELD_MSB                         `MGR_DRAM_ADDRESS_MGR_FIELD_LSB+`MGR_MGR_ID_WIDTH-1
`define MGR_DRAM_ADDRESS_MGR_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_MGR_FIELD_MSB - `MGR_DRAM_ADDRESS_MGR_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_MGR_FIELD_RANGE                        `MGR_DRAM_ADDRESS_MGR_FIELD_MSB : `MGR_DRAM_ADDRESS_MGR_FIELD_LSB

// Useful macros
// extract bank without lsb (for PBC increment in request generation
`define MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_LSB                         `MGR_DRAM_ADDRESS_BANK_FIELD_LSB+1
`define MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_MSB                         `MGR_DRAM_ADDRESS_BANK_FIELD_MSB
`define MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_SIZE                        (`MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_MSB - `MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_LSB +1)
`define MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_RANGE                        `MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_MSB : `MGR_DRAM_ADDRESS_BANK_DIV2_FIELD_LSB



// Field locations based on address formed from access order
// WCBP
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB                         2  // account for byte address
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB+`MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_WORD_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_WORD_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB                         `MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_CHAN_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_LSB                         (`MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB-`MGR_DRAM_LINE_ADDRESS_WIDTH)+1
`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_WORD_FIELD_MSB
`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_LINE_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_LINE_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_LINE_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_LINE_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB                         `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_BANK_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_BANK_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB                         `MGR_DRAM_WCBP_ORDER_BANK_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_MSB                         `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_SIZE                        (`MGR_DRAM_WCBP_ORDER_PAGE_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_PAGE_FIELD_RANGE                        `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_PAGE_FIELD_LSB

// When we increment through addresses when determining memory requests or streaming data, we actually increment bank x2
// SO the address is formed by dropping the bank LSB. SO we need indexes for those cases when the bank lsb is not included in the address
`define MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB             `MGR_DRAM_WCBP_ORDER_CHAN_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB             `MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-2
`define MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_SIZE            (`MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_RANGE            `MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB

`define MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB             `MGR_DRAM_WCBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB+1
`define MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_MSB             `MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_SIZE            (`MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_MSB - `MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB +1)
`define MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_RANGE            `MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_MSB : `MGR_DRAM_WCBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB


// CWBP
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB                         2  // account for byte address
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB+`MGR_DRAM_CHANNEL_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_CHAN_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_LSB

`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_CHAN_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB+`MGR_DRAM_WORD_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_WORD_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_WORD_FIELD_LSB

`ifdef  MGR_DRAM_REQUEST_LINE_LT_CACHELINE
  `define MGR_DRAM_CWBP_ORDER_LINE_FIELD_LSB                         (`MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB-`MGR_DRAM_LINE_ADDRESS_WIDTH)+1
  `define MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB
  `define MGR_DRAM_CWBP_ORDER_LINE_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_LINE_FIELD_LSB +1)
  `define MGR_DRAM_CWBP_ORDER_LINE_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_LINE_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_LINE_FIELD_LSB
`endif

`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_BANK_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_BANK_FIELD_LSB

`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_BANK_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_PAGE_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_PAGE_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_PAGE_FIELD_LSB

// When we increment through addresses when determining memory requests or streaming data, we actually increment bank x2
// SO the address is formed by dropping the bank LSB. SO we need indexes for those cases when the bank lsb is not included in the address
`define MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_WORD_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB+`MGR_DRAM_BANK_ADDRESS_WIDTH-2
`define MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_LSB

`define MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB                         `MGR_DRAM_CWBP_ORDER_BANK_WO_BANK_LSB_FIELD_MSB+1
`define MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_MSB                         `MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB+`MGR_DRAM_PAGE_ADDRESS_WIDTH-1
`define MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_SIZE                        (`MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_MSB - `MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB +1)
`define MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_RANGE                        `MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_MSB : `MGR_DRAM_CWBP_ORDER_PAGE_WO_BANK_LSB_FIELD_LSB

//------------------------------------------------------------------------------------------------------------------------
// The memory requestor will always open the next channel/bank/page based on the current address
// If a memory request provides an entire page, then to determine whether we
// need a request, just form an adrress based on page/bank/channel and increment 
// If a memory request is a partial page (line), then form an address based on PBLC or PBCL
//
// 1) Line same size as page, so only increment page/bank/channel
`ifndef  MGR_DRAM_REQUEST_CLINE_LT_PAGE
  // PBC
  `define MGR_DRAM_PBC_CHAN_FIELD_WIDTH       `MGR_DRAM_CHANNEL_ADDRESS_WIDTH
  `define MGR_DRAM_PBC_CHAN_FIELD_LSB         0
  `define MGR_DRAM_PBC_CHAN_FIELD_MSB         `MGR_DRAM_PBC_CHAN_FIELD_LSB+`MGR_DRAM_PBC_CHAN_FIELD_WIDTH -1
  `define MGR_DRAM_PBC_CHAN_FIELD_SIZE        (`MGR_DRAM_PBC_CHAN_FIELD_MSB - `MGR_DRAM_PBC_CHAN_FIELD_LSB +1)
  `define MGR_DRAM_PBC_CHAN_FIELD_RANGE        `MGR_DRAM_PBC_CHAN_FIELD_MSB : `MGR_DRAM_PBC_CHAN_FIELD_LSB
  
  // Remember, we increment bank/2, so reduce width by 1
  `define MGR_DRAM_PBC_BANK_FIELD_WIDTH       `MGR_DRAM_BANK_ADDRESS_WIDTH-1
  `define MGR_DRAM_PBC_BANK_FIELD_LSB         `MGR_DRAM_PBC_CHAN_FIELD_MSB+1
  `define MGR_DRAM_PBC_BANK_FIELD_MSB         `MGR_DRAM_PBC_BANK_FIELD_LSB+`MGR_DRAM_PBC_BANK_FIELD_WIDTH -1
  `define MGR_DRAM_PBC_BANK_FIELD_SIZE        (`MGR_DRAM_PBC_BANK_FIELD_MSB - `MGR_DRAM_PBC_BANK_FIELD_LSB +1)
  `define MGR_DRAM_PBC_BANK_FIELD_RANGE        `MGR_DRAM_PBC_BANK_FIELD_MSB : `MGR_DRAM_PBC_BANK_FIELD_LSB
  
  `define MGR_DRAM_PBC_PAGE_FIELD_WIDTH       `MGR_DRAM_PAGE_ADDRESS_WIDTH
  `define MGR_DRAM_PBC_PAGE_FIELD_LSB         `MGR_DRAM_PBC_BANK_FIELD_MSB+1
  `define MGR_DRAM_PBC_PAGE_FIELD_MSB         `MGR_DRAM_PBC_PAGE_FIELD_LSB+`MGR_DRAM_PBC_PAGE_FIELD_WIDTH -1
  `define MGR_DRAM_PBC_PAGE_FIELD_SIZE        (`MGR_DRAM_PBC_PAGE_FIELD_MSB - `MGR_DRAM_PBC_PAGE_FIELD_LSB +1)
  `define MGR_DRAM_PBC_PAGE_FIELD_RANGE        `MGR_DRAM_PBC_PAGE_FIELD_MSB : `MGR_DRAM_PBC_PAGE_FIELD_LSB
  
  `define MGR_DRAM_PBC_WIDTH                   `MGR_DRAM_PBC_PAGE_FIELD_WIDTH      \
                                              +`MGR_DRAM_PBC_BANK_FIELD_WIDTH      \
                                              +`MGR_DRAM_PBC_CHAN_FIELD_WIDTH 
                                              
  `define MGR_DRAM_PBC_MSB            `MGR_DRAM_PBC_WIDTH -1
  `define MGR_DRAM_PBC_LSB            0
  `define MGR_DRAM_PBC_SIZE           (`MGR_DRAM_PBC_MSB - `MGR_DRAM_PBC_LSB +1)
  `define MGR_DRAM_PBC_RANGE           `MGR_DRAM_PBC_MSB : `MGR_DRAM_PBC_LSB
`endif
//------------------------------------------------------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------------------------------------------------------
// Other useful macros

`define MGR_DRAM_BANK_DIV2_ADDRESS_WIDTH                       `MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_BANK_DIV2_ADDRESS_MSB                         `MGR_DRAM_BANK_DIV2_ADDRESS_WIDTH-1
`define MGR_DRAM_BANK_DIV2_ADDRESS_LSB                         0
`define MGR_DRAM_BANK_DIV2_ADDRESS_SIZE                        (`MGR_DRAM_BANK_DIV2_ADDRESS_MSB - `MGR_DRAM_BANK_DIV2_ADDRESS_LSB +1)
`define MGR_DRAM_BANK_DIV2_ADDRESS_RANGE                        `MGR_DRAM_BANK_DIV2_ADDRESS_MSB : `MGR_DRAM_BANK_DIV2_ADDRESS_LSB

// we always increment the bank by two, so when we load the counter which increments through the consequtive and jump fields, we will
// actually load the bank field with the bank_address[msb:1] rather than bank_address[lsb:0].
// Then we will insert the lsb into the request bank
`define MGR_DRAM_BANK_ADDRESS_WO_LSB_WIDTH                       `MGR_DRAM_BANK_ADDRESS_WIDTH-1
`define MGR_DRAM_BANK_ADDRESS_WO_LSB_MSB                         `MGR_DRAM_BANK_ADDRESS_MSB
`define MGR_DRAM_BANK_ADDRESS_WO_LSB_LSB                         `MGR_DRAM_BANK_ADDRESS_LSB+1
`define MGR_DRAM_BANK_ADDRESS_WO_LSB_SIZE                        (`MGR_DRAM_BANK_ADDRESS_WO_LSB_MSB - `MGR_DRAM_BANK_ADDRESS_WO_LSB_LSB +1)
`define MGR_DRAM_BANK_ADDRESS_WO_LSB_RANGE                        `MGR_DRAM_BANK_ADDRESS_WO_LSB_MSB : `MGR_DRAM_BANK_ADDRESS_WO_LSB_LSB

//------------------------------------------------------------------------------------------------------------------------------------------------------
//------------------------------------------------------------------------------------------------------------------------------------------------------

// 2) Line smaller than page, so increment either page/bank/channel/line or page/bank/line/channel
`ifdef  MGR_DRAM_REQUEST_CLINE_LT_PAGE

  //----------------------------------------------------------------------------------------------------
  // PBCL
  `define MGR_DRAM_PBCL_CLINE_FIELD_WIDTH       `MGR_DRAM_LINE_ADDRESS_WIDTH 
  `define MGR_DRAM_PBCL_CLINE_FIELD_LSB         0
  `define MGR_DRAM_PBCL_CLINE_FIELD_MSB         `MGR_DRAM_PBCL_CLINE_FIELD_LSB+`MGR_DRAM_PBCL_CLINE_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_CLINE_FIELD_SIZE        (`MGR_DRAM_PBCL_CLINE_FIELD_MSB - `MGR_DRAM_PBCL_CLINE_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_CLINE_FIELD_RANGE        `MGR_DRAM_PBCL_CLINE_FIELD_MSB : `MGR_DRAM_PBCL_CLINE_FIELD_LSB

  `define MGR_DRAM_PBCL_CHAN_FIELD_WIDTH       `MGR_DRAM_CHANNEL_ADDRESS_WIDTH
  `define MGR_DRAM_PBCL_CHAN_FIELD_LSB         `MGR_DRAM_PBCL_CLINE_FIELD_MSB+1
  `define MGR_DRAM_PBCL_CHAN_FIELD_MSB         `MGR_DRAM_PBCL_CHAN_FIELD_LSB+`MGR_DRAM_PBCL_CHAN_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_CHAN_FIELD_SIZE        (`MGR_DRAM_PBCL_CHAN_FIELD_MSB - `MGR_DRAM_PBCL_CHAN_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_CHAN_FIELD_RANGE        `MGR_DRAM_PBCL_CHAN_FIELD_MSB : `MGR_DRAM_PBCL_CHAN_FIELD_LSB
  
  // Remember, we increment bank/2, so reduce width by 1
  `define MGR_DRAM_PBCL_BANK_FIELD_WIDTH       `MGR_DRAM_BANK_ADDRESS_WIDTH-1
  `define MGR_DRAM_PBCL_BANK_FIELD_LSB         `MGR_DRAM_PBCL_CHAN_FIELD_MSB+1
  `define MGR_DRAM_PBCL_BANK_FIELD_MSB         `MGR_DRAM_PBCL_BANK_FIELD_LSB+`MGR_DRAM_PBCL_BANK_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_BANK_FIELD_SIZE        (`MGR_DRAM_PBCL_BANK_FIELD_MSB - `MGR_DRAM_PBCL_BANK_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_BANK_FIELD_RANGE        `MGR_DRAM_PBCL_BANK_FIELD_MSB : `MGR_DRAM_PBCL_BANK_FIELD_LSB
  
  `define MGR_DRAM_PBCL_PAGE_FIELD_WIDTH       `MGR_DRAM_PAGE_ADDRESS_WIDTH
  `define MGR_DRAM_PBCL_PAGE_FIELD_LSB         `MGR_DRAM_PBCL_BANK_FIELD_MSB+1
  `define MGR_DRAM_PBCL_PAGE_FIELD_MSB         `MGR_DRAM_PBCL_PAGE_FIELD_LSB+`MGR_DRAM_PBCL_PAGE_FIELD_WIDTH -1
  `define MGR_DRAM_PBCL_PAGE_FIELD_SIZE        (`MGR_DRAM_PBCL_PAGE_FIELD_MSB - `MGR_DRAM_PBCL_PAGE_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_PAGE_FIELD_RANGE        `MGR_DRAM_PBCL_PAGE_FIELD_MSB : `MGR_DRAM_PBCL_PAGE_FIELD_LSB
  
  `define MGR_DRAM_PBCL_WIDTH                   `MGR_DRAM_PBCL_PAGE_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBCL_BANK_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBCL_CHAN_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBCL_CLINE_FIELD_WIDTH       
  
  
  `define MGR_DRAM_PBCL_MSB            `MGR_DRAM_PBCL_WIDTH -1
  `define MGR_DRAM_PBCL_LSB            0
  `define MGR_DRAM_PBCL_SIZE           (`MGR_DRAM_PBCL_MSB - `MGR_DRAM_PBCL_LSB +1)
  `define MGR_DRAM_PBCL_RANGE           `MGR_DRAM_PBCL_MSB : `MGR_DRAM_PBCL_LSB


  // Other useful macros
  `define MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_LSB         `MGR_DRAM_PBCL_BANK_FIELD_LSB
  `define MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_MSB         `MGR_DRAM_PBCL_BANK_FIELD_MSB-1
  `define MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_SIZE        (`MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_MSB - `MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_LSB +1)
  `define MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_RANGE        `MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_MSB : `MGR_DRAM_PBCL_BANK_WO_MSB_FIELD_LSB

  //----------------------------------------------------------------------------------------------------
  // PBLC
  `define MGR_DRAM_PBLC_CHAN_FIELD_WIDTH       `MGR_DRAM_CHANNEL_ADDRESS_WIDTH
  `define MGR_DRAM_PBLC_CHAN_FIELD_LSB         0
  `define MGR_DRAM_PBLC_CHAN_FIELD_MSB         `MGR_DRAM_PBLC_CHAN_FIELD_LSB+`MGR_DRAM_PBLC_CHAN_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_CHAN_FIELD_SIZE        (`MGR_DRAM_PBLC_CHAN_FIELD_MSB - `MGR_DRAM_PBLC_CHAN_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_CHAN_FIELD_RANGE        `MGR_DRAM_PBLC_CHAN_FIELD_MSB : `MGR_DRAM_PBLC_CHAN_FIELD_LSB
  
  `define MGR_DRAM_PBLC_CLINE_FIELD_WIDTH       `MGR_DRAM_LINE_ADDRESS_WIDTH 
  `define MGR_DRAM_PBLC_CLINE_FIELD_LSB         `MGR_DRAM_PBLC_CHAN_FIELD_MSB+1
  `define MGR_DRAM_PBLC_CLINE_FIELD_MSB         `MGR_DRAM_PBLC_CLINE_FIELD_LSB+`MGR_DRAM_PBLC_CLINE_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_CLINE_FIELD_SIZE        (`MGR_DRAM_PBLC_CLINE_FIELD_MSB - `MGR_DRAM_PBLC_CLINE_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_CLINE_FIELD_RANGE        `MGR_DRAM_PBLC_CLINE_FIELD_MSB : `MGR_DRAM_PBLC_CLINE_FIELD_LSB

  // Remember, we increment bank/2, so reduce width by 1
  `define MGR_DRAM_PBLC_BANK_FIELD_WIDTH       `MGR_DRAM_BANK_ADDRESS_WIDTH-1
  `define MGR_DRAM_PBLC_BANK_FIELD_LSB         `MGR_DRAM_PBLC_CLINE_FIELD_MSB+1
  `define MGR_DRAM_PBLC_BANK_FIELD_MSB         `MGR_DRAM_PBLC_BANK_FIELD_LSB+`MGR_DRAM_PBLC_BANK_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_BANK_FIELD_SIZE        (`MGR_DRAM_PBLC_BANK_FIELD_MSB - `MGR_DRAM_PBLC_BANK_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_BANK_FIELD_RANGE        `MGR_DRAM_PBLC_BANK_FIELD_MSB : `MGR_DRAM_PBLC_BANK_FIELD_LSB
  
  `define MGR_DRAM_PBLC_PAGE_FIELD_WIDTH       `MGR_DRAM_PAGE_ADDRESS_WIDTH
  `define MGR_DRAM_PBLC_PAGE_FIELD_LSB         `MGR_DRAM_PBLC_BANK_FIELD_MSB+1
  `define MGR_DRAM_PBLC_PAGE_FIELD_MSB         `MGR_DRAM_PBLC_PAGE_FIELD_LSB+`MGR_DRAM_PBLC_PAGE_FIELD_WIDTH -1
  `define MGR_DRAM_PBLC_PAGE_FIELD_SIZE        (`MGR_DRAM_PBLC_PAGE_FIELD_MSB - `MGR_DRAM_PBLC_PAGE_FIELD_LSB +1)
  `define MGR_DRAM_PBLC_PAGE_FIELD_RANGE        `MGR_DRAM_PBLC_PAGE_FIELD_MSB : `MGR_DRAM_PBLC_PAGE_FIELD_LSB
  
  `define MGR_DRAM_PBLC_WIDTH                   `MGR_DRAM_PBLC_PAGE_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBLC_BANK_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBLC_CHAN_FIELD_WIDTH      \
                                               +`MGR_DRAM_PBLC_CLINE_FIELD_WIDTH       
  
  
  `define MGR_DRAM_PBLC_MSB            `MGR_DRAM_PBLC_WIDTH -1
  `define MGR_DRAM_PBLC_LSB            0
  `define MGR_DRAM_PBLC_SIZE           (`MGR_DRAM_PBLC_MSB - `MGR_DRAM_PBLC_LSB +1)
  `define MGR_DRAM_PBLC_RANGE           `MGR_DRAM_PBLC_MSB : `MGR_DRAM_PBLC_LSB

`endif


//---------------------------------------------------------------------------------------------------------------------
//---------------------------------------------------------------------------------------------------------------------
// NoC

//---------------------------------------------------------------------------------------------------------------------
// Internal
`define MGR_NOC_INTERNAL_DATA_WIDTH        `MGR_ARRAY_NOC_INTERNAL_DATA_WIDTH
`define MGR_NOC_INTERNAL_DATA_MSB          `MGR_NOC_INTERNAL_DATA_WIDTH-1
`define MGR_NOC_INTERNAL_DATA_LSB          0
`define MGR_NOC_INTERNAL_DATA_RANGE        `MGR_NOC_INTERNAL_DATA_MSB : `MGR_NOC_INTERNAL_DATA_LSB

`define MGR_NOC_INTERNAL_INTF_NUM_WORDS          `MGR_NOC_INTERNAL_DATA_WIDTH/32

`define MGR_NOC_INTERNAL_INTF_NUM_WORDS_WIDTH                       `MGR_NOC_INTERNAL_INTF_NUM_WORDS          
`define MGR_NOC_INTERNAL_INTF_NUM_WORDS_MSB                         `MGR_NOC_INTERNAL_INTF_NUM_WORDS_WIDTH-1
`define MGR_NOC_INTERNAL_INTF_NUM_WORDS_LSB                         0
`define MGR_NOC_INTERNAL_INTF_NUM_WORDS_SIZE                        (`MGR_NOC_INTERNAL_INTF_NUM_WORDS_MSB - `MGR_NOC_INTERNAL_INTF_NUM_WORDS_LSB +1)
`define MGR_NOC_INTERNAL_INTF_NUM_WORDS_RANGE                        `MGR_NOC_INTERNAL_INTF_NUM_WORDS_MSB : `MGR_NOC_INTERNAL_INTF_NUM_WORDS_LSB


//---------------------------------------------------------------------------------------------------------------------
// External
`define MGR_NOC_EXTERNAL_DATA_WIDTH        `MGR_ARRAY_NOC_EXTERNAL_DATA_WIDTH 
`define MGR_NOC_EXTERNAL_DATA_MSB          `MGR_NOC_EXTERNAL_DATA_WIDTH-1
`define MGR_NOC_EXTERNAL_DATA_LSB          0
`define MGR_NOC_EXTERNAL_DATA_RANGE        `MGR_NOC_EXTERNAL_DATA_MSB : `MGR_NOC_EXTERNAL_DATA_LSB


//---------------------------------------------------------------------------------------------------------------------
// MCast group
// - table is 64 entries

`define MGR_NOC_MCAST_GROUP_PTR_DEPTH   64
`define MGR_NOC_MCAST_GROUP_PTR_WIDTH   (`CLOG2(`MGR_NOC_MCAST_GROUP_PTR_DEPTH ))
`define MGR_NOC_MCAST_GROUP_PTR_MSB     `MGR_NOC_MCAST_GROUP_PTR_WIDTH-1
`define MGR_NOC_MCAST_GROUP_PTR_LSB     0
`define MGR_NOC_MCAST_GROUP_PTR_SIZE    (`MGR_NOC_MCAST_GROUP_PTR_MSB - `MGR_NOC_MCAST_GROUP_PTR_LSB +1)
`define MGR_NOC_MCAST_GROUP_PTR_RANGE    `MGR_NOC_MCAST_GROUP_PTR_MSB : `MGR_NOC_MCAST_GROUP_PTR_LSB




`endif
