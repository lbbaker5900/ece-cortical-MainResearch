
   // lane0 from NoC 
   wire                                            sdp__cntl__lane0_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane0_strm_cntl       ; 
   reg                                             cntl__sdp__lane0_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane0_strm_data       ; 
   reg                                             cntl__sdp__lane0_strm_data_valid ; 
   // lane0 to NoC 
   wire                                            cntl__sdp__lane0_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane0_strm_cntl       ; 
   wire                                            sdp__cntl__lane0_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane0_strm_data       ; 
   wire                                            sdp__cntl__lane0_strm_data_valid ; 
   // lane1 from NoC 
   wire                                            sdp__cntl__lane1_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane1_strm_cntl       ; 
   reg                                             cntl__sdp__lane1_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane1_strm_data       ; 
   reg                                             cntl__sdp__lane1_strm_data_valid ; 
   // lane1 to NoC 
   wire                                            cntl__sdp__lane1_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane1_strm_cntl       ; 
   wire                                            sdp__cntl__lane1_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane1_strm_data       ; 
   wire                                            sdp__cntl__lane1_strm_data_valid ; 
   // lane2 from NoC 
   wire                                            sdp__cntl__lane2_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane2_strm_cntl       ; 
   reg                                             cntl__sdp__lane2_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane2_strm_data       ; 
   reg                                             cntl__sdp__lane2_strm_data_valid ; 
   // lane2 to NoC 
   wire                                            cntl__sdp__lane2_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane2_strm_cntl       ; 
   wire                                            sdp__cntl__lane2_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane2_strm_data       ; 
   wire                                            sdp__cntl__lane2_strm_data_valid ; 
   // lane3 from NoC 
   wire                                            sdp__cntl__lane3_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane3_strm_cntl       ; 
   reg                                             cntl__sdp__lane3_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane3_strm_data       ; 
   reg                                             cntl__sdp__lane3_strm_data_valid ; 
   // lane3 to NoC 
   wire                                            cntl__sdp__lane3_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane3_strm_cntl       ; 
   wire                                            sdp__cntl__lane3_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane3_strm_data       ; 
   wire                                            sdp__cntl__lane3_strm_data_valid ; 
   // lane4 from NoC 
   wire                                            sdp__cntl__lane4_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane4_strm_cntl       ; 
   reg                                             cntl__sdp__lane4_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane4_strm_data       ; 
   reg                                             cntl__sdp__lane4_strm_data_valid ; 
   // lane4 to NoC 
   wire                                            cntl__sdp__lane4_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane4_strm_cntl       ; 
   wire                                            sdp__cntl__lane4_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane4_strm_data       ; 
   wire                                            sdp__cntl__lane4_strm_data_valid ; 
   // lane5 from NoC 
   wire                                            sdp__cntl__lane5_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane5_strm_cntl       ; 
   reg                                             cntl__sdp__lane5_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane5_strm_data       ; 
   reg                                             cntl__sdp__lane5_strm_data_valid ; 
   // lane5 to NoC 
   wire                                            cntl__sdp__lane5_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane5_strm_cntl       ; 
   wire                                            sdp__cntl__lane5_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane5_strm_data       ; 
   wire                                            sdp__cntl__lane5_strm_data_valid ; 
   // lane6 from NoC 
   wire                                            sdp__cntl__lane6_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane6_strm_cntl       ; 
   reg                                             cntl__sdp__lane6_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane6_strm_data       ; 
   reg                                             cntl__sdp__lane6_strm_data_valid ; 
   // lane6 to NoC 
   wire                                            cntl__sdp__lane6_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane6_strm_cntl       ; 
   wire                                            sdp__cntl__lane6_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane6_strm_data       ; 
   wire                                            sdp__cntl__lane6_strm_data_valid ; 
   // lane7 from NoC 
   wire                                            sdp__cntl__lane7_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane7_strm_cntl       ; 
   reg                                             cntl__sdp__lane7_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane7_strm_data       ; 
   reg                                             cntl__sdp__lane7_strm_data_valid ; 
   // lane7 to NoC 
   wire                                            cntl__sdp__lane7_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane7_strm_cntl       ; 
   wire                                            sdp__cntl__lane7_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane7_strm_data       ; 
   wire                                            sdp__cntl__lane7_strm_data_valid ; 
   // lane8 from NoC 
   wire                                            sdp__cntl__lane8_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane8_strm_cntl       ; 
   reg                                             cntl__sdp__lane8_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane8_strm_data       ; 
   reg                                             cntl__sdp__lane8_strm_data_valid ; 
   // lane8 to NoC 
   wire                                            cntl__sdp__lane8_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane8_strm_cntl       ; 
   wire                                            sdp__cntl__lane8_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane8_strm_data       ; 
   wire                                            sdp__cntl__lane8_strm_data_valid ; 
   // lane9 from NoC 
   wire                                            sdp__cntl__lane9_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane9_strm_cntl       ; 
   reg                                             cntl__sdp__lane9_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane9_strm_data       ; 
   reg                                             cntl__sdp__lane9_strm_data_valid ; 
   // lane9 to NoC 
   wire                                            cntl__sdp__lane9_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane9_strm_cntl       ; 
   wire                                            sdp__cntl__lane9_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane9_strm_data       ; 
   wire                                            sdp__cntl__lane9_strm_data_valid ; 
   // lane10 from NoC 
   wire                                            sdp__cntl__lane10_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane10_strm_cntl       ; 
   reg                                             cntl__sdp__lane10_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane10_strm_data       ; 
   reg                                             cntl__sdp__lane10_strm_data_valid ; 
   // lane10 to NoC 
   wire                                            cntl__sdp__lane10_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane10_strm_cntl       ; 
   wire                                            sdp__cntl__lane10_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane10_strm_data       ; 
   wire                                            sdp__cntl__lane10_strm_data_valid ; 
   // lane11 from NoC 
   wire                                            sdp__cntl__lane11_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane11_strm_cntl       ; 
   reg                                             cntl__sdp__lane11_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane11_strm_data       ; 
   reg                                             cntl__sdp__lane11_strm_data_valid ; 
   // lane11 to NoC 
   wire                                            cntl__sdp__lane11_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane11_strm_cntl       ; 
   wire                                            sdp__cntl__lane11_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane11_strm_data       ; 
   wire                                            sdp__cntl__lane11_strm_data_valid ; 
   // lane12 from NoC 
   wire                                            sdp__cntl__lane12_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane12_strm_cntl       ; 
   reg                                             cntl__sdp__lane12_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane12_strm_data       ; 
   reg                                             cntl__sdp__lane12_strm_data_valid ; 
   // lane12 to NoC 
   wire                                            cntl__sdp__lane12_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane12_strm_cntl       ; 
   wire                                            sdp__cntl__lane12_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane12_strm_data       ; 
   wire                                            sdp__cntl__lane12_strm_data_valid ; 
   // lane13 from NoC 
   wire                                            sdp__cntl__lane13_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane13_strm_cntl       ; 
   reg                                             cntl__sdp__lane13_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane13_strm_data       ; 
   reg                                             cntl__sdp__lane13_strm_data_valid ; 
   // lane13 to NoC 
   wire                                            cntl__sdp__lane13_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane13_strm_cntl       ; 
   wire                                            sdp__cntl__lane13_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane13_strm_data       ; 
   wire                                            sdp__cntl__lane13_strm_data_valid ; 
   // lane14 from NoC 
   wire                                            sdp__cntl__lane14_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane14_strm_cntl       ; 
   reg                                             cntl__sdp__lane14_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane14_strm_data       ; 
   reg                                             cntl__sdp__lane14_strm_data_valid ; 
   // lane14 to NoC 
   wire                                            cntl__sdp__lane14_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane14_strm_cntl       ; 
   wire                                            sdp__cntl__lane14_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane14_strm_data       ; 
   wire                                            sdp__cntl__lane14_strm_data_valid ; 
   // lane15 from NoC 
   wire                                            sdp__cntl__lane15_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane15_strm_cntl       ; 
   reg                                             cntl__sdp__lane15_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane15_strm_data       ; 
   reg                                             cntl__sdp__lane15_strm_data_valid ; 
   // lane15 to NoC 
   wire                                            cntl__sdp__lane15_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane15_strm_cntl       ; 
   wire                                            sdp__cntl__lane15_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane15_strm_data       ; 
   wire                                            sdp__cntl__lane15_strm_data_valid ; 
   // lane16 from NoC 
   wire                                            sdp__cntl__lane16_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane16_strm_cntl       ; 
   reg                                             cntl__sdp__lane16_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane16_strm_data       ; 
   reg                                             cntl__sdp__lane16_strm_data_valid ; 
   // lane16 to NoC 
   wire                                            cntl__sdp__lane16_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane16_strm_cntl       ; 
   wire                                            sdp__cntl__lane16_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane16_strm_data       ; 
   wire                                            sdp__cntl__lane16_strm_data_valid ; 
   // lane17 from NoC 
   wire                                            sdp__cntl__lane17_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane17_strm_cntl       ; 
   reg                                             cntl__sdp__lane17_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane17_strm_data       ; 
   reg                                             cntl__sdp__lane17_strm_data_valid ; 
   // lane17 to NoC 
   wire                                            cntl__sdp__lane17_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane17_strm_cntl       ; 
   wire                                            sdp__cntl__lane17_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane17_strm_data       ; 
   wire                                            sdp__cntl__lane17_strm_data_valid ; 
   // lane18 from NoC 
   wire                                            sdp__cntl__lane18_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane18_strm_cntl       ; 
   reg                                             cntl__sdp__lane18_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane18_strm_data       ; 
   reg                                             cntl__sdp__lane18_strm_data_valid ; 
   // lane18 to NoC 
   wire                                            cntl__sdp__lane18_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane18_strm_cntl       ; 
   wire                                            sdp__cntl__lane18_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane18_strm_data       ; 
   wire                                            sdp__cntl__lane18_strm_data_valid ; 
   // lane19 from NoC 
   wire                                            sdp__cntl__lane19_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane19_strm_cntl       ; 
   reg                                             cntl__sdp__lane19_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane19_strm_data       ; 
   reg                                             cntl__sdp__lane19_strm_data_valid ; 
   // lane19 to NoC 
   wire                                            cntl__sdp__lane19_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane19_strm_cntl       ; 
   wire                                            sdp__cntl__lane19_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane19_strm_data       ; 
   wire                                            sdp__cntl__lane19_strm_data_valid ; 
   // lane20 from NoC 
   wire                                            sdp__cntl__lane20_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane20_strm_cntl       ; 
   reg                                             cntl__sdp__lane20_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane20_strm_data       ; 
   reg                                             cntl__sdp__lane20_strm_data_valid ; 
   // lane20 to NoC 
   wire                                            cntl__sdp__lane20_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane20_strm_cntl       ; 
   wire                                            sdp__cntl__lane20_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane20_strm_data       ; 
   wire                                            sdp__cntl__lane20_strm_data_valid ; 
   // lane21 from NoC 
   wire                                            sdp__cntl__lane21_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane21_strm_cntl       ; 
   reg                                             cntl__sdp__lane21_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane21_strm_data       ; 
   reg                                             cntl__sdp__lane21_strm_data_valid ; 
   // lane21 to NoC 
   wire                                            cntl__sdp__lane21_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane21_strm_cntl       ; 
   wire                                            sdp__cntl__lane21_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane21_strm_data       ; 
   wire                                            sdp__cntl__lane21_strm_data_valid ; 
   // lane22 from NoC 
   wire                                            sdp__cntl__lane22_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane22_strm_cntl       ; 
   reg                                             cntl__sdp__lane22_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane22_strm_data       ; 
   reg                                             cntl__sdp__lane22_strm_data_valid ; 
   // lane22 to NoC 
   wire                                            cntl__sdp__lane22_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane22_strm_cntl       ; 
   wire                                            sdp__cntl__lane22_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane22_strm_data       ; 
   wire                                            sdp__cntl__lane22_strm_data_valid ; 
   // lane23 from NoC 
   wire                                            sdp__cntl__lane23_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane23_strm_cntl       ; 
   reg                                             cntl__sdp__lane23_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane23_strm_data       ; 
   reg                                             cntl__sdp__lane23_strm_data_valid ; 
   // lane23 to NoC 
   wire                                            cntl__sdp__lane23_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane23_strm_cntl       ; 
   wire                                            sdp__cntl__lane23_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane23_strm_data       ; 
   wire                                            sdp__cntl__lane23_strm_data_valid ; 
   // lane24 from NoC 
   wire                                            sdp__cntl__lane24_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane24_strm_cntl       ; 
   reg                                             cntl__sdp__lane24_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane24_strm_data       ; 
   reg                                             cntl__sdp__lane24_strm_data_valid ; 
   // lane24 to NoC 
   wire                                            cntl__sdp__lane24_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane24_strm_cntl       ; 
   wire                                            sdp__cntl__lane24_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane24_strm_data       ; 
   wire                                            sdp__cntl__lane24_strm_data_valid ; 
   // lane25 from NoC 
   wire                                            sdp__cntl__lane25_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane25_strm_cntl       ; 
   reg                                             cntl__sdp__lane25_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane25_strm_data       ; 
   reg                                             cntl__sdp__lane25_strm_data_valid ; 
   // lane25 to NoC 
   wire                                            cntl__sdp__lane25_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane25_strm_cntl       ; 
   wire                                            sdp__cntl__lane25_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane25_strm_data       ; 
   wire                                            sdp__cntl__lane25_strm_data_valid ; 
   // lane26 from NoC 
   wire                                            sdp__cntl__lane26_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane26_strm_cntl       ; 
   reg                                             cntl__sdp__lane26_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane26_strm_data       ; 
   reg                                             cntl__sdp__lane26_strm_data_valid ; 
   // lane26 to NoC 
   wire                                            cntl__sdp__lane26_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane26_strm_cntl       ; 
   wire                                            sdp__cntl__lane26_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane26_strm_data       ; 
   wire                                            sdp__cntl__lane26_strm_data_valid ; 
   // lane27 from NoC 
   wire                                            sdp__cntl__lane27_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane27_strm_cntl       ; 
   reg                                             cntl__sdp__lane27_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane27_strm_data       ; 
   reg                                             cntl__sdp__lane27_strm_data_valid ; 
   // lane27 to NoC 
   wire                                            cntl__sdp__lane27_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane27_strm_cntl       ; 
   wire                                            sdp__cntl__lane27_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane27_strm_data       ; 
   wire                                            sdp__cntl__lane27_strm_data_valid ; 
   // lane28 from NoC 
   wire                                            sdp__cntl__lane28_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane28_strm_cntl       ; 
   reg                                             cntl__sdp__lane28_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane28_strm_data       ; 
   reg                                             cntl__sdp__lane28_strm_data_valid ; 
   // lane28 to NoC 
   wire                                            cntl__sdp__lane28_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane28_strm_cntl       ; 
   wire                                            sdp__cntl__lane28_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane28_strm_data       ; 
   wire                                            sdp__cntl__lane28_strm_data_valid ; 
   // lane29 from NoC 
   wire                                            sdp__cntl__lane29_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane29_strm_cntl       ; 
   reg                                             cntl__sdp__lane29_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane29_strm_data       ; 
   reg                                             cntl__sdp__lane29_strm_data_valid ; 
   // lane29 to NoC 
   wire                                            cntl__sdp__lane29_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane29_strm_cntl       ; 
   wire                                            sdp__cntl__lane29_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane29_strm_data       ; 
   wire                                            sdp__cntl__lane29_strm_data_valid ; 
   // lane30 from NoC 
   wire                                            sdp__cntl__lane30_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane30_strm_cntl       ; 
   reg                                             cntl__sdp__lane30_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane30_strm_data       ; 
   reg                                             cntl__sdp__lane30_strm_data_valid ; 
   // lane30 to NoC 
   wire                                            cntl__sdp__lane30_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane30_strm_cntl       ; 
   wire                                            sdp__cntl__lane30_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane30_strm_data       ; 
   wire                                            sdp__cntl__lane30_strm_data_valid ; 
   // lane31 from NoC 
   wire                                            sdp__cntl__lane31_strm_ready      ; 
   reg[`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]        cntl__sdp__lane31_strm_cntl       ; 
   reg                                             cntl__sdp__lane31_strm_id         ; 
   reg[`STREAMING_OP_CNTL_DATA_RANGE      ]        cntl__sdp__lane31_strm_data       ; 
   reg                                             cntl__sdp__lane31_strm_data_valid ; 
   // lane31 to NoC 
   wire                                            cntl__sdp__lane31_strm_ready      ; 
   wire [`STREAMING_OP_CNTL_STRM_CNTL_RANGE ]      sdp__cntl__lane31_strm_cntl       ; 
   wire                                            sdp__cntl__lane31_strm_id         ; 
   wire [`STREAMING_OP_CNTL_DATA_RANGE      ]      sdp__cntl__lane31_strm_data       ; 
   wire                                            sdp__cntl__lane31_strm_data_valid ; 
