
        // PE 0, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[0][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[0][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[0][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[0][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[0][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[0][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[0][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[0][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[0][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[0][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[0][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[0][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[0][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[0][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[0][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[0][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[0][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[0][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[0][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[0][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[0][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[0][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[0][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[0][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[0][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[0][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[0][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[0][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[0][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[0][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[0][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[0][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[0][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[0][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[0][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[0][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[0][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[0][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[0][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[0][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[0][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[0][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[0][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[0][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[0][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[0][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[0][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[0][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[0][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[0][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[0][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[0][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[0][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[0][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[0][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[0][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[0][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[0][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[0][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[0][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[0][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[0][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[0][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[0][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[0][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[0][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[0][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[0][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[0][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[0][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[0][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[0][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[0][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[0][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[0][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[0][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[0][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[0][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[0][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[0][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[0][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[0][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[0][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[0][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[0][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[0][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[0][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[0][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[0][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[0][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[0][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[0][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[0][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[0][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[0][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[0][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[0][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[0][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[0][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[0][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[0][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[0][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[0][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[0][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[0][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[0][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[0][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[0][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[0][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[0][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[0][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[0][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[0][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[0][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[0][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[0][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[0][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[0][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[0][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[0][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[0][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[0][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[0][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[0][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[0][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[0][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[0][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[0][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[0][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[0][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[0][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[0][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[0][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[0][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[0][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[0][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[0][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[0][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[0][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[0][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[0][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[0][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[0][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[0][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[0][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[0][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[0][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[0][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[0][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[0][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[0][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[0][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[0][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[0][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[0][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[0][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[0][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[0][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[0][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[0][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[0][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[0][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[0][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[0][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[0][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[0][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[0][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[0][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[0][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[0][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[0][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[0][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[0][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[0][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[0][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[0][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[0][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[0][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[0][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[0][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[0][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[0][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[0][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[0][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[0][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[0][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 0, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[0][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[0][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[0][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[0][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[0].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[0][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[0][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[0].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[0][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[1][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[1][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[1][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[1][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[1][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[1][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[1][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[1][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[1][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[1][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[1][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[1][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[1][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[1][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[1][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[1][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[1][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[1][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[1][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[1][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[1][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[1][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[1][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[1][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[1][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[1][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[1][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[1][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[1][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[1][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[1][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[1][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[1][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[1][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[1][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[1][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[1][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[1][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[1][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[1][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[1][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[1][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[1][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[1][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[1][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[1][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[1][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[1][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[1][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[1][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[1][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[1][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[1][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[1][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[1][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[1][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[1][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[1][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[1][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[1][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[1][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[1][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[1][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[1][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[1][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[1][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[1][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[1][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[1][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[1][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[1][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[1][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[1][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[1][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[1][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[1][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[1][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[1][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[1][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[1][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[1][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[1][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[1][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[1][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[1][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[1][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[1][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[1][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[1][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[1][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[1][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[1][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[1][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[1][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[1][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[1][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[1][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[1][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[1][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[1][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[1][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[1][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[1][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[1][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[1][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[1][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[1][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[1][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[1][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[1][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[1][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[1][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[1][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[1][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[1][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[1][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[1][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[1][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[1][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[1][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[1][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[1][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[1][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[1][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[1][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[1][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[1][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[1][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[1][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[1][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[1][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[1][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[1][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[1][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[1][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[1][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[1][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[1][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[1][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[1][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[1][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[1][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[1][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[1][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[1][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[1][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[1][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[1][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[1][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[1][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[1][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[1][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[1][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[1][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[1][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[1][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[1][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[1][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[1][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[1][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[1][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[1][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[1][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[1][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[1][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[1][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[1][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[1][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[1][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[1][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[1][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[1][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[1][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[1][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[1][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[1][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[1][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[1][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[1][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[1][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[1][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[1][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[1][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[1][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[1][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[1][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 1, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[1][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[1][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[1][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[1][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[1].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[1][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[1][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[1].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[1][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[2][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[2][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[2][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[2][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[2][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[2][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[2][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[2][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[2][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[2][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[2][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[2][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[2][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[2][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[2][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[2][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[2][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[2][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[2][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[2][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[2][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[2][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[2][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[2][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[2][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[2][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[2][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[2][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[2][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[2][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[2][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[2][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[2][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[2][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[2][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[2][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[2][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[2][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[2][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[2][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[2][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[2][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[2][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[2][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[2][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[2][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[2][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[2][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[2][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[2][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[2][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[2][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[2][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[2][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[2][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[2][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[2][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[2][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[2][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[2][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[2][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[2][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[2][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[2][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[2][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[2][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[2][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[2][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[2][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[2][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[2][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[2][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[2][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[2][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[2][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[2][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[2][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[2][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[2][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[2][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[2][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[2][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[2][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[2][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[2][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[2][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[2][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[2][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[2][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[2][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[2][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[2][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[2][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[2][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[2][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[2][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[2][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[2][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[2][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[2][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[2][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[2][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[2][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[2][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[2][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[2][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[2][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[2][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[2][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[2][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[2][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[2][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[2][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[2][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[2][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[2][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[2][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[2][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[2][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[2][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[2][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[2][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[2][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[2][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[2][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[2][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[2][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[2][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[2][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[2][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[2][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[2][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[2][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[2][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[2][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[2][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[2][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[2][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[2][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[2][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[2][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[2][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[2][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[2][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[2][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[2][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[2][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[2][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[2][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[2][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[2][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[2][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[2][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[2][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[2][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[2][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[2][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[2][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[2][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[2][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[2][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[2][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[2][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[2][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[2][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[2][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[2][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[2][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[2][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[2][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[2][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[2][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[2][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[2][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[2][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[2][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[2][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[2][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[2][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[2][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[2][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[2][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[2][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[2][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[2][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[2][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 2, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[2][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[2][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[2][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[2][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[2].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[2][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[2][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[2].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[2][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[3][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[3][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[3][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[3][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[3][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[3][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[3][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[3][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[3][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[3][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[3][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[3][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[3][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[3][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[3][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[3][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[3][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[3][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[3][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[3][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[3][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[3][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[3][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[3][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[3][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[3][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[3][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[3][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[3][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[3][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[3][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[3][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[3][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[3][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[3][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[3][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[3][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[3][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[3][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[3][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[3][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[3][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[3][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[3][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[3][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[3][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[3][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[3][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[3][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[3][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[3][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[3][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[3][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[3][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[3][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[3][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[3][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[3][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[3][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[3][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[3][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[3][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[3][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[3][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[3][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[3][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[3][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[3][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[3][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[3][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[3][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[3][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[3][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[3][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[3][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[3][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[3][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[3][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[3][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[3][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[3][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[3][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[3][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[3][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[3][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[3][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[3][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[3][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[3][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[3][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[3][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[3][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[3][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[3][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[3][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[3][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[3][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[3][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[3][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[3][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[3][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[3][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[3][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[3][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[3][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[3][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[3][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[3][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[3][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[3][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[3][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[3][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[3][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[3][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[3][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[3][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[3][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[3][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[3][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[3][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[3][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[3][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[3][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[3][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[3][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[3][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[3][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[3][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[3][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[3][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[3][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[3][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[3][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[3][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[3][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[3][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[3][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[3][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[3][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[3][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[3][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[3][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[3][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[3][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[3][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[3][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[3][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[3][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[3][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[3][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[3][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[3][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[3][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[3][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[3][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[3][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[3][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[3][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[3][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[3][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[3][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[3][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[3][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[3][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[3][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[3][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[3][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[3][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[3][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[3][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[3][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[3][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[3][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[3][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[3][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[3][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[3][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[3][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[3][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[3][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[3][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[3][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[3][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[3][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[3][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[3][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 3, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[3][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[3][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[3][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[3][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[3].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[3][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[3][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[3].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[3][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[4][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[4][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[4][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[4][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[4][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[4][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[4][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[4][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[4][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[4][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[4][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[4][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[4][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[4][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[4][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[4][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[4][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[4][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[4][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[4][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[4][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[4][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[4][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[4][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[4][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[4][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[4][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[4][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[4][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[4][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[4][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[4][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[4][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[4][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[4][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[4][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[4][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[4][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[4][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[4][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[4][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[4][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[4][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[4][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[4][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[4][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[4][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[4][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[4][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[4][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[4][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[4][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[4][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[4][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[4][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[4][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[4][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[4][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[4][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[4][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[4][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[4][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[4][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[4][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[4][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[4][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[4][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[4][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[4][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[4][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[4][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[4][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[4][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[4][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[4][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[4][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[4][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[4][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[4][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[4][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[4][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[4][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[4][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[4][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[4][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[4][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[4][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[4][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[4][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[4][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[4][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[4][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[4][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[4][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[4][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[4][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[4][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[4][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[4][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[4][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[4][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[4][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[4][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[4][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[4][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[4][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[4][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[4][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[4][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[4][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[4][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[4][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[4][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[4][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[4][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[4][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[4][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[4][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[4][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[4][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[4][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[4][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[4][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[4][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[4][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[4][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[4][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[4][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[4][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[4][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[4][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[4][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[4][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[4][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[4][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[4][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[4][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[4][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[4][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[4][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[4][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[4][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[4][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[4][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[4][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[4][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[4][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[4][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[4][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[4][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[4][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[4][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[4][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[4][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[4][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[4][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[4][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[4][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[4][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[4][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[4][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[4][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[4][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[4][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[4][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[4][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[4][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[4][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[4][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[4][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[4][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[4][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[4][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[4][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[4][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[4][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[4][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[4][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[4][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[4][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[4][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[4][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[4][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[4][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[4][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[4][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 4, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[4][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[4][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[4][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[4][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[4].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[4][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[4][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[4].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[4][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[5][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[5][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[5][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[5][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[5][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[5][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[5][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[5][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[5][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[5][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[5][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[5][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[5][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[5][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[5][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[5][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[5][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[5][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[5][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[5][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[5][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[5][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[5][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[5][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[5][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[5][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[5][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[5][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[5][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[5][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[5][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[5][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[5][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[5][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[5][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[5][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[5][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[5][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[5][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[5][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[5][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[5][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[5][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[5][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[5][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[5][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[5][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[5][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[5][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[5][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[5][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[5][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[5][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[5][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[5][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[5][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[5][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[5][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[5][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[5][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[5][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[5][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[5][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[5][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[5][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[5][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[5][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[5][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[5][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[5][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[5][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[5][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[5][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[5][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[5][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[5][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[5][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[5][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[5][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[5][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[5][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[5][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[5][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[5][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[5][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[5][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[5][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[5][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[5][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[5][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[5][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[5][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[5][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[5][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[5][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[5][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[5][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[5][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[5][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[5][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[5][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[5][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[5][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[5][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[5][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[5][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[5][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[5][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[5][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[5][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[5][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[5][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[5][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[5][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[5][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[5][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[5][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[5][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[5][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[5][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[5][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[5][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[5][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[5][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[5][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[5][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[5][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[5][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[5][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[5][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[5][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[5][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[5][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[5][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[5][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[5][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[5][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[5][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[5][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[5][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[5][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[5][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[5][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[5][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[5][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[5][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[5][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[5][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[5][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[5][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[5][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[5][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[5][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[5][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[5][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[5][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[5][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[5][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[5][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[5][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[5][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[5][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[5][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[5][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[5][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[5][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[5][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[5][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[5][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[5][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[5][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[5][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[5][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[5][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[5][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[5][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[5][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[5][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[5][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[5][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[5][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[5][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[5][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[5][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[5][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[5][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 5, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[5][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[5][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[5][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[5][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[5].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[5][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[5][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[5].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[5][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[6][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[6][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[6][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[6][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[6][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[6][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[6][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[6][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[6][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[6][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[6][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[6][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[6][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[6][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[6][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[6][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[6][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[6][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[6][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[6][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[6][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[6][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[6][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[6][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[6][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[6][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[6][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[6][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[6][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[6][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[6][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[6][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[6][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[6][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[6][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[6][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[6][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[6][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[6][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[6][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[6][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[6][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[6][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[6][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[6][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[6][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[6][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[6][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[6][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[6][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[6][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[6][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[6][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[6][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[6][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[6][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[6][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[6][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[6][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[6][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[6][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[6][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[6][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[6][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[6][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[6][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[6][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[6][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[6][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[6][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[6][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[6][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[6][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[6][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[6][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[6][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[6][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[6][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[6][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[6][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[6][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[6][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[6][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[6][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[6][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[6][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[6][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[6][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[6][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[6][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[6][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[6][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[6][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[6][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[6][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[6][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[6][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[6][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[6][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[6][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[6][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[6][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[6][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[6][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[6][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[6][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[6][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[6][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[6][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[6][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[6][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[6][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[6][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[6][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[6][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[6][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[6][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[6][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[6][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[6][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[6][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[6][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[6][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[6][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[6][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[6][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[6][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[6][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[6][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[6][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[6][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[6][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[6][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[6][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[6][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[6][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[6][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[6][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[6][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[6][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[6][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[6][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[6][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[6][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[6][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[6][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[6][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[6][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[6][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[6][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[6][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[6][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[6][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[6][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[6][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[6][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[6][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[6][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[6][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[6][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[6][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[6][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[6][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[6][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[6][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[6][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[6][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[6][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[6][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[6][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[6][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[6][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[6][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[6][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[6][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[6][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[6][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[6][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[6][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[6][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[6][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[6][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[6][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[6][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[6][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[6][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 6, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[6][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[6][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[6][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[6][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[6].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[6][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[6][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[6].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[6][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[7][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[7][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[7][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[7][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[7][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[7][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[7][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[7][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[7][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[7][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[7][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[7][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[7][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[7][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[7][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[7][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[7][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[7][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[7][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[7][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[7][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[7][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[7][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[7][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[7][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[7][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[7][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[7][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[7][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[7][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[7][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[7][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[7][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[7][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[7][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[7][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[7][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[7][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[7][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[7][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[7][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[7][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[7][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[7][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[7][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[7][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[7][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[7][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[7][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[7][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[7][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[7][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[7][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[7][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[7][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[7][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[7][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[7][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[7][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[7][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[7][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[7][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[7][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[7][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[7][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[7][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[7][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[7][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[7][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[7][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[7][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[7][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[7][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[7][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[7][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[7][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[7][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[7][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[7][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[7][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[7][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[7][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[7][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[7][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[7][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[7][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[7][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[7][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[7][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[7][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[7][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[7][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[7][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[7][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[7][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[7][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[7][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[7][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[7][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[7][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[7][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[7][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[7][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[7][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[7][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[7][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[7][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[7][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[7][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[7][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[7][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[7][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[7][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[7][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[7][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[7][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[7][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[7][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[7][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[7][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[7][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[7][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[7][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[7][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[7][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[7][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[7][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[7][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[7][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[7][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[7][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[7][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[7][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[7][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[7][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[7][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[7][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[7][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[7][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[7][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[7][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[7][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[7][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[7][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[7][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[7][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[7][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[7][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[7][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[7][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[7][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[7][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[7][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[7][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[7][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[7][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[7][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[7][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[7][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[7][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[7][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[7][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[7][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[7][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[7][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[7][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[7][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[7][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[7][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[7][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[7][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[7][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[7][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[7][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[7][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[7][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[7][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[7][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[7][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[7][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[7][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[7][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[7][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[7][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[7][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[7][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 7, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[7][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[7][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[7][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[7][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[7].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[7][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[7][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[7].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[7][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[8][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[8][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[8][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[8][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[8][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[8][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[8][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[8][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[8][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[8][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[8][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[8][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[8][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[8][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[8][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[8][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[8][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[8][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[8][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[8][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[8][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[8][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[8][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[8][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[8][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[8][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[8][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[8][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[8][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[8][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[8][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[8][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[8][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[8][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[8][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[8][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[8][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[8][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[8][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[8][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[8][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[8][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[8][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[8][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[8][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[8][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[8][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[8][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[8][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[8][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[8][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[8][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[8][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[8][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[8][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[8][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[8][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[8][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[8][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[8][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[8][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[8][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[8][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[8][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[8][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[8][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[8][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[8][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[8][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[8][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[8][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[8][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[8][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[8][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[8][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[8][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[8][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[8][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[8][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[8][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[8][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[8][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[8][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[8][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[8][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[8][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[8][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[8][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[8][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[8][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[8][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[8][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[8][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[8][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[8][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[8][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[8][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[8][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[8][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[8][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[8][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[8][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[8][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[8][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[8][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[8][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[8][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[8][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[8][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[8][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[8][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[8][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[8][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[8][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[8][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[8][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[8][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[8][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[8][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[8][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[8][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[8][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[8][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[8][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[8][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[8][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[8][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[8][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[8][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[8][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[8][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[8][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[8][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[8][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[8][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[8][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[8][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[8][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[8][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[8][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[8][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[8][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[8][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[8][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[8][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[8][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[8][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[8][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[8][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[8][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[8][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[8][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[8][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[8][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[8][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[8][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[8][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[8][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[8][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[8][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[8][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[8][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[8][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[8][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[8][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[8][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[8][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[8][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[8][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[8][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[8][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[8][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[8][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[8][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[8][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[8][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[8][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[8][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[8][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[8][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[8][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[8][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[8][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[8][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[8][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[8][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 8, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[8][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[8][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[8][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[8][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[8].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[8][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[8][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[8].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[8][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[9][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[9][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[9][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[9][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[9][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[9][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[9][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[9][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[9][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[9][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[9][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[9][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[9][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[9][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[9][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[9][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[9][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[9][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[9][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[9][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[9][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[9][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[9][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[9][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[9][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[9][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[9][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[9][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[9][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[9][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[9][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[9][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[9][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[9][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[9][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[9][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[9][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[9][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[9][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[9][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[9][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[9][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[9][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[9][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[9][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[9][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[9][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[9][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[9][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[9][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[9][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[9][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[9][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[9][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[9][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[9][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[9][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[9][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[9][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[9][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[9][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[9][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[9][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[9][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[9][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[9][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[9][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[9][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[9][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[9][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[9][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[9][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[9][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[9][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[9][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[9][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[9][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[9][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[9][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[9][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[9][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[9][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[9][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[9][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[9][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[9][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[9][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[9][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[9][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[9][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[9][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[9][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[9][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[9][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[9][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[9][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[9][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[9][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[9][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[9][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[9][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[9][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[9][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[9][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[9][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[9][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[9][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[9][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[9][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[9][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[9][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[9][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[9][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[9][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[9][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[9][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[9][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[9][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[9][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[9][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[9][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[9][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[9][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[9][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[9][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[9][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[9][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[9][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[9][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[9][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[9][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[9][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[9][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[9][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[9][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[9][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[9][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[9][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[9][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[9][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[9][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[9][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[9][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[9][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[9][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[9][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[9][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[9][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[9][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[9][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[9][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[9][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[9][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[9][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[9][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[9][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[9][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[9][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[9][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[9][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[9][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[9][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[9][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[9][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[9][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[9][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[9][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[9][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[9][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[9][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[9][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[9][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[9][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[9][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[9][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[9][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[9][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[9][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[9][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[9][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[9][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[9][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[9][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[9][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[9][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[9][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 9, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[9][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[9][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[9][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[9][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[9].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[9][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[9][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[9].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[9][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[10][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[10][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[10][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[10][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[10][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[10][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[10][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[10][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[10][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[10][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[10][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[10][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[10][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[10][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[10][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[10][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[10][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[10][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[10][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[10][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[10][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[10][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[10][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[10][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[10][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[10][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[10][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[10][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[10][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[10][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[10][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[10][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[10][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[10][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[10][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[10][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[10][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[10][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[10][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[10][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[10][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[10][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[10][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[10][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[10][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[10][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[10][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[10][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[10][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[10][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[10][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[10][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[10][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[10][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[10][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[10][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[10][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[10][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[10][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[10][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[10][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[10][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[10][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[10][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[10][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[10][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[10][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[10][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[10][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[10][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[10][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[10][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[10][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[10][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[10][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[10][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[10][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[10][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[10][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[10][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[10][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[10][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[10][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[10][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[10][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[10][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[10][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[10][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[10][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[10][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[10][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[10][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[10][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[10][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[10][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[10][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[10][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[10][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[10][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[10][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[10][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[10][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[10][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[10][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[10][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[10][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[10][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[10][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[10][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[10][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[10][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[10][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[10][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[10][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[10][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[10][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[10][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[10][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[10][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[10][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[10][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[10][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[10][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[10][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[10][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[10][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[10][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[10][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[10][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[10][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[10][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[10][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[10][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[10][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[10][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[10][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[10][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[10][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[10][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[10][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[10][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[10][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[10][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[10][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[10][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[10][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[10][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[10][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[10][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[10][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[10][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[10][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[10][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[10][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[10][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[10][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[10][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[10][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[10][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[10][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[10][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[10][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[10][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[10][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[10][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[10][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[10][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[10][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[10][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[10][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[10][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[10][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[10][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[10][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[10][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[10][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[10][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[10][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[10][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[10][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[10][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[10][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[10][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[10][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[10][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[10][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 10, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[10][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[10][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[10][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[10][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[10].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[10][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[10][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[10].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[10][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[11][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[11][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[11][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[11][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[11][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[11][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[11][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[11][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[11][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[11][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[11][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[11][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[11][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[11][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[11][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[11][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[11][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[11][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[11][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[11][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[11][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[11][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[11][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[11][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[11][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[11][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[11][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[11][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[11][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[11][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[11][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[11][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[11][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[11][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[11][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[11][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[11][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[11][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[11][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[11][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[11][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[11][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[11][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[11][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[11][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[11][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[11][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[11][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[11][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[11][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[11][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[11][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[11][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[11][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[11][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[11][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[11][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[11][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[11][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[11][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[11][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[11][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[11][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[11][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[11][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[11][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[11][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[11][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[11][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[11][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[11][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[11][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[11][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[11][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[11][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[11][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[11][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[11][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[11][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[11][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[11][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[11][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[11][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[11][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[11][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[11][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[11][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[11][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[11][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[11][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[11][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[11][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[11][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[11][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[11][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[11][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[11][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[11][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[11][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[11][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[11][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[11][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[11][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[11][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[11][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[11][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[11][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[11][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[11][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[11][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[11][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[11][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[11][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[11][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[11][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[11][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[11][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[11][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[11][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[11][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[11][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[11][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[11][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[11][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[11][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[11][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[11][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[11][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[11][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[11][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[11][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[11][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[11][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[11][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[11][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[11][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[11][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[11][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[11][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[11][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[11][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[11][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[11][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[11][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[11][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[11][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[11][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[11][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[11][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[11][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[11][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[11][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[11][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[11][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[11][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[11][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[11][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[11][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[11][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[11][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[11][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[11][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[11][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[11][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[11][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[11][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[11][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[11][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[11][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[11][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[11][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[11][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[11][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[11][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[11][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[11][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[11][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[11][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[11][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[11][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[11][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[11][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[11][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[11][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[11][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[11][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 11, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[11][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[11][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[11][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[11][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[11].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[11][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[11][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[11].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[11][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[12][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[12][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[12][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[12][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[12][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[12][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[12][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[12][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[12][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[12][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[12][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[12][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[12][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[12][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[12][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[12][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[12][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[12][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[12][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[12][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[12][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[12][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[12][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[12][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[12][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[12][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[12][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[12][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[12][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[12][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[12][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[12][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[12][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[12][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[12][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[12][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[12][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[12][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[12][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[12][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[12][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[12][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[12][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[12][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[12][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[12][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[12][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[12][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[12][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[12][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[12][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[12][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[12][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[12][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[12][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[12][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[12][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[12][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[12][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[12][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[12][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[12][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[12][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[12][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[12][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[12][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[12][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[12][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[12][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[12][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[12][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[12][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[12][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[12][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[12][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[12][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[12][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[12][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[12][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[12][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[12][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[12][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[12][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[12][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[12][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[12][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[12][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[12][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[12][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[12][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[12][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[12][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[12][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[12][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[12][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[12][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[12][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[12][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[12][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[12][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[12][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[12][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[12][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[12][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[12][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[12][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[12][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[12][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[12][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[12][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[12][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[12][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[12][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[12][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[12][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[12][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[12][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[12][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[12][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[12][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[12][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[12][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[12][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[12][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[12][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[12][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[12][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[12][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[12][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[12][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[12][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[12][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[12][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[12][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[12][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[12][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[12][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[12][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[12][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[12][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[12][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[12][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[12][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[12][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[12][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[12][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[12][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[12][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[12][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[12][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[12][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[12][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[12][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[12][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[12][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[12][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[12][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[12][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[12][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[12][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[12][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[12][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[12][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[12][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[12][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[12][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[12][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[12][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[12][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[12][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[12][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[12][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[12][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[12][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[12][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[12][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[12][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[12][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[12][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[12][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[12][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[12][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[12][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[12][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[12][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[12][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 12, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[12][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[12][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[12][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[12][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[12].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[12][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[12][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[12].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[12][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[13][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[13][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[13][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[13][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[13][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[13][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[13][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[13][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[13][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[13][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[13][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[13][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[13][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[13][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[13][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[13][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[13][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[13][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[13][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[13][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[13][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[13][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[13][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[13][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[13][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[13][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[13][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[13][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[13][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[13][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[13][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[13][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[13][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[13][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[13][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[13][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[13][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[13][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[13][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[13][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[13][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[13][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[13][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[13][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[13][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[13][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[13][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[13][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[13][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[13][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[13][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[13][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[13][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[13][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[13][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[13][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[13][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[13][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[13][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[13][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[13][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[13][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[13][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[13][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[13][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[13][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[13][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[13][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[13][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[13][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[13][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[13][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[13][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[13][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[13][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[13][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[13][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[13][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[13][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[13][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[13][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[13][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[13][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[13][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[13][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[13][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[13][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[13][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[13][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[13][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[13][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[13][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[13][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[13][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[13][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[13][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[13][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[13][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[13][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[13][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[13][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[13][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[13][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[13][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[13][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[13][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[13][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[13][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[13][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[13][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[13][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[13][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[13][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[13][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[13][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[13][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[13][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[13][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[13][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[13][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[13][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[13][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[13][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[13][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[13][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[13][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[13][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[13][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[13][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[13][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[13][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[13][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[13][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[13][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[13][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[13][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[13][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[13][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[13][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[13][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[13][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[13][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[13][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[13][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[13][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[13][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[13][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[13][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[13][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[13][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[13][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[13][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[13][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[13][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[13][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[13][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[13][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[13][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[13][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[13][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[13][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[13][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[13][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[13][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[13][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[13][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[13][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[13][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[13][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[13][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[13][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[13][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[13][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[13][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[13][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[13][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[13][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[13][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[13][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[13][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[13][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[13][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[13][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[13][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[13][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[13][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 13, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[13][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[13][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[13][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[13][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[13].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[13][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[13][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[13].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[13][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[14][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[14][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[14][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[14][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[14][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[14][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[14][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[14][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[14][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[14][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[14][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[14][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[14][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[14][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[14][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[14][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[14][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[14][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[14][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[14][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[14][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[14][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[14][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[14][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[14][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[14][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[14][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[14][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[14][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[14][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[14][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[14][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[14][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[14][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[14][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[14][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[14][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[14][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[14][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[14][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[14][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[14][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[14][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[14][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[14][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[14][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[14][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[14][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[14][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[14][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[14][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[14][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[14][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[14][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[14][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[14][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[14][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[14][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[14][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[14][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[14][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[14][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[14][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[14][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[14][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[14][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[14][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[14][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[14][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[14][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[14][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[14][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[14][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[14][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[14][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[14][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[14][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[14][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[14][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[14][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[14][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[14][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[14][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[14][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[14][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[14][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[14][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[14][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[14][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[14][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[14][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[14][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[14][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[14][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[14][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[14][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[14][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[14][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[14][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[14][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[14][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[14][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[14][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[14][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[14][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[14][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[14][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[14][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[14][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[14][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[14][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[14][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[14][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[14][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[14][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[14][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[14][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[14][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[14][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[14][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[14][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[14][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[14][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[14][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[14][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[14][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[14][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[14][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[14][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[14][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[14][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[14][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[14][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[14][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[14][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[14][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[14][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[14][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[14][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[14][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[14][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[14][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[14][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[14][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[14][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[14][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[14][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[14][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[14][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[14][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[14][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[14][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[14][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[14][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[14][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[14][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[14][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[14][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[14][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[14][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[14][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[14][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[14][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[14][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[14][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[14][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[14][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[14][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[14][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[14][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[14][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[14][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[14][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[14][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[14][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[14][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[14][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[14][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[14][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[14][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[14][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[14][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[14][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[14][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[14][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[14][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 14, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[14][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[14][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[14][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[14][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[14].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[14][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[14][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[14].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[14][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[15][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[15][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[15][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[15][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[15][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[15][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[15][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[15][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[15][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[15][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[15][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[15][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[15][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[15][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[15][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[15][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[15][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[15][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[15][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[15][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[15][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[15][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[15][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[15][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[15][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[15][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[15][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[15][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[15][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[15][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[15][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[15][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[15][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[15][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[15][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[15][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[15][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[15][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[15][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[15][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[15][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[15][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[15][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[15][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[15][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[15][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[15][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[15][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[15][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[15][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[15][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[15][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[15][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[15][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[15][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[15][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[15][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[15][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[15][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[15][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[15][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[15][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[15][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[15][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[15][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[15][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[15][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[15][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[15][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[15][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[15][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[15][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[15][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[15][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[15][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[15][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[15][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[15][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[15][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[15][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[15][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[15][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[15][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[15][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[15][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[15][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[15][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[15][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[15][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[15][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[15][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[15][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[15][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[15][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[15][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[15][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[15][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[15][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[15][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[15][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[15][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[15][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[15][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[15][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[15][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[15][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[15][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[15][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[15][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[15][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[15][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[15][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[15][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[15][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[15][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[15][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[15][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[15][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[15][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[15][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[15][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[15][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[15][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[15][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[15][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[15][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[15][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[15][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[15][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[15][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[15][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[15][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[15][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[15][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[15][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[15][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[15][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[15][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[15][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[15][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[15][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[15][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[15][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[15][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[15][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[15][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[15][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[15][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[15][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[15][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[15][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[15][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[15][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[15][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[15][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[15][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[15][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[15][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[15][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[15][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[15][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[15][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[15][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[15][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[15][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[15][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[15][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[15][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[15][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[15][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[15][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[15][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[15][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[15][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[15][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[15][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[15][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[15][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[15][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[15][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[15][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[15][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[15][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[15][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[15][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[15][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 15, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[15][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[15][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[15][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[15][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[15].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[15][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[15][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[15].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[15][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[16][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[16][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[16][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[16][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[16][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[16][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[16][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[16][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[16][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[16][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[16][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[16][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[16][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[16][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[16][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[16][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[16][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[16][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[16][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[16][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[16][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[16][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[16][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[16][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[16][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[16][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[16][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[16][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[16][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[16][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[16][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[16][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[16][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[16][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[16][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[16][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[16][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[16][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[16][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[16][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[16][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[16][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[16][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[16][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[16][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[16][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[16][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[16][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[16][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[16][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[16][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[16][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[16][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[16][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[16][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[16][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[16][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[16][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[16][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[16][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[16][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[16][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[16][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[16][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[16][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[16][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[16][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[16][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[16][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[16][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[16][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[16][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[16][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[16][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[16][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[16][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[16][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[16][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[16][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[16][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[16][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[16][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[16][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[16][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[16][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[16][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[16][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[16][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[16][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[16][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[16][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[16][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[16][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[16][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[16][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[16][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[16][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[16][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[16][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[16][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[16][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[16][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[16][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[16][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[16][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[16][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[16][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[16][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[16][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[16][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[16][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[16][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[16][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[16][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[16][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[16][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[16][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[16][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[16][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[16][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[16][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[16][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[16][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[16][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[16][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[16][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[16][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[16][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[16][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[16][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[16][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[16][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[16][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[16][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[16][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[16][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[16][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[16][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[16][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[16][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[16][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[16][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[16][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[16][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[16][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[16][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[16][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[16][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[16][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[16][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[16][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[16][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[16][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[16][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[16][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[16][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[16][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[16][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[16][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[16][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[16][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[16][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[16][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[16][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[16][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[16][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[16][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[16][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[16][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[16][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[16][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[16][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[16][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[16][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[16][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[16][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[16][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[16][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[16][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[16][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[16][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[16][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[16][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[16][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[16][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[16][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 16, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[16][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[16][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[16][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[16][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[16].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[16][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[16][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[16].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[16][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[17][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[17][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[17][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[17][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[17][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[17][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[17][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[17][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[17][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[17][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[17][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[17][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[17][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[17][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[17][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[17][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[17][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[17][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[17][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[17][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[17][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[17][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[17][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[17][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[17][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[17][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[17][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[17][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[17][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[17][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[17][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[17][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[17][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[17][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[17][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[17][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[17][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[17][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[17][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[17][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[17][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[17][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[17][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[17][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[17][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[17][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[17][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[17][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[17][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[17][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[17][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[17][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[17][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[17][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[17][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[17][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[17][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[17][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[17][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[17][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[17][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[17][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[17][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[17][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[17][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[17][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[17][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[17][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[17][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[17][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[17][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[17][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[17][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[17][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[17][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[17][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[17][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[17][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[17][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[17][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[17][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[17][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[17][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[17][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[17][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[17][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[17][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[17][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[17][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[17][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[17][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[17][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[17][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[17][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[17][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[17][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[17][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[17][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[17][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[17][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[17][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[17][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[17][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[17][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[17][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[17][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[17][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[17][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[17][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[17][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[17][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[17][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[17][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[17][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[17][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[17][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[17][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[17][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[17][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[17][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[17][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[17][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[17][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[17][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[17][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[17][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[17][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[17][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[17][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[17][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[17][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[17][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[17][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[17][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[17][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[17][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[17][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[17][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[17][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[17][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[17][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[17][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[17][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[17][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[17][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[17][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[17][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[17][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[17][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[17][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[17][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[17][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[17][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[17][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[17][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[17][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[17][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[17][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[17][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[17][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[17][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[17][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[17][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[17][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[17][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[17][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[17][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[17][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[17][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[17][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[17][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[17][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[17][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[17][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[17][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[17][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[17][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[17][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[17][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[17][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[17][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[17][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[17][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[17][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[17][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[17][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 17, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[17][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[17][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[17][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[17][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[17].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[17][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[17][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[17].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[17][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[18][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[18][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[18][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[18][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[18][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[18][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[18][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[18][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[18][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[18][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[18][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[18][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[18][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[18][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[18][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[18][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[18][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[18][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[18][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[18][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[18][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[18][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[18][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[18][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[18][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[18][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[18][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[18][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[18][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[18][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[18][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[18][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[18][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[18][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[18][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[18][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[18][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[18][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[18][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[18][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[18][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[18][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[18][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[18][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[18][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[18][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[18][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[18][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[18][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[18][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[18][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[18][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[18][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[18][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[18][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[18][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[18][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[18][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[18][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[18][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[18][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[18][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[18][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[18][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[18][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[18][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[18][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[18][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[18][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[18][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[18][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[18][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[18][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[18][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[18][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[18][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[18][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[18][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[18][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[18][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[18][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[18][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[18][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[18][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[18][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[18][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[18][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[18][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[18][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[18][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[18][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[18][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[18][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[18][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[18][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[18][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[18][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[18][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[18][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[18][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[18][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[18][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[18][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[18][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[18][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[18][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[18][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[18][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[18][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[18][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[18][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[18][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[18][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[18][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[18][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[18][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[18][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[18][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[18][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[18][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[18][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[18][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[18][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[18][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[18][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[18][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[18][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[18][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[18][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[18][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[18][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[18][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[18][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[18][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[18][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[18][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[18][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[18][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[18][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[18][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[18][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[18][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[18][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[18][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[18][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[18][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[18][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[18][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[18][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[18][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[18][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[18][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[18][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[18][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[18][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[18][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[18][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[18][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[18][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[18][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[18][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[18][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[18][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[18][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[18][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[18][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[18][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[18][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[18][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[18][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[18][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[18][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[18][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[18][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[18][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[18][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[18][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[18][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[18][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[18][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[18][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[18][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[18][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[18][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[18][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[18][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 18, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[18][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[18][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[18][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[18][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[18].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[18][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[18][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[18].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[18][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[19][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[19][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[19][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[19][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[19][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[19][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[19][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[19][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[19][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[19][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[19][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[19][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[19][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[19][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[19][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[19][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[19][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[19][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[19][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[19][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[19][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[19][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[19][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[19][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[19][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[19][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[19][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[19][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[19][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[19][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[19][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[19][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[19][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[19][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[19][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[19][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[19][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[19][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[19][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[19][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[19][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[19][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[19][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[19][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[19][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[19][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[19][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[19][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[19][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[19][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[19][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[19][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[19][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[19][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[19][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[19][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[19][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[19][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[19][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[19][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[19][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[19][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[19][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[19][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[19][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[19][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[19][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[19][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[19][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[19][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[19][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[19][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[19][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[19][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[19][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[19][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[19][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[19][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[19][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[19][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[19][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[19][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[19][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[19][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[19][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[19][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[19][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[19][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[19][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[19][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[19][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[19][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[19][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[19][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[19][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[19][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[19][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[19][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[19][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[19][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[19][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[19][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[19][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[19][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[19][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[19][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[19][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[19][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[19][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[19][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[19][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[19][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[19][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[19][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[19][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[19][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[19][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[19][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[19][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[19][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[19][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[19][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[19][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[19][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[19][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[19][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[19][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[19][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[19][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[19][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[19][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[19][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[19][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[19][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[19][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[19][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[19][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[19][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[19][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[19][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[19][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[19][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[19][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[19][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[19][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[19][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[19][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[19][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[19][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[19][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[19][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[19][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[19][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[19][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[19][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[19][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[19][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[19][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[19][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[19][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[19][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[19][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[19][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[19][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[19][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[19][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[19][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[19][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[19][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[19][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[19][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[19][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[19][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[19][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[19][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[19][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[19][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[19][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[19][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[19][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[19][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[19][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[19][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[19][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[19][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[19][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 19, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[19][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[19][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[19][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[19][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[19].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[19][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[19][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[19].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[19][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[20][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[20][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[20][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[20][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[20][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[20][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[20][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[20][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[20][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[20][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[20][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[20][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[20][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[20][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[20][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[20][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[20][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[20][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[20][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[20][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[20][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[20][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[20][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[20][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[20][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[20][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[20][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[20][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[20][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[20][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[20][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[20][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[20][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[20][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[20][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[20][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[20][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[20][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[20][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[20][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[20][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[20][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[20][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[20][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[20][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[20][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[20][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[20][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[20][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[20][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[20][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[20][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[20][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[20][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[20][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[20][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[20][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[20][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[20][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[20][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[20][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[20][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[20][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[20][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[20][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[20][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[20][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[20][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[20][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[20][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[20][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[20][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[20][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[20][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[20][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[20][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[20][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[20][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[20][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[20][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[20][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[20][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[20][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[20][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[20][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[20][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[20][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[20][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[20][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[20][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[20][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[20][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[20][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[20][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[20][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[20][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[20][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[20][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[20][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[20][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[20][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[20][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[20][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[20][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[20][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[20][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[20][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[20][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[20][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[20][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[20][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[20][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[20][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[20][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[20][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[20][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[20][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[20][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[20][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[20][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[20][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[20][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[20][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[20][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[20][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[20][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[20][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[20][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[20][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[20][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[20][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[20][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[20][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[20][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[20][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[20][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[20][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[20][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[20][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[20][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[20][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[20][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[20][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[20][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[20][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[20][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[20][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[20][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[20][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[20][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[20][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[20][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[20][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[20][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[20][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[20][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[20][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[20][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[20][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[20][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[20][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[20][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[20][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[20][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[20][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[20][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[20][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[20][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[20][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[20][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[20][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[20][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[20][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[20][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[20][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[20][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[20][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[20][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[20][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[20][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[20][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[20][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[20][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[20][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[20][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[20][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 20, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[20][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[20][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[20][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[20][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[20].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[20][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[20][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[20].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[20][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[21][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[21][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[21][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[21][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[21][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[21][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[21][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[21][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[21][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[21][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[21][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[21][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[21][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[21][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[21][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[21][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[21][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[21][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[21][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[21][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[21][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[21][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[21][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[21][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[21][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[21][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[21][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[21][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[21][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[21][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[21][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[21][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[21][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[21][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[21][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[21][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[21][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[21][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[21][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[21][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[21][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[21][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[21][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[21][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[21][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[21][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[21][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[21][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[21][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[21][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[21][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[21][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[21][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[21][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[21][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[21][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[21][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[21][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[21][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[21][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[21][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[21][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[21][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[21][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[21][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[21][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[21][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[21][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[21][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[21][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[21][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[21][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[21][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[21][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[21][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[21][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[21][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[21][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[21][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[21][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[21][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[21][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[21][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[21][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[21][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[21][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[21][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[21][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[21][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[21][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[21][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[21][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[21][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[21][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[21][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[21][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[21][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[21][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[21][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[21][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[21][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[21][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[21][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[21][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[21][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[21][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[21][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[21][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[21][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[21][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[21][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[21][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[21][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[21][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[21][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[21][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[21][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[21][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[21][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[21][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[21][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[21][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[21][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[21][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[21][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[21][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[21][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[21][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[21][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[21][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[21][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[21][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[21][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[21][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[21][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[21][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[21][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[21][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[21][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[21][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[21][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[21][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[21][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[21][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[21][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[21][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[21][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[21][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[21][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[21][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[21][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[21][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[21][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[21][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[21][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[21][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[21][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[21][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[21][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[21][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[21][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[21][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[21][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[21][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[21][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[21][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[21][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[21][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[21][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[21][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[21][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[21][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[21][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[21][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[21][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[21][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[21][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[21][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[21][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[21][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[21][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[21][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[21][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[21][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[21][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[21][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 21, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[21][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[21][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[21][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[21][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[21].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[21][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[21][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[21].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[21][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[22][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[22][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[22][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[22][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[22][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[22][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[22][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[22][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[22][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[22][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[22][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[22][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[22][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[22][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[22][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[22][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[22][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[22][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[22][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[22][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[22][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[22][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[22][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[22][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[22][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[22][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[22][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[22][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[22][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[22][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[22][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[22][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[22][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[22][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[22][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[22][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[22][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[22][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[22][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[22][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[22][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[22][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[22][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[22][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[22][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[22][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[22][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[22][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[22][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[22][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[22][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[22][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[22][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[22][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[22][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[22][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[22][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[22][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[22][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[22][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[22][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[22][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[22][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[22][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[22][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[22][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[22][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[22][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[22][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[22][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[22][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[22][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[22][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[22][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[22][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[22][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[22][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[22][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[22][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[22][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[22][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[22][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[22][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[22][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[22][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[22][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[22][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[22][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[22][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[22][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[22][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[22][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[22][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[22][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[22][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[22][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[22][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[22][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[22][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[22][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[22][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[22][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[22][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[22][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[22][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[22][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[22][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[22][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[22][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[22][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[22][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[22][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[22][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[22][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[22][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[22][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[22][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[22][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[22][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[22][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[22][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[22][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[22][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[22][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[22][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[22][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[22][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[22][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[22][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[22][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[22][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[22][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[22][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[22][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[22][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[22][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[22][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[22][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[22][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[22][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[22][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[22][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[22][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[22][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[22][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[22][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[22][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[22][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[22][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[22][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[22][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[22][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[22][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[22][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[22][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[22][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[22][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[22][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[22][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[22][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[22][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[22][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[22][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[22][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[22][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[22][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[22][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[22][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[22][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[22][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[22][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[22][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[22][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[22][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[22][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[22][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[22][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[22][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[22][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[22][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[22][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[22][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[22][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[22][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[22][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[22][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 22, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[22][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[22][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[22][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[22][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[22].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[22][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[22][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[22].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[22][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[23][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[23][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[23][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[23][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[23][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[23][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[23][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[23][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[23][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[23][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[23][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[23][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[23][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[23][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[23][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[23][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[23][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[23][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[23][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[23][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[23][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[23][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[23][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[23][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[23][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[23][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[23][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[23][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[23][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[23][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[23][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[23][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[23][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[23][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[23][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[23][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[23][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[23][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[23][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[23][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[23][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[23][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[23][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[23][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[23][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[23][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[23][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[23][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[23][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[23][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[23][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[23][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[23][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[23][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[23][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[23][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[23][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[23][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[23][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[23][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[23][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[23][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[23][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[23][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[23][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[23][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[23][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[23][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[23][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[23][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[23][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[23][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[23][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[23][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[23][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[23][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[23][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[23][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[23][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[23][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[23][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[23][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[23][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[23][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[23][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[23][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[23][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[23][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[23][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[23][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[23][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[23][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[23][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[23][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[23][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[23][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[23][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[23][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[23][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[23][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[23][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[23][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[23][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[23][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[23][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[23][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[23][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[23][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[23][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[23][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[23][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[23][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[23][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[23][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[23][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[23][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[23][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[23][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[23][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[23][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[23][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[23][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[23][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[23][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[23][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[23][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[23][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[23][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[23][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[23][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[23][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[23][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[23][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[23][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[23][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[23][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[23][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[23][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[23][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[23][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[23][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[23][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[23][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[23][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[23][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[23][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[23][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[23][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[23][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[23][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[23][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[23][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[23][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[23][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[23][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[23][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[23][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[23][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[23][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[23][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[23][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[23][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[23][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[23][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[23][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[23][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[23][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[23][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[23][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[23][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[23][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[23][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[23][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[23][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[23][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[23][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[23][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[23][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[23][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[23][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[23][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[23][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[23][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[23][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[23][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[23][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 23, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[23][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[23][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[23][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[23][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[23].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[23][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[23][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[23].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[23][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[24][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[24][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[24][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[24][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[24][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[24][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[24][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[24][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[24][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[24][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[24][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[24][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[24][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[24][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[24][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[24][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[24][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[24][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[24][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[24][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[24][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[24][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[24][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[24][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[24][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[24][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[24][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[24][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[24][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[24][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[24][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[24][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[24][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[24][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[24][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[24][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[24][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[24][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[24][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[24][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[24][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[24][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[24][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[24][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[24][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[24][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[24][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[24][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[24][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[24][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[24][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[24][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[24][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[24][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[24][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[24][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[24][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[24][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[24][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[24][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[24][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[24][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[24][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[24][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[24][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[24][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[24][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[24][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[24][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[24][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[24][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[24][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[24][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[24][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[24][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[24][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[24][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[24][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[24][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[24][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[24][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[24][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[24][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[24][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[24][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[24][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[24][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[24][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[24][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[24][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[24][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[24][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[24][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[24][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[24][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[24][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[24][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[24][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[24][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[24][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[24][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[24][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[24][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[24][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[24][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[24][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[24][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[24][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[24][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[24][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[24][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[24][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[24][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[24][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[24][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[24][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[24][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[24][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[24][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[24][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[24][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[24][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[24][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[24][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[24][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[24][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[24][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[24][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[24][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[24][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[24][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[24][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[24][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[24][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[24][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[24][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[24][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[24][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[24][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[24][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[24][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[24][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[24][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[24][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[24][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[24][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[24][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[24][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[24][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[24][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[24][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[24][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[24][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[24][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[24][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[24][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[24][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[24][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[24][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[24][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[24][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[24][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[24][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[24][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[24][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[24][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[24][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[24][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[24][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[24][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[24][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[24][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[24][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[24][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[24][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[24][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[24][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[24][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[24][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[24][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[24][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[24][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[24][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[24][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[24][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[24][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 24, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[24][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[24][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[24][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[24][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[24].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[24][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[24][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[24].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[24][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[25][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[25][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[25][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[25][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[25][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[25][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[25][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[25][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[25][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[25][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[25][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[25][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[25][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[25][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[25][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[25][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[25][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[25][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[25][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[25][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[25][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[25][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[25][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[25][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[25][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[25][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[25][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[25][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[25][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[25][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[25][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[25][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[25][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[25][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[25][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[25][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[25][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[25][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[25][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[25][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[25][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[25][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[25][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[25][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[25][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[25][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[25][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[25][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[25][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[25][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[25][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[25][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[25][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[25][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[25][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[25][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[25][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[25][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[25][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[25][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[25][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[25][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[25][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[25][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[25][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[25][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[25][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[25][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[25][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[25][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[25][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[25][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[25][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[25][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[25][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[25][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[25][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[25][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[25][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[25][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[25][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[25][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[25][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[25][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[25][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[25][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[25][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[25][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[25][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[25][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[25][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[25][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[25][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[25][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[25][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[25][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[25][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[25][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[25][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[25][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[25][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[25][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[25][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[25][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[25][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[25][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[25][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[25][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[25][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[25][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[25][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[25][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[25][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[25][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[25][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[25][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[25][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[25][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[25][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[25][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[25][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[25][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[25][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[25][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[25][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[25][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[25][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[25][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[25][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[25][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[25][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[25][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[25][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[25][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[25][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[25][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[25][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[25][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[25][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[25][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[25][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[25][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[25][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[25][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[25][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[25][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[25][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[25][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[25][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[25][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[25][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[25][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[25][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[25][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[25][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[25][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[25][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[25][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[25][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[25][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[25][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[25][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[25][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[25][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[25][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[25][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[25][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[25][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[25][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[25][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[25][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[25][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[25][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[25][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[25][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[25][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[25][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[25][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[25][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[25][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[25][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[25][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[25][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[25][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[25][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[25][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 25, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[25][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[25][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[25][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[25][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[25].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[25][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[25][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[25].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[25][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[26][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[26][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[26][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[26][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[26][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[26][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[26][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[26][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[26][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[26][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[26][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[26][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[26][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[26][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[26][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[26][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[26][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[26][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[26][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[26][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[26][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[26][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[26][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[26][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[26][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[26][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[26][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[26][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[26][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[26][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[26][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[26][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[26][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[26][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[26][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[26][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[26][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[26][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[26][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[26][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[26][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[26][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[26][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[26][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[26][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[26][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[26][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[26][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[26][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[26][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[26][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[26][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[26][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[26][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[26][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[26][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[26][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[26][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[26][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[26][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[26][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[26][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[26][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[26][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[26][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[26][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[26][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[26][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[26][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[26][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[26][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[26][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[26][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[26][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[26][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[26][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[26][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[26][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[26][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[26][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[26][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[26][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[26][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[26][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[26][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[26][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[26][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[26][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[26][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[26][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[26][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[26][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[26][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[26][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[26][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[26][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[26][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[26][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[26][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[26][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[26][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[26][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[26][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[26][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[26][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[26][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[26][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[26][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[26][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[26][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[26][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[26][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[26][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[26][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[26][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[26][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[26][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[26][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[26][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[26][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[26][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[26][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[26][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[26][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[26][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[26][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[26][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[26][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[26][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[26][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[26][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[26][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[26][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[26][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[26][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[26][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[26][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[26][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[26][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[26][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[26][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[26][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[26][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[26][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[26][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[26][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[26][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[26][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[26][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[26][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[26][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[26][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[26][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[26][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[26][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[26][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[26][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[26][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[26][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[26][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[26][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[26][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[26][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[26][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[26][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[26][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[26][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[26][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[26][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[26][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[26][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[26][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[26][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[26][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[26][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[26][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[26][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[26][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[26][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[26][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[26][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[26][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[26][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[26][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[26][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[26][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 26, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[26][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[26][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[26][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[26][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[26].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[26][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[26][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[26].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[26][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[27][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[27][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[27][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[27][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[27][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[27][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[27][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[27][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[27][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[27][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[27][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[27][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[27][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[27][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[27][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[27][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[27][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[27][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[27][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[27][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[27][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[27][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[27][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[27][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[27][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[27][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[27][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[27][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[27][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[27][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[27][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[27][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[27][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[27][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[27][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[27][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[27][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[27][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[27][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[27][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[27][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[27][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[27][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[27][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[27][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[27][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[27][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[27][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[27][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[27][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[27][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[27][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[27][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[27][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[27][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[27][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[27][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[27][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[27][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[27][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[27][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[27][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[27][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[27][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[27][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[27][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[27][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[27][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[27][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[27][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[27][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[27][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[27][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[27][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[27][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[27][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[27][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[27][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[27][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[27][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[27][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[27][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[27][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[27][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[27][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[27][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[27][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[27][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[27][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[27][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[27][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[27][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[27][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[27][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[27][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[27][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[27][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[27][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[27][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[27][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[27][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[27][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[27][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[27][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[27][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[27][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[27][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[27][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[27][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[27][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[27][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[27][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[27][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[27][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[27][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[27][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[27][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[27][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[27][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[27][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[27][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[27][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[27][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[27][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[27][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[27][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[27][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[27][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[27][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[27][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[27][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[27][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[27][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[27][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[27][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[27][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[27][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[27][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[27][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[27][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[27][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[27][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[27][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[27][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[27][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[27][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[27][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[27][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[27][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[27][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[27][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[27][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[27][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[27][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[27][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[27][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[27][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[27][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[27][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[27][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[27][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[27][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[27][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[27][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[27][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[27][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[27][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[27][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[27][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[27][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[27][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[27][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[27][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[27][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[27][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[27][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[27][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[27][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[27][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[27][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[27][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[27][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[27][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[27][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[27][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[27][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 27, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[27][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[27][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[27][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[27][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[27].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[27][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[27][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[27].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[27][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[28][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[28][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[28][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[28][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[28][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[28][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[28][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[28][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[28][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[28][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[28][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[28][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[28][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[28][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[28][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[28][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[28][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[28][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[28][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[28][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[28][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[28][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[28][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[28][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[28][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[28][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[28][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[28][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[28][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[28][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[28][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[28][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[28][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[28][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[28][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[28][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[28][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[28][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[28][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[28][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[28][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[28][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[28][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[28][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[28][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[28][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[28][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[28][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[28][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[28][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[28][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[28][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[28][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[28][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[28][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[28][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[28][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[28][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[28][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[28][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[28][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[28][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[28][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[28][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[28][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[28][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[28][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[28][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[28][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[28][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[28][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[28][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[28][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[28][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[28][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[28][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[28][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[28][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[28][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[28][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[28][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[28][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[28][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[28][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[28][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[28][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[28][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[28][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[28][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[28][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[28][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[28][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[28][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[28][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[28][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[28][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[28][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[28][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[28][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[28][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[28][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[28][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[28][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[28][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[28][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[28][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[28][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[28][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[28][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[28][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[28][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[28][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[28][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[28][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[28][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[28][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[28][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[28][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[28][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[28][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[28][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[28][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[28][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[28][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[28][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[28][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[28][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[28][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[28][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[28][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[28][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[28][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[28][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[28][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[28][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[28][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[28][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[28][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[28][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[28][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[28][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[28][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[28][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[28][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[28][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[28][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[28][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[28][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[28][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[28][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[28][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[28][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[28][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[28][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[28][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[28][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[28][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[28][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[28][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[28][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[28][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[28][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[28][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[28][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[28][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[28][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[28][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[28][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[28][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[28][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[28][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[28][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[28][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[28][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[28][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[28][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[28][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[28][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[28][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[28][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[28][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[28][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[28][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[28][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[28][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[28][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 28, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[28][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[28][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[28][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[28][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[28].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[28][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[28][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[28].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[28][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[29][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[29][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[29][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[29][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[29][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[29][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[29][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[29][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[29][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[29][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[29][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[29][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[29][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[29][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[29][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[29][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[29][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[29][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[29][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[29][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[29][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[29][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[29][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[29][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[29][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[29][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[29][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[29][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[29][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[29][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[29][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[29][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[29][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[29][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[29][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[29][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[29][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[29][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[29][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[29][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[29][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[29][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[29][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[29][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[29][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[29][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[29][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[29][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[29][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[29][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[29][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[29][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[29][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[29][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[29][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[29][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[29][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[29][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[29][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[29][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[29][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[29][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[29][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[29][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[29][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[29][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[29][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[29][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[29][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[29][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[29][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[29][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[29][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[29][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[29][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[29][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[29][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[29][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[29][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[29][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[29][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[29][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[29][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[29][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[29][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[29][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[29][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[29][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[29][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[29][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[29][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[29][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[29][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[29][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[29][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[29][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[29][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[29][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[29][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[29][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[29][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[29][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[29][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[29][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[29][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[29][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[29][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[29][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[29][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[29][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[29][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[29][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[29][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[29][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[29][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[29][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[29][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[29][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[29][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[29][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[29][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[29][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[29][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[29][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[29][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[29][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[29][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[29][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[29][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[29][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[29][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[29][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[29][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[29][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[29][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[29][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[29][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[29][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[29][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[29][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[29][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[29][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[29][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[29][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[29][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[29][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[29][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[29][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[29][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[29][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[29][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[29][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[29][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[29][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[29][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[29][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[29][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[29][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[29][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[29][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[29][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[29][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[29][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[29][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[29][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[29][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[29][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[29][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[29][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[29][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[29][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[29][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[29][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[29][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[29][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[29][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[29][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[29][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[29][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[29][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[29][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[29][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[29][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[29][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[29][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[29][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 29, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[29][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[29][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[29][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[29][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[29].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[29][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[29][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[29].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[29][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[30][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[30][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[30][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[30][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[30][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[30][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[30][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[30][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[30][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[30][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[30][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[30][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[30][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[30][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[30][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[30][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[30][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[30][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[30][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[30][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[30][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[30][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[30][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[30][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[30][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[30][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[30][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[30][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[30][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[30][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[30][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[30][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[30][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[30][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[30][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[30][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[30][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[30][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[30][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[30][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[30][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[30][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[30][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[30][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[30][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[30][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[30][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[30][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[30][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[30][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[30][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[30][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[30][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[30][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[30][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[30][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[30][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[30][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[30][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[30][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[30][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[30][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[30][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[30][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[30][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[30][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[30][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[30][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[30][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[30][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[30][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[30][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[30][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[30][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[30][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[30][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[30][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[30][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[30][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[30][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[30][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[30][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[30][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[30][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[30][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[30][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[30][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[30][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[30][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[30][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[30][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[30][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[30][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[30][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[30][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[30][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[30][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[30][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[30][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[30][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[30][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[30][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[30][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[30][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[30][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[30][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[30][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[30][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[30][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[30][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[30][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[30][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[30][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[30][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[30][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[30][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[30][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[30][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[30][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[30][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[30][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[30][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[30][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[30][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[30][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[30][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[30][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[30][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[30][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[30][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[30][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[30][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[30][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[30][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[30][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[30][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[30][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[30][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[30][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[30][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[30][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[30][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[30][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[30][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[30][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[30][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[30][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[30][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[30][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[30][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[30][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[30][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[30][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[30][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[30][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[30][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[30][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[30][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[30][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[30][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[30][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[30][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[30][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[30][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[30][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[30][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[30][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[30][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[30][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[30][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[30][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[30][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[30][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[30][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[30][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[30][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[30][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[30][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[30][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[30][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[30][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[30][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[30][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[30][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[30][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[30][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 30, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[30][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[30][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[30][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[30][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[30].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[30][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[30][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[30].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[30][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[31][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[31][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[31][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[31][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[31][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[31][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[31][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[31][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[31][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[31][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[31][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[31][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[31][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[31][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[31][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[31][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[31][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[31][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[31][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[31][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[31][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[31][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[31][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[31][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[31][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[31][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[31][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[31][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[31][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[31][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[31][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[31][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[31][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[31][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[31][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[31][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[31][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[31][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[31][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[31][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[31][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[31][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[31][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[31][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[31][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[31][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[31][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[31][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[31][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[31][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[31][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[31][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[31][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[31][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[31][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[31][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[31][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[31][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[31][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[31][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[31][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[31][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[31][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[31][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[31][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[31][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[31][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[31][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[31][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[31][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[31][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[31][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[31][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[31][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[31][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[31][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[31][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[31][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[31][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[31][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[31][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[31][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[31][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[31][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[31][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[31][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[31][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[31][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[31][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[31][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[31][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[31][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[31][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[31][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[31][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[31][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[31][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[31][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[31][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[31][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[31][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[31][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[31][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[31][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[31][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[31][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[31][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[31][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[31][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[31][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[31][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[31][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[31][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[31][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[31][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[31][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[31][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[31][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[31][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[31][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[31][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[31][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[31][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[31][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[31][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[31][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[31][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[31][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[31][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[31][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[31][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[31][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[31][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[31][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[31][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[31][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[31][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[31][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[31][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[31][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[31][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[31][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[31][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[31][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[31][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[31][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[31][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[31][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[31][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[31][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[31][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[31][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[31][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[31][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[31][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[31][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[31][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[31][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[31][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[31][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[31][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[31][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[31][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[31][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[31][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[31][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[31][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[31][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[31][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[31][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[31][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[31][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[31][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[31][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[31][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[31][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[31][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[31][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[31][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[31][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[31][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[31][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[31][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[31][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[31][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[31][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 31, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[31][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[31][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[31][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[31][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[31].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[31][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[31][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[31].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[31][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[32][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[32][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[32][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[32][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[32][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[32][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[32][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[32][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[32][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[32][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[32][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[32][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[32][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[32][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[32][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[32][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[32][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[32][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[32][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[32][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[32][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[32][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[32][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[32][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[32][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[32][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[32][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[32][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[32][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[32][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[32][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[32][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[32][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[32][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[32][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[32][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[32][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[32][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[32][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[32][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[32][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[32][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[32][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[32][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[32][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[32][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[32][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[32][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[32][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[32][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[32][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[32][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[32][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[32][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[32][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[32][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[32][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[32][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[32][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[32][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[32][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[32][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[32][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[32][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[32][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[32][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[32][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[32][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[32][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[32][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[32][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[32][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[32][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[32][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[32][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[32][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[32][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[32][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[32][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[32][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[32][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[32][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[32][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[32][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[32][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[32][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[32][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[32][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[32][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[32][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[32][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[32][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[32][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[32][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[32][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[32][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[32][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[32][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[32][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[32][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[32][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[32][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[32][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[32][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[32][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[32][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[32][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[32][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[32][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[32][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[32][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[32][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[32][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[32][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[32][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[32][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[32][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[32][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[32][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[32][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[32][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[32][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[32][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[32][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[32][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[32][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[32][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[32][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[32][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[32][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[32][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[32][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[32][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[32][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[32][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[32][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[32][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[32][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[32][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[32][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[32][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[32][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[32][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[32][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[32][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[32][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[32][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[32][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[32][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[32][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[32][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[32][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[32][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[32][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[32][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[32][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[32][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[32][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[32][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[32][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[32][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[32][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[32][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[32][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[32][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[32][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[32][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[32][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[32][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[32][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[32][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[32][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[32][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[32][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[32][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[32][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[32][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[32][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[32][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[32][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[32][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[32][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[32][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[32][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[32][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[32][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 32, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[32][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[32][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[32][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[32][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[32].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[32][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[32][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[32].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[32][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[33][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[33][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[33][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[33][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[33][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[33][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[33][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[33][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[33][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[33][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[33][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[33][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[33][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[33][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[33][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[33][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[33][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[33][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[33][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[33][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[33][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[33][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[33][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[33][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[33][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[33][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[33][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[33][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[33][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[33][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[33][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[33][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[33][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[33][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[33][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[33][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[33][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[33][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[33][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[33][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[33][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[33][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[33][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[33][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[33][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[33][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[33][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[33][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[33][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[33][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[33][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[33][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[33][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[33][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[33][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[33][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[33][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[33][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[33][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[33][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[33][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[33][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[33][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[33][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[33][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[33][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[33][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[33][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[33][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[33][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[33][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[33][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[33][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[33][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[33][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[33][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[33][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[33][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[33][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[33][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[33][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[33][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[33][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[33][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[33][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[33][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[33][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[33][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[33][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[33][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[33][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[33][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[33][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[33][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[33][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[33][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[33][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[33][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[33][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[33][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[33][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[33][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[33][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[33][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[33][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[33][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[33][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[33][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[33][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[33][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[33][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[33][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[33][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[33][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[33][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[33][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[33][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[33][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[33][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[33][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[33][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[33][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[33][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[33][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[33][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[33][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[33][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[33][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[33][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[33][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[33][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[33][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[33][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[33][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[33][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[33][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[33][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[33][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[33][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[33][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[33][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[33][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[33][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[33][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[33][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[33][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[33][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[33][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[33][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[33][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[33][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[33][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[33][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[33][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[33][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[33][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[33][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[33][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[33][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[33][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[33][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[33][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[33][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[33][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[33][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[33][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[33][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[33][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[33][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[33][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[33][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[33][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[33][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[33][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[33][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[33][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[33][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[33][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[33][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[33][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[33][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[33][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[33][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[33][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[33][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[33][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 33, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[33][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[33][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[33][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[33][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[33].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[33][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[33][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[33].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[33][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[34][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[34][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[34][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[34][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[34][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[34][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[34][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[34][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[34][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[34][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[34][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[34][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[34][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[34][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[34][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[34][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[34][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[34][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[34][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[34][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[34][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[34][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[34][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[34][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[34][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[34][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[34][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[34][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[34][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[34][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[34][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[34][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[34][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[34][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[34][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[34][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[34][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[34][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[34][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[34][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[34][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[34][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[34][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[34][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[34][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[34][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[34][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[34][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[34][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[34][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[34][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[34][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[34][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[34][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[34][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[34][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[34][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[34][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[34][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[34][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[34][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[34][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[34][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[34][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[34][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[34][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[34][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[34][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[34][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[34][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[34][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[34][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[34][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[34][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[34][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[34][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[34][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[34][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[34][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[34][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[34][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[34][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[34][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[34][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[34][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[34][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[34][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[34][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[34][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[34][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[34][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[34][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[34][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[34][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[34][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[34][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[34][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[34][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[34][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[34][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[34][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[34][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[34][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[34][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[34][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[34][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[34][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[34][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[34][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[34][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[34][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[34][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[34][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[34][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[34][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[34][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[34][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[34][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[34][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[34][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[34][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[34][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[34][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[34][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[34][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[34][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[34][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[34][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[34][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[34][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[34][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[34][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[34][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[34][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[34][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[34][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[34][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[34][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[34][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[34][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[34][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[34][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[34][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[34][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[34][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[34][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[34][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[34][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[34][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[34][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[34][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[34][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[34][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[34][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[34][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[34][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[34][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[34][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[34][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[34][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[34][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[34][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[34][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[34][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[34][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[34][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[34][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[34][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[34][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[34][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[34][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[34][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[34][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[34][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[34][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[34][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[34][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[34][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[34][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[34][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[34][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[34][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[34][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[34][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[34][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[34][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 34, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[34][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[34][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[34][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[34][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[34].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[34][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[34][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[34].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[34][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[35][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[35][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[35][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[35][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[35][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[35][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[35][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[35][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[35][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[35][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[35][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[35][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[35][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[35][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[35][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[35][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[35][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[35][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[35][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[35][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[35][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[35][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[35][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[35][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[35][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[35][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[35][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[35][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[35][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[35][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[35][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[35][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[35][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[35][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[35][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[35][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[35][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[35][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[35][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[35][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[35][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[35][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[35][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[35][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[35][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[35][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[35][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[35][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[35][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[35][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[35][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[35][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[35][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[35][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[35][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[35][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[35][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[35][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[35][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[35][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[35][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[35][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[35][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[35][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[35][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[35][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[35][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[35][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[35][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[35][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[35][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[35][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[35][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[35][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[35][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[35][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[35][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[35][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[35][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[35][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[35][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[35][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[35][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[35][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[35][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[35][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[35][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[35][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[35][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[35][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[35][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[35][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[35][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[35][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[35][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[35][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[35][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[35][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[35][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[35][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[35][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[35][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[35][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[35][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[35][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[35][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[35][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[35][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[35][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[35][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[35][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[35][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[35][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[35][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[35][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[35][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[35][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[35][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[35][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[35][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[35][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[35][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[35][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[35][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[35][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[35][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[35][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[35][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[35][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[35][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[35][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[35][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[35][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[35][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[35][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[35][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[35][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[35][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[35][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[35][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[35][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[35][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[35][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[35][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[35][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[35][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[35][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[35][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[35][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[35][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[35][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[35][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[35][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[35][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[35][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[35][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[35][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[35][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[35][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[35][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[35][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[35][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[35][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[35][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[35][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[35][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[35][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[35][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[35][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[35][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[35][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[35][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[35][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[35][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[35][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[35][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[35][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[35][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[35][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[35][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[35][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[35][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[35][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[35][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[35][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[35][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 35, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[35][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[35][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[35][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[35][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[35].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[35][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[35][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[35].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[35][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[36][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[36][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[36][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[36][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[36][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[36][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[36][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[36][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[36][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[36][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[36][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[36][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[36][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[36][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[36][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[36][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[36][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[36][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[36][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[36][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[36][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[36][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[36][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[36][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[36][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[36][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[36][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[36][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[36][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[36][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[36][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[36][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[36][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[36][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[36][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[36][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[36][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[36][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[36][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[36][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[36][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[36][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[36][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[36][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[36][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[36][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[36][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[36][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[36][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[36][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[36][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[36][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[36][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[36][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[36][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[36][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[36][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[36][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[36][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[36][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[36][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[36][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[36][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[36][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[36][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[36][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[36][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[36][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[36][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[36][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[36][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[36][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[36][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[36][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[36][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[36][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[36][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[36][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[36][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[36][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[36][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[36][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[36][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[36][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[36][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[36][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[36][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[36][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[36][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[36][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[36][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[36][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[36][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[36][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[36][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[36][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[36][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[36][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[36][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[36][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[36][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[36][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[36][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[36][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[36][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[36][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[36][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[36][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[36][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[36][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[36][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[36][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[36][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[36][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[36][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[36][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[36][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[36][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[36][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[36][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[36][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[36][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[36][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[36][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[36][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[36][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[36][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[36][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[36][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[36][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[36][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[36][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[36][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[36][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[36][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[36][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[36][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[36][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[36][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[36][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[36][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[36][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[36][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[36][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[36][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[36][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[36][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[36][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[36][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[36][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[36][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[36][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[36][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[36][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[36][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[36][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[36][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[36][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[36][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[36][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[36][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[36][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[36][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[36][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[36][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[36][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[36][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[36][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[36][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[36][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[36][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[36][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[36][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[36][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[36][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[36][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[36][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[36][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[36][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[36][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[36][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[36][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[36][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[36][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[36][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[36][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 36, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[36][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[36][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[36][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[36][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[36].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[36][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[36][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[36].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[36][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[37][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[37][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[37][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[37][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[37][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[37][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[37][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[37][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[37][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[37][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[37][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[37][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[37][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[37][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[37][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[37][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[37][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[37][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[37][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[37][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[37][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[37][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[37][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[37][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[37][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[37][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[37][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[37][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[37][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[37][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[37][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[37][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[37][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[37][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[37][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[37][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[37][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[37][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[37][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[37][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[37][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[37][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[37][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[37][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[37][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[37][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[37][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[37][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[37][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[37][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[37][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[37][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[37][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[37][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[37][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[37][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[37][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[37][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[37][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[37][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[37][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[37][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[37][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[37][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[37][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[37][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[37][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[37][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[37][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[37][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[37][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[37][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[37][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[37][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[37][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[37][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[37][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[37][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[37][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[37][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[37][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[37][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[37][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[37][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[37][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[37][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[37][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[37][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[37][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[37][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[37][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[37][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[37][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[37][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[37][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[37][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[37][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[37][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[37][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[37][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[37][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[37][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[37][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[37][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[37][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[37][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[37][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[37][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[37][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[37][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[37][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[37][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[37][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[37][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[37][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[37][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[37][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[37][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[37][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[37][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[37][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[37][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[37][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[37][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[37][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[37][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[37][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[37][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[37][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[37][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[37][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[37][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[37][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[37][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[37][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[37][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[37][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[37][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[37][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[37][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[37][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[37][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[37][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[37][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[37][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[37][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[37][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[37][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[37][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[37][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[37][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[37][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[37][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[37][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[37][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[37][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[37][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[37][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[37][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[37][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[37][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[37][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[37][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[37][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[37][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[37][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[37][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[37][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[37][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[37][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[37][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[37][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[37][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[37][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[37][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[37][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[37][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[37][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[37][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[37][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[37][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[37][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[37][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[37][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[37][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[37][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 37, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[37][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[37][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[37][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[37][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[37].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[37][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[37][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[37].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[37][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[38][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[38][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[38][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[38][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[38][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[38][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[38][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[38][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[38][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[38][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[38][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[38][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[38][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[38][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[38][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[38][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[38][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[38][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[38][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[38][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[38][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[38][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[38][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[38][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[38][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[38][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[38][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[38][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[38][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[38][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[38][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[38][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[38][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[38][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[38][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[38][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[38][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[38][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[38][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[38][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[38][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[38][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[38][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[38][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[38][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[38][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[38][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[38][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[38][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[38][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[38][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[38][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[38][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[38][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[38][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[38][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[38][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[38][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[38][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[38][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[38][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[38][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[38][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[38][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[38][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[38][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[38][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[38][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[38][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[38][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[38][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[38][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[38][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[38][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[38][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[38][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[38][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[38][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[38][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[38][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[38][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[38][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[38][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[38][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[38][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[38][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[38][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[38][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[38][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[38][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[38][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[38][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[38][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[38][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[38][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[38][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[38][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[38][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[38][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[38][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[38][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[38][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[38][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[38][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[38][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[38][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[38][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[38][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[38][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[38][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[38][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[38][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[38][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[38][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[38][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[38][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[38][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[38][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[38][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[38][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[38][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[38][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[38][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[38][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[38][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[38][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[38][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[38][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[38][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[38][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[38][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[38][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[38][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[38][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[38][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[38][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[38][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[38][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[38][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[38][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[38][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[38][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[38][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[38][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[38][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[38][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[38][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[38][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[38][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[38][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[38][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[38][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[38][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[38][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[38][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[38][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[38][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[38][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[38][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[38][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[38][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[38][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[38][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[38][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[38][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[38][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[38][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[38][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[38][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[38][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[38][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[38][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[38][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[38][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[38][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[38][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[38][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[38][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[38][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[38][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[38][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[38][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[38][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[38][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[38][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[38][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 38, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[38][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[38][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[38][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[38][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[38].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[38][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[38][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[38].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[38][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[39][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[39][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[39][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[39][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[39][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[39][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[39][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[39][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[39][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[39][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[39][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[39][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[39][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[39][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[39][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[39][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[39][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[39][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[39][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[39][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[39][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[39][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[39][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[39][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[39][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[39][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[39][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[39][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[39][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[39][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[39][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[39][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[39][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[39][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[39][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[39][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[39][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[39][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[39][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[39][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[39][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[39][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[39][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[39][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[39][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[39][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[39][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[39][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[39][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[39][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[39][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[39][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[39][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[39][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[39][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[39][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[39][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[39][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[39][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[39][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[39][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[39][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[39][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[39][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[39][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[39][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[39][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[39][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[39][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[39][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[39][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[39][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[39][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[39][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[39][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[39][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[39][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[39][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[39][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[39][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[39][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[39][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[39][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[39][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[39][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[39][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[39][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[39][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[39][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[39][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[39][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[39][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[39][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[39][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[39][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[39][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[39][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[39][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[39][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[39][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[39][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[39][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[39][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[39][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[39][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[39][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[39][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[39][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[39][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[39][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[39][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[39][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[39][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[39][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[39][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[39][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[39][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[39][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[39][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[39][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[39][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[39][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[39][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[39][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[39][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[39][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[39][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[39][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[39][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[39][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[39][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[39][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[39][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[39][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[39][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[39][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[39][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[39][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[39][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[39][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[39][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[39][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[39][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[39][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[39][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[39][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[39][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[39][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[39][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[39][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[39][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[39][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[39][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[39][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[39][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[39][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[39][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[39][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[39][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[39][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[39][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[39][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[39][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[39][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[39][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[39][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[39][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[39][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[39][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[39][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[39][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[39][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[39][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[39][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[39][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[39][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[39][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[39][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[39][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[39][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[39][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[39][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[39][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[39][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[39][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[39][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 39, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[39][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[39][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[39][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[39][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[39].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[39][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[39][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[39].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[39][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[40][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[40][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[40][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[40][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[40][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[40][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[40][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[40][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[40][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[40][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[40][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[40][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[40][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[40][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[40][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[40][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[40][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[40][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[40][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[40][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[40][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[40][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[40][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[40][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[40][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[40][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[40][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[40][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[40][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[40][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[40][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[40][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[40][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[40][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[40][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[40][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[40][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[40][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[40][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[40][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[40][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[40][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[40][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[40][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[40][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[40][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[40][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[40][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[40][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[40][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[40][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[40][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[40][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[40][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[40][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[40][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[40][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[40][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[40][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[40][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[40][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[40][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[40][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[40][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[40][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[40][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[40][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[40][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[40][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[40][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[40][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[40][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[40][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[40][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[40][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[40][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[40][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[40][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[40][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[40][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[40][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[40][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[40][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[40][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[40][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[40][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[40][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[40][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[40][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[40][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[40][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[40][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[40][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[40][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[40][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[40][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[40][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[40][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[40][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[40][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[40][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[40][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[40][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[40][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[40][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[40][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[40][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[40][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[40][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[40][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[40][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[40][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[40][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[40][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[40][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[40][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[40][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[40][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[40][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[40][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[40][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[40][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[40][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[40][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[40][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[40][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[40][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[40][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[40][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[40][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[40][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[40][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[40][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[40][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[40][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[40][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[40][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[40][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[40][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[40][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[40][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[40][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[40][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[40][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[40][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[40][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[40][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[40][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[40][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[40][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[40][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[40][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[40][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[40][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[40][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[40][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[40][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[40][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[40][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[40][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[40][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[40][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[40][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[40][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[40][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[40][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[40][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[40][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[40][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[40][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[40][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[40][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[40][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[40][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[40][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[40][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[40][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[40][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[40][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[40][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[40][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[40][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[40][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[40][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[40][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[40][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 40, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[40][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[40][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[40][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[40][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[40].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[40][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[40][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[40].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[40][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[41][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[41][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[41][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[41][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[41][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[41][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[41][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[41][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[41][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[41][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[41][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[41][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[41][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[41][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[41][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[41][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[41][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[41][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[41][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[41][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[41][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[41][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[41][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[41][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[41][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[41][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[41][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[41][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[41][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[41][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[41][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[41][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[41][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[41][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[41][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[41][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[41][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[41][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[41][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[41][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[41][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[41][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[41][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[41][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[41][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[41][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[41][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[41][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[41][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[41][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[41][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[41][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[41][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[41][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[41][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[41][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[41][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[41][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[41][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[41][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[41][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[41][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[41][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[41][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[41][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[41][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[41][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[41][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[41][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[41][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[41][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[41][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[41][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[41][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[41][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[41][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[41][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[41][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[41][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[41][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[41][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[41][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[41][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[41][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[41][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[41][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[41][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[41][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[41][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[41][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[41][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[41][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[41][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[41][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[41][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[41][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[41][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[41][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[41][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[41][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[41][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[41][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[41][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[41][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[41][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[41][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[41][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[41][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[41][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[41][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[41][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[41][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[41][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[41][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[41][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[41][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[41][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[41][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[41][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[41][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[41][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[41][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[41][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[41][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[41][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[41][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[41][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[41][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[41][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[41][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[41][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[41][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[41][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[41][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[41][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[41][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[41][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[41][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[41][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[41][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[41][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[41][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[41][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[41][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[41][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[41][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[41][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[41][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[41][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[41][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[41][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[41][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[41][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[41][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[41][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[41][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[41][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[41][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[41][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[41][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[41][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[41][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[41][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[41][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[41][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[41][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[41][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[41][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[41][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[41][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[41][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[41][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[41][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[41][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[41][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[41][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[41][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[41][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[41][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[41][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[41][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[41][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[41][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[41][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[41][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[41][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 41, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[41][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[41][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[41][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[41][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[41].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[41][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[41][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[41].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[41][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[42][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[42][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[42][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[42][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[42][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[42][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[42][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[42][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[42][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[42][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[42][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[42][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[42][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[42][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[42][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[42][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[42][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[42][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[42][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[42][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[42][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[42][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[42][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[42][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[42][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[42][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[42][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[42][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[42][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[42][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[42][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[42][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[42][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[42][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[42][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[42][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[42][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[42][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[42][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[42][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[42][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[42][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[42][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[42][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[42][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[42][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[42][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[42][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[42][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[42][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[42][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[42][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[42][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[42][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[42][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[42][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[42][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[42][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[42][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[42][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[42][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[42][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[42][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[42][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[42][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[42][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[42][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[42][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[42][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[42][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[42][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[42][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[42][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[42][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[42][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[42][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[42][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[42][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[42][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[42][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[42][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[42][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[42][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[42][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[42][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[42][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[42][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[42][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[42][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[42][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[42][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[42][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[42][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[42][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[42][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[42][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[42][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[42][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[42][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[42][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[42][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[42][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[42][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[42][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[42][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[42][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[42][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[42][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[42][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[42][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[42][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[42][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[42][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[42][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[42][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[42][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[42][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[42][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[42][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[42][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[42][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[42][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[42][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[42][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[42][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[42][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[42][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[42][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[42][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[42][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[42][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[42][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[42][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[42][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[42][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[42][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[42][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[42][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[42][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[42][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[42][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[42][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[42][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[42][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[42][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[42][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[42][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[42][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[42][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[42][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[42][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[42][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[42][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[42][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[42][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[42][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[42][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[42][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[42][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[42][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[42][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[42][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[42][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[42][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[42][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[42][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[42][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[42][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[42][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[42][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[42][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[42][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[42][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[42][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[42][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[42][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[42][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[42][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[42][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[42][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[42][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[42][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[42][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[42][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[42][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[42][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 42, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[42][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[42][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[42][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[42][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[42].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[42][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[42][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[42].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[42][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[43][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[43][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[43][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[43][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[43][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[43][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[43][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[43][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[43][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[43][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[43][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[43][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[43][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[43][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[43][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[43][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[43][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[43][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[43][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[43][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[43][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[43][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[43][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[43][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[43][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[43][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[43][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[43][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[43][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[43][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[43][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[43][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[43][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[43][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[43][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[43][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[43][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[43][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[43][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[43][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[43][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[43][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[43][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[43][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[43][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[43][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[43][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[43][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[43][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[43][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[43][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[43][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[43][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[43][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[43][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[43][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[43][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[43][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[43][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[43][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[43][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[43][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[43][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[43][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[43][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[43][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[43][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[43][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[43][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[43][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[43][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[43][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[43][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[43][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[43][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[43][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[43][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[43][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[43][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[43][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[43][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[43][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[43][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[43][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[43][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[43][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[43][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[43][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[43][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[43][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[43][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[43][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[43][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[43][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[43][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[43][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[43][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[43][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[43][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[43][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[43][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[43][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[43][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[43][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[43][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[43][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[43][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[43][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[43][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[43][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[43][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[43][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[43][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[43][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[43][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[43][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[43][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[43][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[43][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[43][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[43][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[43][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[43][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[43][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[43][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[43][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[43][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[43][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[43][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[43][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[43][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[43][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[43][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[43][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[43][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[43][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[43][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[43][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[43][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[43][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[43][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[43][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[43][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[43][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[43][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[43][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[43][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[43][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[43][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[43][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[43][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[43][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[43][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[43][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[43][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[43][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[43][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[43][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[43][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[43][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[43][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[43][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[43][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[43][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[43][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[43][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[43][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[43][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[43][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[43][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[43][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[43][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[43][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[43][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[43][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[43][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[43][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[43][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[43][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[43][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[43][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[43][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[43][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[43][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[43][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[43][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 43, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[43][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[43][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[43][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[43][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[43].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[43][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[43][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[43].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[43][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[44][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[44][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[44][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[44][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[44][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[44][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[44][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[44][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[44][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[44][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[44][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[44][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[44][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[44][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[44][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[44][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[44][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[44][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[44][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[44][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[44][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[44][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[44][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[44][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[44][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[44][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[44][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[44][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[44][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[44][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[44][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[44][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[44][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[44][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[44][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[44][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[44][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[44][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[44][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[44][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[44][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[44][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[44][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[44][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[44][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[44][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[44][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[44][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[44][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[44][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[44][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[44][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[44][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[44][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[44][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[44][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[44][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[44][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[44][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[44][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[44][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[44][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[44][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[44][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[44][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[44][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[44][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[44][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[44][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[44][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[44][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[44][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[44][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[44][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[44][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[44][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[44][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[44][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[44][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[44][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[44][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[44][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[44][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[44][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[44][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[44][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[44][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[44][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[44][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[44][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[44][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[44][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[44][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[44][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[44][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[44][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[44][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[44][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[44][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[44][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[44][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[44][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[44][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[44][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[44][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[44][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[44][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[44][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[44][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[44][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[44][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[44][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[44][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[44][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[44][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[44][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[44][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[44][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[44][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[44][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[44][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[44][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[44][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[44][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[44][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[44][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[44][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[44][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[44][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[44][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[44][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[44][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[44][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[44][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[44][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[44][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[44][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[44][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[44][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[44][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[44][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[44][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[44][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[44][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[44][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[44][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[44][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[44][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[44][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[44][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[44][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[44][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[44][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[44][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[44][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[44][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[44][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[44][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[44][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[44][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[44][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[44][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[44][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[44][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[44][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[44][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[44][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[44][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[44][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[44][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[44][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[44][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[44][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[44][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[44][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[44][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[44][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[44][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[44][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[44][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[44][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[44][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[44][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[44][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[44][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[44][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 44, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[44][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[44][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[44][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[44][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[44].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[44][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[44][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[44].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[44][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[45][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[45][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[45][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[45][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[45][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[45][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[45][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[45][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[45][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[45][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[45][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[45][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[45][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[45][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[45][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[45][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[45][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[45][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[45][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[45][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[45][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[45][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[45][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[45][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[45][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[45][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[45][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[45][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[45][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[45][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[45][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[45][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[45][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[45][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[45][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[45][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[45][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[45][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[45][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[45][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[45][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[45][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[45][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[45][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[45][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[45][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[45][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[45][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[45][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[45][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[45][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[45][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[45][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[45][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[45][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[45][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[45][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[45][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[45][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[45][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[45][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[45][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[45][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[45][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[45][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[45][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[45][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[45][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[45][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[45][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[45][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[45][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[45][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[45][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[45][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[45][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[45][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[45][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[45][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[45][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[45][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[45][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[45][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[45][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[45][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[45][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[45][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[45][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[45][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[45][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[45][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[45][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[45][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[45][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[45][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[45][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[45][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[45][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[45][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[45][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[45][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[45][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[45][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[45][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[45][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[45][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[45][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[45][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[45][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[45][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[45][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[45][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[45][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[45][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[45][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[45][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[45][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[45][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[45][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[45][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[45][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[45][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[45][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[45][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[45][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[45][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[45][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[45][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[45][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[45][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[45][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[45][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[45][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[45][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[45][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[45][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[45][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[45][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[45][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[45][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[45][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[45][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[45][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[45][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[45][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[45][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[45][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[45][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[45][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[45][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[45][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[45][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[45][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[45][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[45][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[45][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[45][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[45][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[45][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[45][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[45][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[45][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[45][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[45][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[45][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[45][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[45][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[45][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[45][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[45][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[45][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[45][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[45][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[45][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[45][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[45][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[45][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[45][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[45][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[45][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[45][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[45][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[45][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[45][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[45][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[45][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 45, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[45][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[45][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[45][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[45][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[45].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[45][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[45][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[45].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[45][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[46][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[46][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[46][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[46][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[46][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[46][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[46][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[46][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[46][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[46][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[46][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[46][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[46][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[46][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[46][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[46][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[46][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[46][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[46][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[46][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[46][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[46][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[46][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[46][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[46][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[46][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[46][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[46][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[46][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[46][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[46][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[46][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[46][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[46][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[46][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[46][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[46][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[46][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[46][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[46][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[46][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[46][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[46][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[46][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[46][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[46][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[46][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[46][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[46][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[46][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[46][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[46][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[46][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[46][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[46][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[46][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[46][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[46][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[46][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[46][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[46][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[46][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[46][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[46][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[46][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[46][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[46][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[46][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[46][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[46][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[46][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[46][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[46][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[46][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[46][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[46][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[46][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[46][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[46][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[46][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[46][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[46][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[46][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[46][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[46][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[46][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[46][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[46][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[46][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[46][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[46][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[46][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[46][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[46][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[46][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[46][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[46][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[46][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[46][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[46][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[46][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[46][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[46][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[46][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[46][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[46][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[46][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[46][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[46][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[46][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[46][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[46][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[46][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[46][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[46][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[46][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[46][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[46][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[46][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[46][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[46][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[46][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[46][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[46][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[46][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[46][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[46][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[46][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[46][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[46][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[46][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[46][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[46][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[46][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[46][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[46][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[46][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[46][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[46][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[46][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[46][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[46][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[46][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[46][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[46][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[46][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[46][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[46][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[46][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[46][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[46][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[46][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[46][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[46][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[46][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[46][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[46][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[46][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[46][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[46][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[46][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[46][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[46][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[46][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[46][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[46][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[46][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[46][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[46][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[46][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[46][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[46][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[46][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[46][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[46][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[46][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[46][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[46][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[46][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[46][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[46][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[46][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[46][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[46][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[46][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[46][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 46, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[46][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[46][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[46][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[46][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[46].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[46][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[46][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[46].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[46][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[47][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[47][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[47][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[47][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[47][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[47][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[47][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[47][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[47][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[47][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[47][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[47][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[47][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[47][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[47][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[47][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[47][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[47][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[47][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[47][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[47][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[47][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[47][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[47][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[47][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[47][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[47][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[47][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[47][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[47][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[47][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[47][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[47][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[47][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[47][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[47][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[47][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[47][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[47][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[47][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[47][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[47][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[47][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[47][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[47][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[47][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[47][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[47][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[47][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[47][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[47][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[47][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[47][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[47][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[47][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[47][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[47][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[47][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[47][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[47][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[47][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[47][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[47][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[47][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[47][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[47][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[47][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[47][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[47][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[47][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[47][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[47][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[47][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[47][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[47][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[47][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[47][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[47][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[47][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[47][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[47][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[47][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[47][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[47][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[47][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[47][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[47][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[47][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[47][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[47][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[47][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[47][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[47][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[47][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[47][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[47][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[47][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[47][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[47][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[47][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[47][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[47][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[47][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[47][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[47][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[47][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[47][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[47][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[47][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[47][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[47][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[47][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[47][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[47][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[47][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[47][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[47][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[47][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[47][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[47][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[47][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[47][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[47][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[47][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[47][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[47][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[47][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[47][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[47][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[47][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[47][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[47][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[47][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[47][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[47][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[47][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[47][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[47][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[47][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[47][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[47][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[47][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[47][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[47][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[47][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[47][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[47][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[47][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[47][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[47][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[47][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[47][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[47][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[47][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[47][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[47][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[47][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[47][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[47][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[47][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[47][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[47][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[47][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[47][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[47][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[47][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[47][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[47][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[47][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[47][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[47][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[47][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[47][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[47][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[47][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[47][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[47][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[47][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[47][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[47][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[47][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[47][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[47][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[47][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[47][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[47][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 47, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[47][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[47][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[47][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[47][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[47].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[47][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[47][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[47].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[47][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[48][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[48][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[48][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[48][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[48][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[48][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[48][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[48][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[48][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[48][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[48][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[48][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[48][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[48][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[48][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[48][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[48][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[48][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[48][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[48][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[48][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[48][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[48][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[48][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[48][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[48][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[48][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[48][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[48][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[48][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[48][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[48][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[48][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[48][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[48][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[48][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[48][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[48][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[48][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[48][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[48][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[48][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[48][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[48][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[48][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[48][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[48][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[48][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[48][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[48][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[48][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[48][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[48][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[48][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[48][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[48][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[48][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[48][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[48][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[48][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[48][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[48][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[48][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[48][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[48][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[48][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[48][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[48][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[48][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[48][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[48][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[48][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[48][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[48][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[48][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[48][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[48][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[48][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[48][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[48][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[48][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[48][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[48][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[48][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[48][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[48][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[48][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[48][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[48][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[48][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[48][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[48][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[48][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[48][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[48][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[48][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[48][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[48][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[48][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[48][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[48][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[48][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[48][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[48][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[48][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[48][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[48][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[48][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[48][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[48][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[48][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[48][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[48][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[48][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[48][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[48][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[48][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[48][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[48][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[48][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[48][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[48][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[48][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[48][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[48][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[48][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[48][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[48][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[48][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[48][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[48][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[48][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[48][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[48][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[48][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[48][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[48][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[48][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[48][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[48][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[48][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[48][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[48][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[48][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[48][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[48][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[48][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[48][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[48][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[48][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[48][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[48][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[48][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[48][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[48][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[48][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[48][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[48][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[48][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[48][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[48][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[48][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[48][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[48][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[48][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[48][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[48][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[48][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[48][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[48][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[48][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[48][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[48][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[48][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[48][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[48][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[48][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[48][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[48][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[48][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[48][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[48][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[48][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[48][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[48][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[48][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 48, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[48][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[48][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[48][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[48][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[48].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[48][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[48][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[48].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[48][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[49][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[49][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[49][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[49][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[49][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[49][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[49][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[49][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[49][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[49][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[49][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[49][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[49][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[49][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[49][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[49][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[49][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[49][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[49][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[49][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[49][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[49][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[49][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[49][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[49][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[49][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[49][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[49][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[49][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[49][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[49][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[49][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[49][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[49][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[49][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[49][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[49][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[49][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[49][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[49][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[49][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[49][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[49][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[49][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[49][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[49][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[49][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[49][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[49][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[49][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[49][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[49][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[49][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[49][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[49][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[49][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[49][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[49][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[49][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[49][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[49][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[49][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[49][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[49][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[49][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[49][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[49][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[49][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[49][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[49][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[49][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[49][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[49][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[49][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[49][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[49][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[49][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[49][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[49][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[49][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[49][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[49][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[49][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[49][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[49][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[49][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[49][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[49][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[49][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[49][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[49][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[49][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[49][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[49][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[49][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[49][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[49][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[49][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[49][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[49][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[49][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[49][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[49][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[49][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[49][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[49][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[49][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[49][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[49][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[49][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[49][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[49][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[49][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[49][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[49][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[49][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[49][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[49][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[49][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[49][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[49][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[49][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[49][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[49][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[49][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[49][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[49][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[49][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[49][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[49][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[49][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[49][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[49][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[49][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[49][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[49][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[49][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[49][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[49][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[49][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[49][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[49][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[49][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[49][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[49][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[49][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[49][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[49][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[49][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[49][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[49][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[49][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[49][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[49][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[49][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[49][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[49][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[49][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[49][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[49][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[49][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[49][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[49][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[49][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[49][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[49][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[49][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[49][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[49][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[49][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[49][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[49][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[49][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[49][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[49][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[49][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[49][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[49][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[49][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[49][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[49][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[49][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[49][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[49][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[49][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[49][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 49, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[49][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[49][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[49][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[49][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[49].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[49][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[49][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[49].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[49][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[50][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[50][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[50][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[50][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[50][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[50][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[50][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[50][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[50][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[50][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[50][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[50][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[50][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[50][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[50][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[50][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[50][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[50][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[50][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[50][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[50][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[50][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[50][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[50][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[50][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[50][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[50][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[50][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[50][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[50][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[50][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[50][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[50][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[50][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[50][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[50][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[50][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[50][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[50][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[50][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[50][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[50][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[50][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[50][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[50][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[50][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[50][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[50][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[50][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[50][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[50][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[50][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[50][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[50][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[50][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[50][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[50][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[50][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[50][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[50][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[50][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[50][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[50][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[50][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[50][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[50][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[50][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[50][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[50][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[50][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[50][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[50][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[50][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[50][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[50][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[50][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[50][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[50][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[50][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[50][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[50][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[50][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[50][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[50][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[50][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[50][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[50][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[50][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[50][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[50][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[50][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[50][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[50][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[50][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[50][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[50][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[50][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[50][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[50][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[50][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[50][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[50][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[50][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[50][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[50][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[50][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[50][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[50][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[50][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[50][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[50][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[50][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[50][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[50][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[50][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[50][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[50][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[50][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[50][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[50][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[50][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[50][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[50][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[50][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[50][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[50][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[50][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[50][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[50][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[50][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[50][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[50][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[50][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[50][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[50][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[50][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[50][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[50][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[50][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[50][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[50][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[50][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[50][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[50][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[50][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[50][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[50][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[50][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[50][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[50][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[50][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[50][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[50][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[50][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[50][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[50][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[50][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[50][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[50][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[50][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[50][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[50][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[50][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[50][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[50][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[50][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[50][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[50][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[50][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[50][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[50][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[50][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[50][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[50][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[50][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[50][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[50][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[50][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[50][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[50][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[50][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[50][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[50][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[50][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[50][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[50][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 50, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[50][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[50][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[50][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[50][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[50].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[50][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[50][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[50].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[50][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[51][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[51][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[51][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[51][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[51][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[51][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[51][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[51][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[51][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[51][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[51][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[51][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[51][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[51][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[51][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[51][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[51][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[51][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[51][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[51][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[51][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[51][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[51][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[51][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[51][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[51][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[51][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[51][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[51][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[51][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[51][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[51][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[51][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[51][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[51][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[51][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[51][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[51][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[51][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[51][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[51][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[51][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[51][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[51][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[51][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[51][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[51][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[51][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[51][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[51][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[51][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[51][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[51][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[51][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[51][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[51][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[51][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[51][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[51][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[51][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[51][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[51][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[51][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[51][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[51][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[51][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[51][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[51][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[51][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[51][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[51][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[51][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[51][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[51][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[51][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[51][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[51][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[51][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[51][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[51][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[51][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[51][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[51][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[51][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[51][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[51][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[51][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[51][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[51][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[51][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[51][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[51][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[51][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[51][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[51][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[51][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[51][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[51][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[51][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[51][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[51][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[51][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[51][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[51][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[51][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[51][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[51][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[51][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[51][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[51][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[51][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[51][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[51][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[51][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[51][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[51][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[51][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[51][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[51][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[51][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[51][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[51][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[51][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[51][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[51][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[51][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[51][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[51][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[51][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[51][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[51][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[51][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[51][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[51][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[51][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[51][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[51][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[51][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[51][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[51][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[51][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[51][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[51][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[51][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[51][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[51][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[51][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[51][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[51][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[51][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[51][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[51][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[51][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[51][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[51][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[51][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[51][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[51][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[51][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[51][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[51][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[51][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[51][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[51][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[51][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[51][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[51][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[51][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[51][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[51][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[51][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[51][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[51][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[51][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[51][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[51][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[51][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[51][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[51][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[51][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[51][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[51][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[51][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[51][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[51][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[51][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 51, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[51][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[51][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[51][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[51][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[51].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[51][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[51][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[51].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[51][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[52][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[52][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[52][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[52][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[52][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[52][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[52][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[52][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[52][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[52][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[52][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[52][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[52][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[52][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[52][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[52][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[52][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[52][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[52][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[52][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[52][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[52][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[52][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[52][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[52][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[52][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[52][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[52][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[52][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[52][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[52][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[52][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[52][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[52][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[52][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[52][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[52][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[52][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[52][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[52][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[52][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[52][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[52][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[52][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[52][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[52][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[52][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[52][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[52][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[52][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[52][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[52][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[52][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[52][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[52][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[52][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[52][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[52][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[52][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[52][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[52][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[52][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[52][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[52][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[52][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[52][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[52][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[52][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[52][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[52][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[52][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[52][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[52][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[52][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[52][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[52][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[52][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[52][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[52][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[52][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[52][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[52][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[52][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[52][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[52][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[52][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[52][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[52][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[52][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[52][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[52][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[52][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[52][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[52][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[52][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[52][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[52][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[52][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[52][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[52][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[52][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[52][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[52][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[52][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[52][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[52][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[52][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[52][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[52][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[52][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[52][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[52][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[52][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[52][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[52][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[52][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[52][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[52][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[52][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[52][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[52][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[52][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[52][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[52][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[52][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[52][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[52][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[52][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[52][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[52][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[52][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[52][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[52][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[52][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[52][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[52][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[52][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[52][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[52][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[52][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[52][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[52][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[52][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[52][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[52][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[52][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[52][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[52][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[52][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[52][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[52][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[52][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[52][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[52][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[52][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[52][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[52][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[52][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[52][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[52][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[52][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[52][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[52][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[52][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[52][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[52][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[52][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[52][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[52][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[52][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[52][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[52][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[52][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[52][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[52][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[52][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[52][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[52][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[52][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[52][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[52][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[52][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[52][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[52][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[52][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[52][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 52, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[52][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[52][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[52][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[52][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[52].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[52][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[52][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[52].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[52][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[53][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[53][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[53][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[53][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[53][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[53][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[53][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[53][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[53][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[53][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[53][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[53][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[53][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[53][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[53][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[53][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[53][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[53][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[53][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[53][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[53][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[53][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[53][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[53][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[53][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[53][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[53][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[53][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[53][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[53][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[53][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[53][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[53][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[53][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[53][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[53][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[53][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[53][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[53][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[53][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[53][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[53][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[53][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[53][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[53][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[53][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[53][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[53][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[53][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[53][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[53][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[53][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[53][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[53][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[53][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[53][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[53][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[53][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[53][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[53][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[53][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[53][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[53][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[53][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[53][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[53][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[53][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[53][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[53][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[53][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[53][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[53][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[53][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[53][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[53][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[53][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[53][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[53][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[53][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[53][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[53][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[53][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[53][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[53][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[53][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[53][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[53][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[53][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[53][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[53][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[53][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[53][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[53][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[53][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[53][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[53][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[53][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[53][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[53][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[53][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[53][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[53][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[53][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[53][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[53][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[53][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[53][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[53][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[53][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[53][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[53][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[53][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[53][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[53][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[53][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[53][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[53][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[53][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[53][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[53][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[53][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[53][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[53][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[53][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[53][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[53][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[53][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[53][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[53][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[53][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[53][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[53][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[53][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[53][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[53][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[53][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[53][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[53][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[53][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[53][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[53][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[53][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[53][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[53][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[53][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[53][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[53][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[53][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[53][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[53][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[53][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[53][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[53][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[53][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[53][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[53][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[53][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[53][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[53][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[53][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[53][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[53][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[53][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[53][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[53][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[53][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[53][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[53][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[53][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[53][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[53][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[53][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[53][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[53][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[53][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[53][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[53][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[53][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[53][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[53][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[53][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[53][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[53][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[53][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[53][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[53][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 53, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[53][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[53][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[53][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[53][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[53].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[53][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[53][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[53].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[53][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[54][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[54][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[54][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[54][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[54][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[54][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[54][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[54][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[54][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[54][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[54][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[54][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[54][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[54][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[54][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[54][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[54][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[54][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[54][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[54][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[54][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[54][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[54][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[54][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[54][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[54][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[54][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[54][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[54][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[54][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[54][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[54][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[54][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[54][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[54][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[54][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[54][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[54][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[54][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[54][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[54][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[54][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[54][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[54][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[54][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[54][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[54][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[54][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[54][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[54][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[54][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[54][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[54][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[54][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[54][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[54][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[54][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[54][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[54][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[54][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[54][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[54][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[54][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[54][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[54][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[54][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[54][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[54][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[54][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[54][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[54][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[54][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[54][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[54][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[54][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[54][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[54][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[54][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[54][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[54][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[54][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[54][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[54][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[54][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[54][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[54][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[54][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[54][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[54][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[54][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[54][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[54][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[54][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[54][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[54][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[54][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[54][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[54][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[54][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[54][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[54][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[54][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[54][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[54][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[54][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[54][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[54][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[54][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[54][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[54][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[54][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[54][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[54][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[54][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[54][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[54][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[54][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[54][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[54][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[54][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[54][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[54][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[54][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[54][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[54][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[54][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[54][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[54][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[54][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[54][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[54][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[54][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[54][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[54][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[54][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[54][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[54][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[54][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[54][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[54][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[54][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[54][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[54][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[54][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[54][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[54][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[54][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[54][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[54][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[54][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[54][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[54][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[54][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[54][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[54][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[54][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[54][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[54][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[54][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[54][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[54][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[54][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[54][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[54][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[54][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[54][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[54][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[54][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[54][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[54][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[54][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[54][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[54][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[54][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[54][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[54][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[54][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[54][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[54][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[54][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[54][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[54][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[54][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[54][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[54][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[54][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 54, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[54][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[54][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[54][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[54][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[54].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[54][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[54][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[54].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[54][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[55][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[55][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[55][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[55][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[55][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[55][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[55][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[55][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[55][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[55][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[55][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[55][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[55][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[55][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[55][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[55][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[55][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[55][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[55][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[55][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[55][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[55][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[55][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[55][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[55][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[55][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[55][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[55][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[55][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[55][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[55][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[55][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[55][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[55][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[55][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[55][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[55][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[55][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[55][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[55][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[55][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[55][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[55][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[55][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[55][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[55][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[55][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[55][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[55][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[55][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[55][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[55][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[55][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[55][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[55][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[55][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[55][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[55][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[55][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[55][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[55][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[55][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[55][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[55][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[55][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[55][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[55][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[55][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[55][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[55][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[55][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[55][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[55][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[55][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[55][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[55][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[55][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[55][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[55][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[55][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[55][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[55][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[55][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[55][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[55][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[55][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[55][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[55][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[55][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[55][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[55][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[55][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[55][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[55][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[55][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[55][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[55][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[55][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[55][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[55][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[55][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[55][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[55][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[55][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[55][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[55][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[55][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[55][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[55][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[55][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[55][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[55][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[55][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[55][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[55][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[55][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[55][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[55][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[55][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[55][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[55][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[55][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[55][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[55][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[55][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[55][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[55][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[55][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[55][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[55][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[55][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[55][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[55][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[55][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[55][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[55][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[55][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[55][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[55][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[55][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[55][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[55][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[55][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[55][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[55][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[55][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[55][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[55][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[55][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[55][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[55][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[55][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[55][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[55][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[55][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[55][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[55][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[55][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[55][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[55][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[55][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[55][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[55][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[55][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[55][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[55][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[55][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[55][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[55][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[55][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[55][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[55][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[55][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[55][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[55][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[55][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[55][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[55][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[55][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[55][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[55][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[55][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[55][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[55][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[55][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[55][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 55, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[55][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[55][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[55][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[55][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[55].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[55][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[55][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[55].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[55][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[56][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[56][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[56][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[56][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[56][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[56][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[56][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[56][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[56][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[56][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[56][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[56][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[56][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[56][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[56][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[56][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[56][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[56][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[56][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[56][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[56][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[56][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[56][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[56][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[56][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[56][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[56][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[56][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[56][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[56][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[56][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[56][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[56][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[56][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[56][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[56][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[56][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[56][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[56][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[56][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[56][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[56][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[56][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[56][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[56][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[56][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[56][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[56][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[56][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[56][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[56][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[56][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[56][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[56][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[56][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[56][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[56][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[56][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[56][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[56][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[56][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[56][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[56][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[56][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[56][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[56][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[56][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[56][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[56][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[56][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[56][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[56][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[56][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[56][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[56][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[56][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[56][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[56][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[56][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[56][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[56][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[56][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[56][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[56][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[56][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[56][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[56][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[56][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[56][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[56][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[56][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[56][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[56][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[56][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[56][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[56][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[56][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[56][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[56][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[56][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[56][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[56][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[56][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[56][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[56][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[56][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[56][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[56][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[56][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[56][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[56][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[56][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[56][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[56][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[56][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[56][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[56][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[56][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[56][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[56][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[56][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[56][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[56][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[56][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[56][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[56][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[56][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[56][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[56][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[56][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[56][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[56][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[56][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[56][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[56][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[56][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[56][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[56][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[56][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[56][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[56][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[56][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[56][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[56][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[56][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[56][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[56][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[56][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[56][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[56][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[56][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[56][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[56][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[56][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[56][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[56][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[56][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[56][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[56][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[56][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[56][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[56][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[56][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[56][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[56][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[56][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[56][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[56][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[56][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[56][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[56][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[56][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[56][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[56][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[56][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[56][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[56][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[56][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[56][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[56][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[56][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[56][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[56][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[56][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[56][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[56][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 56, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[56][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[56][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[56][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[56][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[56].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[56][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[56][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[56].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[56][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[57][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[57][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[57][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[57][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[57][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[57][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[57][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[57][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[57][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[57][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[57][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[57][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[57][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[57][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[57][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[57][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[57][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[57][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[57][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[57][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[57][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[57][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[57][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[57][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[57][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[57][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[57][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[57][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[57][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[57][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[57][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[57][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[57][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[57][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[57][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[57][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[57][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[57][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[57][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[57][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[57][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[57][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[57][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[57][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[57][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[57][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[57][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[57][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[57][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[57][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[57][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[57][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[57][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[57][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[57][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[57][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[57][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[57][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[57][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[57][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[57][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[57][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[57][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[57][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[57][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[57][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[57][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[57][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[57][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[57][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[57][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[57][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[57][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[57][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[57][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[57][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[57][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[57][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[57][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[57][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[57][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[57][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[57][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[57][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[57][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[57][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[57][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[57][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[57][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[57][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[57][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[57][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[57][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[57][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[57][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[57][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[57][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[57][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[57][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[57][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[57][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[57][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[57][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[57][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[57][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[57][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[57][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[57][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[57][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[57][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[57][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[57][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[57][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[57][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[57][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[57][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[57][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[57][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[57][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[57][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[57][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[57][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[57][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[57][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[57][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[57][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[57][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[57][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[57][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[57][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[57][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[57][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[57][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[57][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[57][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[57][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[57][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[57][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[57][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[57][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[57][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[57][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[57][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[57][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[57][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[57][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[57][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[57][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[57][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[57][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[57][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[57][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[57][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[57][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[57][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[57][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[57][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[57][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[57][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[57][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[57][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[57][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[57][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[57][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[57][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[57][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[57][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[57][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[57][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[57][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[57][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[57][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[57][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[57][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[57][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[57][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[57][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[57][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[57][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[57][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[57][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[57][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[57][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[57][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[57][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[57][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 57, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[57][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[57][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[57][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[57][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[57].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[57][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[57][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[57].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[57][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[58][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[58][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[58][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[58][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[58][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[58][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[58][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[58][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[58][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[58][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[58][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[58][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[58][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[58][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[58][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[58][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[58][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[58][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[58][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[58][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[58][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[58][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[58][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[58][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[58][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[58][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[58][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[58][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[58][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[58][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[58][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[58][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[58][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[58][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[58][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[58][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[58][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[58][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[58][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[58][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[58][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[58][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[58][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[58][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[58][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[58][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[58][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[58][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[58][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[58][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[58][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[58][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[58][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[58][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[58][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[58][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[58][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[58][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[58][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[58][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[58][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[58][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[58][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[58][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[58][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[58][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[58][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[58][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[58][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[58][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[58][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[58][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[58][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[58][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[58][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[58][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[58][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[58][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[58][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[58][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[58][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[58][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[58][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[58][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[58][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[58][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[58][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[58][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[58][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[58][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[58][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[58][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[58][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[58][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[58][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[58][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[58][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[58][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[58][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[58][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[58][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[58][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[58][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[58][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[58][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[58][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[58][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[58][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[58][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[58][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[58][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[58][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[58][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[58][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[58][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[58][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[58][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[58][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[58][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[58][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[58][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[58][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[58][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[58][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[58][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[58][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[58][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[58][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[58][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[58][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[58][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[58][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[58][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[58][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[58][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[58][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[58][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[58][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[58][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[58][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[58][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[58][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[58][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[58][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[58][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[58][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[58][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[58][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[58][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[58][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[58][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[58][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[58][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[58][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[58][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[58][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[58][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[58][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[58][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[58][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[58][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[58][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[58][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[58][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[58][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[58][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[58][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[58][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[58][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[58][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[58][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[58][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[58][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[58][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[58][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[58][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[58][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[58][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[58][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[58][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[58][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[58][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[58][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[58][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[58][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[58][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 58, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[58][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[58][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[58][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[58][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[58].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[58][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[58][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[58].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[58][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[59][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[59][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[59][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[59][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[59][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[59][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[59][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[59][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[59][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[59][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[59][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[59][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[59][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[59][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[59][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[59][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[59][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[59][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[59][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[59][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[59][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[59][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[59][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[59][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[59][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[59][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[59][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[59][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[59][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[59][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[59][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[59][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[59][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[59][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[59][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[59][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[59][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[59][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[59][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[59][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[59][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[59][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[59][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[59][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[59][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[59][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[59][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[59][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[59][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[59][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[59][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[59][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[59][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[59][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[59][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[59][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[59][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[59][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[59][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[59][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[59][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[59][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[59][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[59][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[59][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[59][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[59][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[59][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[59][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[59][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[59][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[59][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[59][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[59][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[59][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[59][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[59][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[59][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[59][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[59][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[59][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[59][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[59][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[59][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[59][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[59][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[59][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[59][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[59][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[59][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[59][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[59][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[59][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[59][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[59][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[59][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[59][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[59][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[59][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[59][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[59][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[59][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[59][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[59][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[59][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[59][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[59][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[59][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[59][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[59][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[59][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[59][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[59][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[59][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[59][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[59][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[59][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[59][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[59][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[59][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[59][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[59][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[59][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[59][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[59][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[59][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[59][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[59][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[59][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[59][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[59][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[59][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[59][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[59][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[59][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[59][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[59][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[59][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[59][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[59][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[59][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[59][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[59][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[59][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[59][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[59][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[59][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[59][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[59][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[59][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[59][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[59][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[59][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[59][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[59][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[59][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[59][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[59][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[59][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[59][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[59][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[59][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[59][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[59][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[59][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[59][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[59][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[59][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[59][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[59][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[59][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[59][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[59][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[59][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[59][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[59][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[59][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[59][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[59][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[59][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[59][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[59][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[59][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[59][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[59][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[59][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 59, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[59][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[59][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[59][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[59][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[59].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[59][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[59][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[59].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[59][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[60][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[60][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[60][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[60][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[60][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[60][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[60][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[60][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[60][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[60][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[60][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[60][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[60][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[60][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[60][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[60][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[60][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[60][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[60][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[60][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[60][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[60][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[60][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[60][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[60][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[60][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[60][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[60][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[60][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[60][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[60][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[60][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[60][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[60][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[60][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[60][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[60][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[60][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[60][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[60][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[60][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[60][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[60][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[60][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[60][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[60][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[60][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[60][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[60][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[60][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[60][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[60][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[60][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[60][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[60][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[60][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[60][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[60][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[60][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[60][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[60][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[60][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[60][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[60][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[60][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[60][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[60][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[60][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[60][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[60][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[60][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[60][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[60][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[60][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[60][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[60][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[60][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[60][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[60][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[60][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[60][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[60][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[60][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[60][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[60][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[60][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[60][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[60][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[60][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[60][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[60][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[60][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[60][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[60][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[60][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[60][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[60][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[60][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[60][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[60][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[60][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[60][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[60][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[60][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[60][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[60][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[60][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[60][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[60][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[60][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[60][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[60][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[60][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[60][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[60][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[60][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[60][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[60][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[60][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[60][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[60][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[60][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[60][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[60][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[60][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[60][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[60][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[60][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[60][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[60][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[60][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[60][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[60][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[60][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[60][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[60][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[60][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[60][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[60][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[60][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[60][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[60][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[60][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[60][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[60][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[60][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[60][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[60][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[60][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[60][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[60][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[60][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[60][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[60][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[60][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[60][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[60][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[60][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[60][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[60][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[60][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[60][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[60][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[60][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[60][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[60][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[60][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[60][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[60][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[60][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[60][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[60][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[60][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[60][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[60][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[60][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[60][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[60][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[60][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[60][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[60][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[60][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[60][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[60][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[60][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[60][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 60, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[60][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[60][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[60][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[60][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[60].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[60][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[60][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[60].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[60][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[61][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[61][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[61][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[61][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[61][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[61][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[61][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[61][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[61][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[61][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[61][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[61][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[61][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[61][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[61][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[61][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[61][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[61][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[61][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[61][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[61][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[61][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[61][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[61][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[61][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[61][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[61][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[61][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[61][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[61][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[61][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[61][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[61][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[61][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[61][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[61][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[61][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[61][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[61][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[61][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[61][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[61][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[61][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[61][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[61][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[61][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[61][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[61][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[61][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[61][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[61][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[61][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[61][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[61][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[61][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[61][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[61][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[61][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[61][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[61][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[61][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[61][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[61][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[61][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[61][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[61][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[61][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[61][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[61][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[61][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[61][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[61][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[61][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[61][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[61][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[61][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[61][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[61][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[61][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[61][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[61][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[61][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[61][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[61][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[61][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[61][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[61][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[61][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[61][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[61][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[61][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[61][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[61][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[61][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[61][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[61][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[61][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[61][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[61][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[61][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[61][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[61][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[61][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[61][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[61][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[61][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[61][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[61][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[61][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[61][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[61][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[61][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[61][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[61][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[61][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[61][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[61][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[61][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[61][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[61][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[61][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[61][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[61][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[61][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[61][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[61][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[61][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[61][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[61][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[61][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[61][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[61][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[61][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[61][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[61][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[61][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[61][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[61][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[61][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[61][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[61][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[61][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[61][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[61][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[61][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[61][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[61][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[61][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[61][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[61][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[61][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[61][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[61][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[61][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[61][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[61][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[61][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[61][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[61][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[61][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[61][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[61][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[61][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[61][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[61][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[61][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[61][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[61][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[61][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[61][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[61][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[61][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[61][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[61][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[61][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[61][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[61][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[61][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[61][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[61][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[61][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[61][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[61][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[61][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[61][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[61][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 61, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[61][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[61][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[61][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[61][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[61].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[61][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[61][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[61].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[61][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[62][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[62][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[62][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[62][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[62][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[62][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[62][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[62][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[62][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[62][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[62][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[62][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[62][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[62][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[62][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[62][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[62][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[62][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[62][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[62][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[62][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[62][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[62][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[62][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[62][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[62][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[62][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[62][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[62][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[62][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[62][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[62][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[62][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[62][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[62][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[62][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[62][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[62][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[62][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[62][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[62][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[62][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[62][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[62][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[62][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[62][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[62][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[62][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[62][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[62][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[62][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[62][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[62][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[62][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[62][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[62][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[62][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[62][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[62][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[62][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[62][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[62][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[62][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[62][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[62][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[62][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[62][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[62][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[62][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[62][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[62][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[62][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[62][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[62][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[62][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[62][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[62][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[62][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[62][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[62][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[62][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[62][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[62][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[62][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[62][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[62][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[62][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[62][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[62][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[62][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[62][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[62][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[62][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[62][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[62][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[62][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[62][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[62][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[62][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[62][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[62][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[62][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[62][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[62][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[62][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[62][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[62][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[62][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[62][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[62][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[62][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[62][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[62][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[62][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[62][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[62][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[62][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[62][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[62][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[62][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[62][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[62][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[62][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[62][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[62][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[62][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[62][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[62][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[62][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[62][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[62][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[62][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[62][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[62][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[62][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[62][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[62][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[62][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[62][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[62][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[62][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[62][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[62][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[62][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[62][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[62][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[62][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[62][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[62][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[62][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[62][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[62][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[62][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[62][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[62][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[62][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[62][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[62][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[62][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[62][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[62][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[62][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[62][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[62][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[62][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[62][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[62][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[62][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[62][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[62][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[62][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[62][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[62][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[62][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[62][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[62][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[62][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[62][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[62][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[62][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[62][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[62][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[62][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[62][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[62][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[62][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 62, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[62][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[62][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[62][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[62][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[62].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[62][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[62][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[62].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[62][31].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 0                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][0].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane0_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane0_strm0_cntl          =   DownstreamStackBusLane[63][0].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane0_strm0_data          =   DownstreamStackBusLane[63][0].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane0_strm0_data_valid    =   DownstreamStackBusLane[63][0].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][0].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane0_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane0_strm1_cntl          =   DownstreamStackBusLane[63][0].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane0_strm1_data          =   DownstreamStackBusLane[63][0].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane0_strm1_data_valid    =   DownstreamStackBusLane[63][0].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 1                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][1].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane1_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane1_strm0_cntl          =   DownstreamStackBusLane[63][1].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane1_strm0_data          =   DownstreamStackBusLane[63][1].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane1_strm0_data_valid    =   DownstreamStackBusLane[63][1].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][1].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane1_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane1_strm1_cntl          =   DownstreamStackBusLane[63][1].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane1_strm1_data          =   DownstreamStackBusLane[63][1].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane1_strm1_data_valid    =   DownstreamStackBusLane[63][1].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 2                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][2].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane2_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane2_strm0_cntl          =   DownstreamStackBusLane[63][2].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane2_strm0_data          =   DownstreamStackBusLane[63][2].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane2_strm0_data_valid    =   DownstreamStackBusLane[63][2].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][2].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane2_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane2_strm1_cntl          =   DownstreamStackBusLane[63][2].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane2_strm1_data          =   DownstreamStackBusLane[63][2].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane2_strm1_data_valid    =   DownstreamStackBusLane[63][2].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 3                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][3].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane3_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane3_strm0_cntl          =   DownstreamStackBusLane[63][3].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane3_strm0_data          =   DownstreamStackBusLane[63][3].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane3_strm0_data_valid    =   DownstreamStackBusLane[63][3].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][3].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane3_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane3_strm1_cntl          =   DownstreamStackBusLane[63][3].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane3_strm1_data          =   DownstreamStackBusLane[63][3].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane3_strm1_data_valid    =   DownstreamStackBusLane[63][3].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 4                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][4].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane4_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane4_strm0_cntl          =   DownstreamStackBusLane[63][4].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane4_strm0_data          =   DownstreamStackBusLane[63][4].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane4_strm0_data_valid    =   DownstreamStackBusLane[63][4].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][4].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane4_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane4_strm1_cntl          =   DownstreamStackBusLane[63][4].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane4_strm1_data          =   DownstreamStackBusLane[63][4].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane4_strm1_data_valid    =   DownstreamStackBusLane[63][4].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 5                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][5].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane5_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane5_strm0_cntl          =   DownstreamStackBusLane[63][5].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane5_strm0_data          =   DownstreamStackBusLane[63][5].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane5_strm0_data_valid    =   DownstreamStackBusLane[63][5].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][5].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane5_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane5_strm1_cntl          =   DownstreamStackBusLane[63][5].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane5_strm1_data          =   DownstreamStackBusLane[63][5].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane5_strm1_data_valid    =   DownstreamStackBusLane[63][5].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 6                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][6].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane6_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane6_strm0_cntl          =   DownstreamStackBusLane[63][6].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane6_strm0_data          =   DownstreamStackBusLane[63][6].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane6_strm0_data_valid    =   DownstreamStackBusLane[63][6].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][6].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane6_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane6_strm1_cntl          =   DownstreamStackBusLane[63][6].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane6_strm1_data          =   DownstreamStackBusLane[63][6].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane6_strm1_data_valid    =   DownstreamStackBusLane[63][6].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 7                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][7].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane7_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane7_strm0_cntl          =   DownstreamStackBusLane[63][7].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane7_strm0_data          =   DownstreamStackBusLane[63][7].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane7_strm0_data_valid    =   DownstreamStackBusLane[63][7].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][7].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane7_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane7_strm1_cntl          =   DownstreamStackBusLane[63][7].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane7_strm1_data          =   DownstreamStackBusLane[63][7].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane7_strm1_data_valid    =   DownstreamStackBusLane[63][7].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 8                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][8].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane8_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane8_strm0_cntl          =   DownstreamStackBusLane[63][8].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane8_strm0_data          =   DownstreamStackBusLane[63][8].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane8_strm0_data_valid    =   DownstreamStackBusLane[63][8].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][8].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane8_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane8_strm1_cntl          =   DownstreamStackBusLane[63][8].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane8_strm1_data          =   DownstreamStackBusLane[63][8].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane8_strm1_data_valid    =   DownstreamStackBusLane[63][8].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 9                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][9].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane9_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane9_strm0_cntl          =   DownstreamStackBusLane[63][9].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane9_strm0_data          =   DownstreamStackBusLane[63][9].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane9_strm0_data_valid    =   DownstreamStackBusLane[63][9].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][9].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane9_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane9_strm1_cntl          =   DownstreamStackBusLane[63][9].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane9_strm1_data          =   DownstreamStackBusLane[63][9].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane9_strm1_data_valid    =   DownstreamStackBusLane[63][9].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 10                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][10].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane10_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane10_strm0_cntl          =   DownstreamStackBusLane[63][10].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane10_strm0_data          =   DownstreamStackBusLane[63][10].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane10_strm0_data_valid    =   DownstreamStackBusLane[63][10].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][10].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane10_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane10_strm1_cntl          =   DownstreamStackBusLane[63][10].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane10_strm1_data          =   DownstreamStackBusLane[63][10].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane10_strm1_data_valid    =   DownstreamStackBusLane[63][10].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 11                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][11].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane11_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane11_strm0_cntl          =   DownstreamStackBusLane[63][11].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane11_strm0_data          =   DownstreamStackBusLane[63][11].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane11_strm0_data_valid    =   DownstreamStackBusLane[63][11].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][11].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane11_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane11_strm1_cntl          =   DownstreamStackBusLane[63][11].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane11_strm1_data          =   DownstreamStackBusLane[63][11].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane11_strm1_data_valid    =   DownstreamStackBusLane[63][11].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 12                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][12].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane12_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane12_strm0_cntl          =   DownstreamStackBusLane[63][12].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane12_strm0_data          =   DownstreamStackBusLane[63][12].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane12_strm0_data_valid    =   DownstreamStackBusLane[63][12].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][12].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane12_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane12_strm1_cntl          =   DownstreamStackBusLane[63][12].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane12_strm1_data          =   DownstreamStackBusLane[63][12].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane12_strm1_data_valid    =   DownstreamStackBusLane[63][12].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 13                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][13].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane13_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane13_strm0_cntl          =   DownstreamStackBusLane[63][13].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane13_strm0_data          =   DownstreamStackBusLane[63][13].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane13_strm0_data_valid    =   DownstreamStackBusLane[63][13].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][13].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane13_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane13_strm1_cntl          =   DownstreamStackBusLane[63][13].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane13_strm1_data          =   DownstreamStackBusLane[63][13].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane13_strm1_data_valid    =   DownstreamStackBusLane[63][13].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 14                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][14].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane14_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane14_strm0_cntl          =   DownstreamStackBusLane[63][14].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane14_strm0_data          =   DownstreamStackBusLane[63][14].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane14_strm0_data_valid    =   DownstreamStackBusLane[63][14].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][14].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane14_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane14_strm1_cntl          =   DownstreamStackBusLane[63][14].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane14_strm1_data          =   DownstreamStackBusLane[63][14].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane14_strm1_data_valid    =   DownstreamStackBusLane[63][14].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 15                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][15].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane15_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane15_strm0_cntl          =   DownstreamStackBusLane[63][15].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane15_strm0_data          =   DownstreamStackBusLane[63][15].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane15_strm0_data_valid    =   DownstreamStackBusLane[63][15].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][15].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane15_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane15_strm1_cntl          =   DownstreamStackBusLane[63][15].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane15_strm1_data          =   DownstreamStackBusLane[63][15].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane15_strm1_data_valid    =   DownstreamStackBusLane[63][15].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 16                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][16].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane16_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane16_strm0_cntl          =   DownstreamStackBusLane[63][16].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane16_strm0_data          =   DownstreamStackBusLane[63][16].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane16_strm0_data_valid    =   DownstreamStackBusLane[63][16].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][16].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane16_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane16_strm1_cntl          =   DownstreamStackBusLane[63][16].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane16_strm1_data          =   DownstreamStackBusLane[63][16].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane16_strm1_data_valid    =   DownstreamStackBusLane[63][16].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 17                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][17].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane17_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane17_strm0_cntl          =   DownstreamStackBusLane[63][17].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane17_strm0_data          =   DownstreamStackBusLane[63][17].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane17_strm0_data_valid    =   DownstreamStackBusLane[63][17].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][17].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane17_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane17_strm1_cntl          =   DownstreamStackBusLane[63][17].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane17_strm1_data          =   DownstreamStackBusLane[63][17].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane17_strm1_data_valid    =   DownstreamStackBusLane[63][17].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 18                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][18].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane18_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane18_strm0_cntl          =   DownstreamStackBusLane[63][18].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane18_strm0_data          =   DownstreamStackBusLane[63][18].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane18_strm0_data_valid    =   DownstreamStackBusLane[63][18].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][18].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane18_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane18_strm1_cntl          =   DownstreamStackBusLane[63][18].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane18_strm1_data          =   DownstreamStackBusLane[63][18].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane18_strm1_data_valid    =   DownstreamStackBusLane[63][18].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 19                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][19].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane19_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane19_strm0_cntl          =   DownstreamStackBusLane[63][19].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane19_strm0_data          =   DownstreamStackBusLane[63][19].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane19_strm0_data_valid    =   DownstreamStackBusLane[63][19].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][19].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane19_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane19_strm1_cntl          =   DownstreamStackBusLane[63][19].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane19_strm1_data          =   DownstreamStackBusLane[63][19].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane19_strm1_data_valid    =   DownstreamStackBusLane[63][19].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 20                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][20].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane20_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane20_strm0_cntl          =   DownstreamStackBusLane[63][20].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane20_strm0_data          =   DownstreamStackBusLane[63][20].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane20_strm0_data_valid    =   DownstreamStackBusLane[63][20].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][20].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane20_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane20_strm1_cntl          =   DownstreamStackBusLane[63][20].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane20_strm1_data          =   DownstreamStackBusLane[63][20].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane20_strm1_data_valid    =   DownstreamStackBusLane[63][20].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 21                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][21].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane21_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane21_strm0_cntl          =   DownstreamStackBusLane[63][21].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane21_strm0_data          =   DownstreamStackBusLane[63][21].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane21_strm0_data_valid    =   DownstreamStackBusLane[63][21].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][21].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane21_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane21_strm1_cntl          =   DownstreamStackBusLane[63][21].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane21_strm1_data          =   DownstreamStackBusLane[63][21].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane21_strm1_data_valid    =   DownstreamStackBusLane[63][21].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 22                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][22].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane22_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane22_strm0_cntl          =   DownstreamStackBusLane[63][22].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane22_strm0_data          =   DownstreamStackBusLane[63][22].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane22_strm0_data_valid    =   DownstreamStackBusLane[63][22].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][22].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane22_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane22_strm1_cntl          =   DownstreamStackBusLane[63][22].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane22_strm1_data          =   DownstreamStackBusLane[63][22].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane22_strm1_data_valid    =   DownstreamStackBusLane[63][22].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 23                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][23].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane23_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane23_strm0_cntl          =   DownstreamStackBusLane[63][23].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane23_strm0_data          =   DownstreamStackBusLane[63][23].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane23_strm0_data_valid    =   DownstreamStackBusLane[63][23].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][23].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane23_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane23_strm1_cntl          =   DownstreamStackBusLane[63][23].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane23_strm1_data          =   DownstreamStackBusLane[63][23].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane23_strm1_data_valid    =   DownstreamStackBusLane[63][23].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 24                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][24].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane24_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane24_strm0_cntl          =   DownstreamStackBusLane[63][24].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane24_strm0_data          =   DownstreamStackBusLane[63][24].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane24_strm0_data_valid    =   DownstreamStackBusLane[63][24].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][24].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane24_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane24_strm1_cntl          =   DownstreamStackBusLane[63][24].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane24_strm1_data          =   DownstreamStackBusLane[63][24].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane24_strm1_data_valid    =   DownstreamStackBusLane[63][24].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 25                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][25].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane25_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane25_strm0_cntl          =   DownstreamStackBusLane[63][25].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane25_strm0_data          =   DownstreamStackBusLane[63][25].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane25_strm0_data_valid    =   DownstreamStackBusLane[63][25].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][25].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane25_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane25_strm1_cntl          =   DownstreamStackBusLane[63][25].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane25_strm1_data          =   DownstreamStackBusLane[63][25].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane25_strm1_data_valid    =   DownstreamStackBusLane[63][25].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 26                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][26].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane26_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane26_strm0_cntl          =   DownstreamStackBusLane[63][26].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane26_strm0_data          =   DownstreamStackBusLane[63][26].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane26_strm0_data_valid    =   DownstreamStackBusLane[63][26].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][26].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane26_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane26_strm1_cntl          =   DownstreamStackBusLane[63][26].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane26_strm1_data          =   DownstreamStackBusLane[63][26].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane26_strm1_data_valid    =   DownstreamStackBusLane[63][26].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 27                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][27].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane27_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane27_strm0_cntl          =   DownstreamStackBusLane[63][27].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane27_strm0_data          =   DownstreamStackBusLane[63][27].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane27_strm0_data_valid    =   DownstreamStackBusLane[63][27].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][27].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane27_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane27_strm1_cntl          =   DownstreamStackBusLane[63][27].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane27_strm1_data          =   DownstreamStackBusLane[63][27].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane27_strm1_data_valid    =   DownstreamStackBusLane[63][27].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 28                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][28].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane28_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane28_strm0_cntl          =   DownstreamStackBusLane[63][28].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane28_strm0_data          =   DownstreamStackBusLane[63][28].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane28_strm0_data_valid    =   DownstreamStackBusLane[63][28].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][28].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane28_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane28_strm1_cntl          =   DownstreamStackBusLane[63][28].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane28_strm1_data          =   DownstreamStackBusLane[63][28].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane28_strm1_data_valid    =   DownstreamStackBusLane[63][28].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 29                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][29].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane29_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane29_strm0_cntl          =   DownstreamStackBusLane[63][29].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane29_strm0_data          =   DownstreamStackBusLane[63][29].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane29_strm0_data_valid    =   DownstreamStackBusLane[63][29].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][29].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane29_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane29_strm1_cntl          =   DownstreamStackBusLane[63][29].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane29_strm1_data          =   DownstreamStackBusLane[63][29].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane29_strm1_data_valid    =   DownstreamStackBusLane[63][29].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 30                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][30].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane30_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane30_strm0_cntl          =   DownstreamStackBusLane[63][30].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane30_strm0_data          =   DownstreamStackBusLane[63][30].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane30_strm0_data_valid    =   DownstreamStackBusLane[63][30].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][30].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane30_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane30_strm1_cntl          =   DownstreamStackBusLane[63][30].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane30_strm1_data          =   DownstreamStackBusLane[63][30].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane30_strm1_data_valid    =   DownstreamStackBusLane[63][30].std__pe__lane_strm1_data_valid    ;      
        
        // PE 63, Lane 31                 
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][31].pe__std__lane_strm0_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane31_strm0_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane31_strm0_cntl          =   DownstreamStackBusLane[63][31].std__pe__lane_strm0_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane31_strm0_data          =   DownstreamStackBusLane[63][31].std__pe__lane_strm0_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane31_strm0_data_valid    =   DownstreamStackBusLane[63][31].std__pe__lane_strm0_data_valid    ;      
        
        //  - doesnt seem to work if you use cb_test for observed signals 
        assign DownstreamStackBusLane[63][31].pe__std__lane_strm1_ready                         =   system_inst.manager_array_inst.mgr_inst[63].std__mgr__lane31_strm1_ready ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane31_strm1_cntl          =   DownstreamStackBusLane[63][31].std__pe__lane_strm1_cntl          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane31_strm1_data          =   DownstreamStackBusLane[63][31].std__pe__lane_strm1_data          ;      
        assign system_inst.manager_array_inst.mgr_inst[63].mgr__std__lane31_strm1_data_valid    =   DownstreamStackBusLane[63][31].std__pe__lane_strm1_data_valid    ;      
        