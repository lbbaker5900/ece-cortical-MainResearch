
  assign stOp_lane[0].scntl__stOp__operation    = scntl__sdp__lane0_stOp_operation   ;
  assign stOp_lane[0].scntl__stOp__strm0_source       = scntl__sdp__lane0_strm0_stOp_source      ;
  assign stOp_lane[0].scntl__stOp__strm0_destination  = scntl__sdp__lane0_strm0_stOp_destination ;
  assign stOp_lane[0].scntl__stOp__strm1_source       = scntl__sdp__lane0_strm1_stOp_source      ;
  assign stOp_lane[0].scntl__stOp__strm1_destination  = scntl__sdp__lane0_strm1_stOp_destination ;
  assign stOp_lane[0].scntl__stOp__strm0_enable       = scntl__sdp__lane0_strm0_stOp_enable      ;
  assign sdp__scntl__lane0_strm0_stOp_ready           = stOp_lane[0].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane0_strm0_stOp_complete        = stOp_lane[0].stOp__scntl__strm0_complete ;
  assign stOp_lane[0].scntl__stOp__strm1_enable       = scntl__sdp__lane0_strm1_stOp_enable      ;
  assign sdp__scntl__lane0_strm1_stOp_ready           = stOp_lane[0].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane0_strm1_stOp_complete        = stOp_lane[0].stOp__scntl__strm1_complete ;
  assign stOp_lane[1].scntl__stOp__operation    = scntl__sdp__lane1_stOp_operation   ;
  assign stOp_lane[1].scntl__stOp__strm0_source       = scntl__sdp__lane1_strm0_stOp_source      ;
  assign stOp_lane[1].scntl__stOp__strm0_destination  = scntl__sdp__lane1_strm0_stOp_destination ;
  assign stOp_lane[1].scntl__stOp__strm1_source       = scntl__sdp__lane1_strm1_stOp_source      ;
  assign stOp_lane[1].scntl__stOp__strm1_destination  = scntl__sdp__lane1_strm1_stOp_destination ;
  assign stOp_lane[1].scntl__stOp__strm0_enable       = scntl__sdp__lane1_strm0_stOp_enable      ;
  assign sdp__scntl__lane1_strm0_stOp_ready           = stOp_lane[1].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane1_strm0_stOp_complete        = stOp_lane[1].stOp__scntl__strm0_complete ;
  assign stOp_lane[1].scntl__stOp__strm1_enable       = scntl__sdp__lane1_strm1_stOp_enable      ;
  assign sdp__scntl__lane1_strm1_stOp_ready           = stOp_lane[1].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane1_strm1_stOp_complete        = stOp_lane[1].stOp__scntl__strm1_complete ;
  assign stOp_lane[2].scntl__stOp__operation    = scntl__sdp__lane2_stOp_operation   ;
  assign stOp_lane[2].scntl__stOp__strm0_source       = scntl__sdp__lane2_strm0_stOp_source      ;
  assign stOp_lane[2].scntl__stOp__strm0_destination  = scntl__sdp__lane2_strm0_stOp_destination ;
  assign stOp_lane[2].scntl__stOp__strm1_source       = scntl__sdp__lane2_strm1_stOp_source      ;
  assign stOp_lane[2].scntl__stOp__strm1_destination  = scntl__sdp__lane2_strm1_stOp_destination ;
  assign stOp_lane[2].scntl__stOp__strm0_enable       = scntl__sdp__lane2_strm0_stOp_enable      ;
  assign sdp__scntl__lane2_strm0_stOp_ready           = stOp_lane[2].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane2_strm0_stOp_complete        = stOp_lane[2].stOp__scntl__strm0_complete ;
  assign stOp_lane[2].scntl__stOp__strm1_enable       = scntl__sdp__lane2_strm1_stOp_enable      ;
  assign sdp__scntl__lane2_strm1_stOp_ready           = stOp_lane[2].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane2_strm1_stOp_complete        = stOp_lane[2].stOp__scntl__strm1_complete ;
  assign stOp_lane[3].scntl__stOp__operation    = scntl__sdp__lane3_stOp_operation   ;
  assign stOp_lane[3].scntl__stOp__strm0_source       = scntl__sdp__lane3_strm0_stOp_source      ;
  assign stOp_lane[3].scntl__stOp__strm0_destination  = scntl__sdp__lane3_strm0_stOp_destination ;
  assign stOp_lane[3].scntl__stOp__strm1_source       = scntl__sdp__lane3_strm1_stOp_source      ;
  assign stOp_lane[3].scntl__stOp__strm1_destination  = scntl__sdp__lane3_strm1_stOp_destination ;
  assign stOp_lane[3].scntl__stOp__strm0_enable       = scntl__sdp__lane3_strm0_stOp_enable      ;
  assign sdp__scntl__lane3_strm0_stOp_ready           = stOp_lane[3].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane3_strm0_stOp_complete        = stOp_lane[3].stOp__scntl__strm0_complete ;
  assign stOp_lane[3].scntl__stOp__strm1_enable       = scntl__sdp__lane3_strm1_stOp_enable      ;
  assign sdp__scntl__lane3_strm1_stOp_ready           = stOp_lane[3].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane3_strm1_stOp_complete        = stOp_lane[3].stOp__scntl__strm1_complete ;
  assign stOp_lane[4].scntl__stOp__operation    = scntl__sdp__lane4_stOp_operation   ;
  assign stOp_lane[4].scntl__stOp__strm0_source       = scntl__sdp__lane4_strm0_stOp_source      ;
  assign stOp_lane[4].scntl__stOp__strm0_destination  = scntl__sdp__lane4_strm0_stOp_destination ;
  assign stOp_lane[4].scntl__stOp__strm1_source       = scntl__sdp__lane4_strm1_stOp_source      ;
  assign stOp_lane[4].scntl__stOp__strm1_destination  = scntl__sdp__lane4_strm1_stOp_destination ;
  assign stOp_lane[4].scntl__stOp__strm0_enable       = scntl__sdp__lane4_strm0_stOp_enable      ;
  assign sdp__scntl__lane4_strm0_stOp_ready           = stOp_lane[4].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane4_strm0_stOp_complete        = stOp_lane[4].stOp__scntl__strm0_complete ;
  assign stOp_lane[4].scntl__stOp__strm1_enable       = scntl__sdp__lane4_strm1_stOp_enable      ;
  assign sdp__scntl__lane4_strm1_stOp_ready           = stOp_lane[4].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane4_strm1_stOp_complete        = stOp_lane[4].stOp__scntl__strm1_complete ;
  assign stOp_lane[5].scntl__stOp__operation    = scntl__sdp__lane5_stOp_operation   ;
  assign stOp_lane[5].scntl__stOp__strm0_source       = scntl__sdp__lane5_strm0_stOp_source      ;
  assign stOp_lane[5].scntl__stOp__strm0_destination  = scntl__sdp__lane5_strm0_stOp_destination ;
  assign stOp_lane[5].scntl__stOp__strm1_source       = scntl__sdp__lane5_strm1_stOp_source      ;
  assign stOp_lane[5].scntl__stOp__strm1_destination  = scntl__sdp__lane5_strm1_stOp_destination ;
  assign stOp_lane[5].scntl__stOp__strm0_enable       = scntl__sdp__lane5_strm0_stOp_enable      ;
  assign sdp__scntl__lane5_strm0_stOp_ready           = stOp_lane[5].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane5_strm0_stOp_complete        = stOp_lane[5].stOp__scntl__strm0_complete ;
  assign stOp_lane[5].scntl__stOp__strm1_enable       = scntl__sdp__lane5_strm1_stOp_enable      ;
  assign sdp__scntl__lane5_strm1_stOp_ready           = stOp_lane[5].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane5_strm1_stOp_complete        = stOp_lane[5].stOp__scntl__strm1_complete ;
  assign stOp_lane[6].scntl__stOp__operation    = scntl__sdp__lane6_stOp_operation   ;
  assign stOp_lane[6].scntl__stOp__strm0_source       = scntl__sdp__lane6_strm0_stOp_source      ;
  assign stOp_lane[6].scntl__stOp__strm0_destination  = scntl__sdp__lane6_strm0_stOp_destination ;
  assign stOp_lane[6].scntl__stOp__strm1_source       = scntl__sdp__lane6_strm1_stOp_source      ;
  assign stOp_lane[6].scntl__stOp__strm1_destination  = scntl__sdp__lane6_strm1_stOp_destination ;
  assign stOp_lane[6].scntl__stOp__strm0_enable       = scntl__sdp__lane6_strm0_stOp_enable      ;
  assign sdp__scntl__lane6_strm0_stOp_ready           = stOp_lane[6].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane6_strm0_stOp_complete        = stOp_lane[6].stOp__scntl__strm0_complete ;
  assign stOp_lane[6].scntl__stOp__strm1_enable       = scntl__sdp__lane6_strm1_stOp_enable      ;
  assign sdp__scntl__lane6_strm1_stOp_ready           = stOp_lane[6].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane6_strm1_stOp_complete        = stOp_lane[6].stOp__scntl__strm1_complete ;
  assign stOp_lane[7].scntl__stOp__operation    = scntl__sdp__lane7_stOp_operation   ;
  assign stOp_lane[7].scntl__stOp__strm0_source       = scntl__sdp__lane7_strm0_stOp_source      ;
  assign stOp_lane[7].scntl__stOp__strm0_destination  = scntl__sdp__lane7_strm0_stOp_destination ;
  assign stOp_lane[7].scntl__stOp__strm1_source       = scntl__sdp__lane7_strm1_stOp_source      ;
  assign stOp_lane[7].scntl__stOp__strm1_destination  = scntl__sdp__lane7_strm1_stOp_destination ;
  assign stOp_lane[7].scntl__stOp__strm0_enable       = scntl__sdp__lane7_strm0_stOp_enable      ;
  assign sdp__scntl__lane7_strm0_stOp_ready           = stOp_lane[7].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane7_strm0_stOp_complete        = stOp_lane[7].stOp__scntl__strm0_complete ;
  assign stOp_lane[7].scntl__stOp__strm1_enable       = scntl__sdp__lane7_strm1_stOp_enable      ;
  assign sdp__scntl__lane7_strm1_stOp_ready           = stOp_lane[7].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane7_strm1_stOp_complete        = stOp_lane[7].stOp__scntl__strm1_complete ;
  assign stOp_lane[8].scntl__stOp__operation    = scntl__sdp__lane8_stOp_operation   ;
  assign stOp_lane[8].scntl__stOp__strm0_source       = scntl__sdp__lane8_strm0_stOp_source      ;
  assign stOp_lane[8].scntl__stOp__strm0_destination  = scntl__sdp__lane8_strm0_stOp_destination ;
  assign stOp_lane[8].scntl__stOp__strm1_source       = scntl__sdp__lane8_strm1_stOp_source      ;
  assign stOp_lane[8].scntl__stOp__strm1_destination  = scntl__sdp__lane8_strm1_stOp_destination ;
  assign stOp_lane[8].scntl__stOp__strm0_enable       = scntl__sdp__lane8_strm0_stOp_enable      ;
  assign sdp__scntl__lane8_strm0_stOp_ready           = stOp_lane[8].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane8_strm0_stOp_complete        = stOp_lane[8].stOp__scntl__strm0_complete ;
  assign stOp_lane[8].scntl__stOp__strm1_enable       = scntl__sdp__lane8_strm1_stOp_enable      ;
  assign sdp__scntl__lane8_strm1_stOp_ready           = stOp_lane[8].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane8_strm1_stOp_complete        = stOp_lane[8].stOp__scntl__strm1_complete ;
  assign stOp_lane[9].scntl__stOp__operation    = scntl__sdp__lane9_stOp_operation   ;
  assign stOp_lane[9].scntl__stOp__strm0_source       = scntl__sdp__lane9_strm0_stOp_source      ;
  assign stOp_lane[9].scntl__stOp__strm0_destination  = scntl__sdp__lane9_strm0_stOp_destination ;
  assign stOp_lane[9].scntl__stOp__strm1_source       = scntl__sdp__lane9_strm1_stOp_source      ;
  assign stOp_lane[9].scntl__stOp__strm1_destination  = scntl__sdp__lane9_strm1_stOp_destination ;
  assign stOp_lane[9].scntl__stOp__strm0_enable       = scntl__sdp__lane9_strm0_stOp_enable      ;
  assign sdp__scntl__lane9_strm0_stOp_ready           = stOp_lane[9].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane9_strm0_stOp_complete        = stOp_lane[9].stOp__scntl__strm0_complete ;
  assign stOp_lane[9].scntl__stOp__strm1_enable       = scntl__sdp__lane9_strm1_stOp_enable      ;
  assign sdp__scntl__lane9_strm1_stOp_ready           = stOp_lane[9].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane9_strm1_stOp_complete        = stOp_lane[9].stOp__scntl__strm1_complete ;
  assign stOp_lane[10].scntl__stOp__operation    = scntl__sdp__lane10_stOp_operation   ;
  assign stOp_lane[10].scntl__stOp__strm0_source       = scntl__sdp__lane10_strm0_stOp_source      ;
  assign stOp_lane[10].scntl__stOp__strm0_destination  = scntl__sdp__lane10_strm0_stOp_destination ;
  assign stOp_lane[10].scntl__stOp__strm1_source       = scntl__sdp__lane10_strm1_stOp_source      ;
  assign stOp_lane[10].scntl__stOp__strm1_destination  = scntl__sdp__lane10_strm1_stOp_destination ;
  assign stOp_lane[10].scntl__stOp__strm0_enable       = scntl__sdp__lane10_strm0_stOp_enable      ;
  assign sdp__scntl__lane10_strm0_stOp_ready           = stOp_lane[10].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane10_strm0_stOp_complete        = stOp_lane[10].stOp__scntl__strm0_complete ;
  assign stOp_lane[10].scntl__stOp__strm1_enable       = scntl__sdp__lane10_strm1_stOp_enable      ;
  assign sdp__scntl__lane10_strm1_stOp_ready           = stOp_lane[10].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane10_strm1_stOp_complete        = stOp_lane[10].stOp__scntl__strm1_complete ;
  assign stOp_lane[11].scntl__stOp__operation    = scntl__sdp__lane11_stOp_operation   ;
  assign stOp_lane[11].scntl__stOp__strm0_source       = scntl__sdp__lane11_strm0_stOp_source      ;
  assign stOp_lane[11].scntl__stOp__strm0_destination  = scntl__sdp__lane11_strm0_stOp_destination ;
  assign stOp_lane[11].scntl__stOp__strm1_source       = scntl__sdp__lane11_strm1_stOp_source      ;
  assign stOp_lane[11].scntl__stOp__strm1_destination  = scntl__sdp__lane11_strm1_stOp_destination ;
  assign stOp_lane[11].scntl__stOp__strm0_enable       = scntl__sdp__lane11_strm0_stOp_enable      ;
  assign sdp__scntl__lane11_strm0_stOp_ready           = stOp_lane[11].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane11_strm0_stOp_complete        = stOp_lane[11].stOp__scntl__strm0_complete ;
  assign stOp_lane[11].scntl__stOp__strm1_enable       = scntl__sdp__lane11_strm1_stOp_enable      ;
  assign sdp__scntl__lane11_strm1_stOp_ready           = stOp_lane[11].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane11_strm1_stOp_complete        = stOp_lane[11].stOp__scntl__strm1_complete ;
  assign stOp_lane[12].scntl__stOp__operation    = scntl__sdp__lane12_stOp_operation   ;
  assign stOp_lane[12].scntl__stOp__strm0_source       = scntl__sdp__lane12_strm0_stOp_source      ;
  assign stOp_lane[12].scntl__stOp__strm0_destination  = scntl__sdp__lane12_strm0_stOp_destination ;
  assign stOp_lane[12].scntl__stOp__strm1_source       = scntl__sdp__lane12_strm1_stOp_source      ;
  assign stOp_lane[12].scntl__stOp__strm1_destination  = scntl__sdp__lane12_strm1_stOp_destination ;
  assign stOp_lane[12].scntl__stOp__strm0_enable       = scntl__sdp__lane12_strm0_stOp_enable      ;
  assign sdp__scntl__lane12_strm0_stOp_ready           = stOp_lane[12].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane12_strm0_stOp_complete        = stOp_lane[12].stOp__scntl__strm0_complete ;
  assign stOp_lane[12].scntl__stOp__strm1_enable       = scntl__sdp__lane12_strm1_stOp_enable      ;
  assign sdp__scntl__lane12_strm1_stOp_ready           = stOp_lane[12].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane12_strm1_stOp_complete        = stOp_lane[12].stOp__scntl__strm1_complete ;
  assign stOp_lane[13].scntl__stOp__operation    = scntl__sdp__lane13_stOp_operation   ;
  assign stOp_lane[13].scntl__stOp__strm0_source       = scntl__sdp__lane13_strm0_stOp_source      ;
  assign stOp_lane[13].scntl__stOp__strm0_destination  = scntl__sdp__lane13_strm0_stOp_destination ;
  assign stOp_lane[13].scntl__stOp__strm1_source       = scntl__sdp__lane13_strm1_stOp_source      ;
  assign stOp_lane[13].scntl__stOp__strm1_destination  = scntl__sdp__lane13_strm1_stOp_destination ;
  assign stOp_lane[13].scntl__stOp__strm0_enable       = scntl__sdp__lane13_strm0_stOp_enable      ;
  assign sdp__scntl__lane13_strm0_stOp_ready           = stOp_lane[13].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane13_strm0_stOp_complete        = stOp_lane[13].stOp__scntl__strm0_complete ;
  assign stOp_lane[13].scntl__stOp__strm1_enable       = scntl__sdp__lane13_strm1_stOp_enable      ;
  assign sdp__scntl__lane13_strm1_stOp_ready           = stOp_lane[13].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane13_strm1_stOp_complete        = stOp_lane[13].stOp__scntl__strm1_complete ;
  assign stOp_lane[14].scntl__stOp__operation    = scntl__sdp__lane14_stOp_operation   ;
  assign stOp_lane[14].scntl__stOp__strm0_source       = scntl__sdp__lane14_strm0_stOp_source      ;
  assign stOp_lane[14].scntl__stOp__strm0_destination  = scntl__sdp__lane14_strm0_stOp_destination ;
  assign stOp_lane[14].scntl__stOp__strm1_source       = scntl__sdp__lane14_strm1_stOp_source      ;
  assign stOp_lane[14].scntl__stOp__strm1_destination  = scntl__sdp__lane14_strm1_stOp_destination ;
  assign stOp_lane[14].scntl__stOp__strm0_enable       = scntl__sdp__lane14_strm0_stOp_enable      ;
  assign sdp__scntl__lane14_strm0_stOp_ready           = stOp_lane[14].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane14_strm0_stOp_complete        = stOp_lane[14].stOp__scntl__strm0_complete ;
  assign stOp_lane[14].scntl__stOp__strm1_enable       = scntl__sdp__lane14_strm1_stOp_enable      ;
  assign sdp__scntl__lane14_strm1_stOp_ready           = stOp_lane[14].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane14_strm1_stOp_complete        = stOp_lane[14].stOp__scntl__strm1_complete ;
  assign stOp_lane[15].scntl__stOp__operation    = scntl__sdp__lane15_stOp_operation   ;
  assign stOp_lane[15].scntl__stOp__strm0_source       = scntl__sdp__lane15_strm0_stOp_source      ;
  assign stOp_lane[15].scntl__stOp__strm0_destination  = scntl__sdp__lane15_strm0_stOp_destination ;
  assign stOp_lane[15].scntl__stOp__strm1_source       = scntl__sdp__lane15_strm1_stOp_source      ;
  assign stOp_lane[15].scntl__stOp__strm1_destination  = scntl__sdp__lane15_strm1_stOp_destination ;
  assign stOp_lane[15].scntl__stOp__strm0_enable       = scntl__sdp__lane15_strm0_stOp_enable      ;
  assign sdp__scntl__lane15_strm0_stOp_ready           = stOp_lane[15].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane15_strm0_stOp_complete        = stOp_lane[15].stOp__scntl__strm0_complete ;
  assign stOp_lane[15].scntl__stOp__strm1_enable       = scntl__sdp__lane15_strm1_stOp_enable      ;
  assign sdp__scntl__lane15_strm1_stOp_ready           = stOp_lane[15].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane15_strm1_stOp_complete        = stOp_lane[15].stOp__scntl__strm1_complete ;
  assign stOp_lane[16].scntl__stOp__operation    = scntl__sdp__lane16_stOp_operation   ;
  assign stOp_lane[16].scntl__stOp__strm0_source       = scntl__sdp__lane16_strm0_stOp_source      ;
  assign stOp_lane[16].scntl__stOp__strm0_destination  = scntl__sdp__lane16_strm0_stOp_destination ;
  assign stOp_lane[16].scntl__stOp__strm1_source       = scntl__sdp__lane16_strm1_stOp_source      ;
  assign stOp_lane[16].scntl__stOp__strm1_destination  = scntl__sdp__lane16_strm1_stOp_destination ;
  assign stOp_lane[16].scntl__stOp__strm0_enable       = scntl__sdp__lane16_strm0_stOp_enable      ;
  assign sdp__scntl__lane16_strm0_stOp_ready           = stOp_lane[16].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane16_strm0_stOp_complete        = stOp_lane[16].stOp__scntl__strm0_complete ;
  assign stOp_lane[16].scntl__stOp__strm1_enable       = scntl__sdp__lane16_strm1_stOp_enable      ;
  assign sdp__scntl__lane16_strm1_stOp_ready           = stOp_lane[16].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane16_strm1_stOp_complete        = stOp_lane[16].stOp__scntl__strm1_complete ;
  assign stOp_lane[17].scntl__stOp__operation    = scntl__sdp__lane17_stOp_operation   ;
  assign stOp_lane[17].scntl__stOp__strm0_source       = scntl__sdp__lane17_strm0_stOp_source      ;
  assign stOp_lane[17].scntl__stOp__strm0_destination  = scntl__sdp__lane17_strm0_stOp_destination ;
  assign stOp_lane[17].scntl__stOp__strm1_source       = scntl__sdp__lane17_strm1_stOp_source      ;
  assign stOp_lane[17].scntl__stOp__strm1_destination  = scntl__sdp__lane17_strm1_stOp_destination ;
  assign stOp_lane[17].scntl__stOp__strm0_enable       = scntl__sdp__lane17_strm0_stOp_enable      ;
  assign sdp__scntl__lane17_strm0_stOp_ready           = stOp_lane[17].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane17_strm0_stOp_complete        = stOp_lane[17].stOp__scntl__strm0_complete ;
  assign stOp_lane[17].scntl__stOp__strm1_enable       = scntl__sdp__lane17_strm1_stOp_enable      ;
  assign sdp__scntl__lane17_strm1_stOp_ready           = stOp_lane[17].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane17_strm1_stOp_complete        = stOp_lane[17].stOp__scntl__strm1_complete ;
  assign stOp_lane[18].scntl__stOp__operation    = scntl__sdp__lane18_stOp_operation   ;
  assign stOp_lane[18].scntl__stOp__strm0_source       = scntl__sdp__lane18_strm0_stOp_source      ;
  assign stOp_lane[18].scntl__stOp__strm0_destination  = scntl__sdp__lane18_strm0_stOp_destination ;
  assign stOp_lane[18].scntl__stOp__strm1_source       = scntl__sdp__lane18_strm1_stOp_source      ;
  assign stOp_lane[18].scntl__stOp__strm1_destination  = scntl__sdp__lane18_strm1_stOp_destination ;
  assign stOp_lane[18].scntl__stOp__strm0_enable       = scntl__sdp__lane18_strm0_stOp_enable      ;
  assign sdp__scntl__lane18_strm0_stOp_ready           = stOp_lane[18].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane18_strm0_stOp_complete        = stOp_lane[18].stOp__scntl__strm0_complete ;
  assign stOp_lane[18].scntl__stOp__strm1_enable       = scntl__sdp__lane18_strm1_stOp_enable      ;
  assign sdp__scntl__lane18_strm1_stOp_ready           = stOp_lane[18].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane18_strm1_stOp_complete        = stOp_lane[18].stOp__scntl__strm1_complete ;
  assign stOp_lane[19].scntl__stOp__operation    = scntl__sdp__lane19_stOp_operation   ;
  assign stOp_lane[19].scntl__stOp__strm0_source       = scntl__sdp__lane19_strm0_stOp_source      ;
  assign stOp_lane[19].scntl__stOp__strm0_destination  = scntl__sdp__lane19_strm0_stOp_destination ;
  assign stOp_lane[19].scntl__stOp__strm1_source       = scntl__sdp__lane19_strm1_stOp_source      ;
  assign stOp_lane[19].scntl__stOp__strm1_destination  = scntl__sdp__lane19_strm1_stOp_destination ;
  assign stOp_lane[19].scntl__stOp__strm0_enable       = scntl__sdp__lane19_strm0_stOp_enable      ;
  assign sdp__scntl__lane19_strm0_stOp_ready           = stOp_lane[19].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane19_strm0_stOp_complete        = stOp_lane[19].stOp__scntl__strm0_complete ;
  assign stOp_lane[19].scntl__stOp__strm1_enable       = scntl__sdp__lane19_strm1_stOp_enable      ;
  assign sdp__scntl__lane19_strm1_stOp_ready           = stOp_lane[19].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane19_strm1_stOp_complete        = stOp_lane[19].stOp__scntl__strm1_complete ;
  assign stOp_lane[20].scntl__stOp__operation    = scntl__sdp__lane20_stOp_operation   ;
  assign stOp_lane[20].scntl__stOp__strm0_source       = scntl__sdp__lane20_strm0_stOp_source      ;
  assign stOp_lane[20].scntl__stOp__strm0_destination  = scntl__sdp__lane20_strm0_stOp_destination ;
  assign stOp_lane[20].scntl__stOp__strm1_source       = scntl__sdp__lane20_strm1_stOp_source      ;
  assign stOp_lane[20].scntl__stOp__strm1_destination  = scntl__sdp__lane20_strm1_stOp_destination ;
  assign stOp_lane[20].scntl__stOp__strm0_enable       = scntl__sdp__lane20_strm0_stOp_enable      ;
  assign sdp__scntl__lane20_strm0_stOp_ready           = stOp_lane[20].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane20_strm0_stOp_complete        = stOp_lane[20].stOp__scntl__strm0_complete ;
  assign stOp_lane[20].scntl__stOp__strm1_enable       = scntl__sdp__lane20_strm1_stOp_enable      ;
  assign sdp__scntl__lane20_strm1_stOp_ready           = stOp_lane[20].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane20_strm1_stOp_complete        = stOp_lane[20].stOp__scntl__strm1_complete ;
  assign stOp_lane[21].scntl__stOp__operation    = scntl__sdp__lane21_stOp_operation   ;
  assign stOp_lane[21].scntl__stOp__strm0_source       = scntl__sdp__lane21_strm0_stOp_source      ;
  assign stOp_lane[21].scntl__stOp__strm0_destination  = scntl__sdp__lane21_strm0_stOp_destination ;
  assign stOp_lane[21].scntl__stOp__strm1_source       = scntl__sdp__lane21_strm1_stOp_source      ;
  assign stOp_lane[21].scntl__stOp__strm1_destination  = scntl__sdp__lane21_strm1_stOp_destination ;
  assign stOp_lane[21].scntl__stOp__strm0_enable       = scntl__sdp__lane21_strm0_stOp_enable      ;
  assign sdp__scntl__lane21_strm0_stOp_ready           = stOp_lane[21].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane21_strm0_stOp_complete        = stOp_lane[21].stOp__scntl__strm0_complete ;
  assign stOp_lane[21].scntl__stOp__strm1_enable       = scntl__sdp__lane21_strm1_stOp_enable      ;
  assign sdp__scntl__lane21_strm1_stOp_ready           = stOp_lane[21].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane21_strm1_stOp_complete        = stOp_lane[21].stOp__scntl__strm1_complete ;
  assign stOp_lane[22].scntl__stOp__operation    = scntl__sdp__lane22_stOp_operation   ;
  assign stOp_lane[22].scntl__stOp__strm0_source       = scntl__sdp__lane22_strm0_stOp_source      ;
  assign stOp_lane[22].scntl__stOp__strm0_destination  = scntl__sdp__lane22_strm0_stOp_destination ;
  assign stOp_lane[22].scntl__stOp__strm1_source       = scntl__sdp__lane22_strm1_stOp_source      ;
  assign stOp_lane[22].scntl__stOp__strm1_destination  = scntl__sdp__lane22_strm1_stOp_destination ;
  assign stOp_lane[22].scntl__stOp__strm0_enable       = scntl__sdp__lane22_strm0_stOp_enable      ;
  assign sdp__scntl__lane22_strm0_stOp_ready           = stOp_lane[22].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane22_strm0_stOp_complete        = stOp_lane[22].stOp__scntl__strm0_complete ;
  assign stOp_lane[22].scntl__stOp__strm1_enable       = scntl__sdp__lane22_strm1_stOp_enable      ;
  assign sdp__scntl__lane22_strm1_stOp_ready           = stOp_lane[22].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane22_strm1_stOp_complete        = stOp_lane[22].stOp__scntl__strm1_complete ;
  assign stOp_lane[23].scntl__stOp__operation    = scntl__sdp__lane23_stOp_operation   ;
  assign stOp_lane[23].scntl__stOp__strm0_source       = scntl__sdp__lane23_strm0_stOp_source      ;
  assign stOp_lane[23].scntl__stOp__strm0_destination  = scntl__sdp__lane23_strm0_stOp_destination ;
  assign stOp_lane[23].scntl__stOp__strm1_source       = scntl__sdp__lane23_strm1_stOp_source      ;
  assign stOp_lane[23].scntl__stOp__strm1_destination  = scntl__sdp__lane23_strm1_stOp_destination ;
  assign stOp_lane[23].scntl__stOp__strm0_enable       = scntl__sdp__lane23_strm0_stOp_enable      ;
  assign sdp__scntl__lane23_strm0_stOp_ready           = stOp_lane[23].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane23_strm0_stOp_complete        = stOp_lane[23].stOp__scntl__strm0_complete ;
  assign stOp_lane[23].scntl__stOp__strm1_enable       = scntl__sdp__lane23_strm1_stOp_enable      ;
  assign sdp__scntl__lane23_strm1_stOp_ready           = stOp_lane[23].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane23_strm1_stOp_complete        = stOp_lane[23].stOp__scntl__strm1_complete ;
  assign stOp_lane[24].scntl__stOp__operation    = scntl__sdp__lane24_stOp_operation   ;
  assign stOp_lane[24].scntl__stOp__strm0_source       = scntl__sdp__lane24_strm0_stOp_source      ;
  assign stOp_lane[24].scntl__stOp__strm0_destination  = scntl__sdp__lane24_strm0_stOp_destination ;
  assign stOp_lane[24].scntl__stOp__strm1_source       = scntl__sdp__lane24_strm1_stOp_source      ;
  assign stOp_lane[24].scntl__stOp__strm1_destination  = scntl__sdp__lane24_strm1_stOp_destination ;
  assign stOp_lane[24].scntl__stOp__strm0_enable       = scntl__sdp__lane24_strm0_stOp_enable      ;
  assign sdp__scntl__lane24_strm0_stOp_ready           = stOp_lane[24].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane24_strm0_stOp_complete        = stOp_lane[24].stOp__scntl__strm0_complete ;
  assign stOp_lane[24].scntl__stOp__strm1_enable       = scntl__sdp__lane24_strm1_stOp_enable      ;
  assign sdp__scntl__lane24_strm1_stOp_ready           = stOp_lane[24].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane24_strm1_stOp_complete        = stOp_lane[24].stOp__scntl__strm1_complete ;
  assign stOp_lane[25].scntl__stOp__operation    = scntl__sdp__lane25_stOp_operation   ;
  assign stOp_lane[25].scntl__stOp__strm0_source       = scntl__sdp__lane25_strm0_stOp_source      ;
  assign stOp_lane[25].scntl__stOp__strm0_destination  = scntl__sdp__lane25_strm0_stOp_destination ;
  assign stOp_lane[25].scntl__stOp__strm1_source       = scntl__sdp__lane25_strm1_stOp_source      ;
  assign stOp_lane[25].scntl__stOp__strm1_destination  = scntl__sdp__lane25_strm1_stOp_destination ;
  assign stOp_lane[25].scntl__stOp__strm0_enable       = scntl__sdp__lane25_strm0_stOp_enable      ;
  assign sdp__scntl__lane25_strm0_stOp_ready           = stOp_lane[25].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane25_strm0_stOp_complete        = stOp_lane[25].stOp__scntl__strm0_complete ;
  assign stOp_lane[25].scntl__stOp__strm1_enable       = scntl__sdp__lane25_strm1_stOp_enable      ;
  assign sdp__scntl__lane25_strm1_stOp_ready           = stOp_lane[25].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane25_strm1_stOp_complete        = stOp_lane[25].stOp__scntl__strm1_complete ;
  assign stOp_lane[26].scntl__stOp__operation    = scntl__sdp__lane26_stOp_operation   ;
  assign stOp_lane[26].scntl__stOp__strm0_source       = scntl__sdp__lane26_strm0_stOp_source      ;
  assign stOp_lane[26].scntl__stOp__strm0_destination  = scntl__sdp__lane26_strm0_stOp_destination ;
  assign stOp_lane[26].scntl__stOp__strm1_source       = scntl__sdp__lane26_strm1_stOp_source      ;
  assign stOp_lane[26].scntl__stOp__strm1_destination  = scntl__sdp__lane26_strm1_stOp_destination ;
  assign stOp_lane[26].scntl__stOp__strm0_enable       = scntl__sdp__lane26_strm0_stOp_enable      ;
  assign sdp__scntl__lane26_strm0_stOp_ready           = stOp_lane[26].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane26_strm0_stOp_complete        = stOp_lane[26].stOp__scntl__strm0_complete ;
  assign stOp_lane[26].scntl__stOp__strm1_enable       = scntl__sdp__lane26_strm1_stOp_enable      ;
  assign sdp__scntl__lane26_strm1_stOp_ready           = stOp_lane[26].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane26_strm1_stOp_complete        = stOp_lane[26].stOp__scntl__strm1_complete ;
  assign stOp_lane[27].scntl__stOp__operation    = scntl__sdp__lane27_stOp_operation   ;
  assign stOp_lane[27].scntl__stOp__strm0_source       = scntl__sdp__lane27_strm0_stOp_source      ;
  assign stOp_lane[27].scntl__stOp__strm0_destination  = scntl__sdp__lane27_strm0_stOp_destination ;
  assign stOp_lane[27].scntl__stOp__strm1_source       = scntl__sdp__lane27_strm1_stOp_source      ;
  assign stOp_lane[27].scntl__stOp__strm1_destination  = scntl__sdp__lane27_strm1_stOp_destination ;
  assign stOp_lane[27].scntl__stOp__strm0_enable       = scntl__sdp__lane27_strm0_stOp_enable      ;
  assign sdp__scntl__lane27_strm0_stOp_ready           = stOp_lane[27].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane27_strm0_stOp_complete        = stOp_lane[27].stOp__scntl__strm0_complete ;
  assign stOp_lane[27].scntl__stOp__strm1_enable       = scntl__sdp__lane27_strm1_stOp_enable      ;
  assign sdp__scntl__lane27_strm1_stOp_ready           = stOp_lane[27].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane27_strm1_stOp_complete        = stOp_lane[27].stOp__scntl__strm1_complete ;
  assign stOp_lane[28].scntl__stOp__operation    = scntl__sdp__lane28_stOp_operation   ;
  assign stOp_lane[28].scntl__stOp__strm0_source       = scntl__sdp__lane28_strm0_stOp_source      ;
  assign stOp_lane[28].scntl__stOp__strm0_destination  = scntl__sdp__lane28_strm0_stOp_destination ;
  assign stOp_lane[28].scntl__stOp__strm1_source       = scntl__sdp__lane28_strm1_stOp_source      ;
  assign stOp_lane[28].scntl__stOp__strm1_destination  = scntl__sdp__lane28_strm1_stOp_destination ;
  assign stOp_lane[28].scntl__stOp__strm0_enable       = scntl__sdp__lane28_strm0_stOp_enable      ;
  assign sdp__scntl__lane28_strm0_stOp_ready           = stOp_lane[28].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane28_strm0_stOp_complete        = stOp_lane[28].stOp__scntl__strm0_complete ;
  assign stOp_lane[28].scntl__stOp__strm1_enable       = scntl__sdp__lane28_strm1_stOp_enable      ;
  assign sdp__scntl__lane28_strm1_stOp_ready           = stOp_lane[28].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane28_strm1_stOp_complete        = stOp_lane[28].stOp__scntl__strm1_complete ;
  assign stOp_lane[29].scntl__stOp__operation    = scntl__sdp__lane29_stOp_operation   ;
  assign stOp_lane[29].scntl__stOp__strm0_source       = scntl__sdp__lane29_strm0_stOp_source      ;
  assign stOp_lane[29].scntl__stOp__strm0_destination  = scntl__sdp__lane29_strm0_stOp_destination ;
  assign stOp_lane[29].scntl__stOp__strm1_source       = scntl__sdp__lane29_strm1_stOp_source      ;
  assign stOp_lane[29].scntl__stOp__strm1_destination  = scntl__sdp__lane29_strm1_stOp_destination ;
  assign stOp_lane[29].scntl__stOp__strm0_enable       = scntl__sdp__lane29_strm0_stOp_enable      ;
  assign sdp__scntl__lane29_strm0_stOp_ready           = stOp_lane[29].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane29_strm0_stOp_complete        = stOp_lane[29].stOp__scntl__strm0_complete ;
  assign stOp_lane[29].scntl__stOp__strm1_enable       = scntl__sdp__lane29_strm1_stOp_enable      ;
  assign sdp__scntl__lane29_strm1_stOp_ready           = stOp_lane[29].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane29_strm1_stOp_complete        = stOp_lane[29].stOp__scntl__strm1_complete ;
  assign stOp_lane[30].scntl__stOp__operation    = scntl__sdp__lane30_stOp_operation   ;
  assign stOp_lane[30].scntl__stOp__strm0_source       = scntl__sdp__lane30_strm0_stOp_source      ;
  assign stOp_lane[30].scntl__stOp__strm0_destination  = scntl__sdp__lane30_strm0_stOp_destination ;
  assign stOp_lane[30].scntl__stOp__strm1_source       = scntl__sdp__lane30_strm1_stOp_source      ;
  assign stOp_lane[30].scntl__stOp__strm1_destination  = scntl__sdp__lane30_strm1_stOp_destination ;
  assign stOp_lane[30].scntl__stOp__strm0_enable       = scntl__sdp__lane30_strm0_stOp_enable      ;
  assign sdp__scntl__lane30_strm0_stOp_ready           = stOp_lane[30].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane30_strm0_stOp_complete        = stOp_lane[30].stOp__scntl__strm0_complete ;
  assign stOp_lane[30].scntl__stOp__strm1_enable       = scntl__sdp__lane30_strm1_stOp_enable      ;
  assign sdp__scntl__lane30_strm1_stOp_ready           = stOp_lane[30].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane30_strm1_stOp_complete        = stOp_lane[30].stOp__scntl__strm1_complete ;
  assign stOp_lane[31].scntl__stOp__operation    = scntl__sdp__lane31_stOp_operation   ;
  assign stOp_lane[31].scntl__stOp__strm0_source       = scntl__sdp__lane31_strm0_stOp_source      ;
  assign stOp_lane[31].scntl__stOp__strm0_destination  = scntl__sdp__lane31_strm0_stOp_destination ;
  assign stOp_lane[31].scntl__stOp__strm1_source       = scntl__sdp__lane31_strm1_stOp_source      ;
  assign stOp_lane[31].scntl__stOp__strm1_destination  = scntl__sdp__lane31_strm1_stOp_destination ;
  assign stOp_lane[31].scntl__stOp__strm0_enable       = scntl__sdp__lane31_strm0_stOp_enable      ;
  assign sdp__scntl__lane31_strm0_stOp_ready           = stOp_lane[31].stOp__scntl__strm0_ready    ;
  assign sdp__scntl__lane31_strm0_stOp_complete        = stOp_lane[31].stOp__scntl__strm0_complete ;
  assign stOp_lane[31].scntl__stOp__strm1_enable       = scntl__sdp__lane31_strm1_stOp_enable      ;
  assign sdp__scntl__lane31_strm1_stOp_ready           = stOp_lane[31].stOp__scntl__strm1_ready    ;
  assign sdp__scntl__lane31_strm1_stOp_complete        = stOp_lane[31].stOp__scntl__strm1_complete ;
