
            begin
                @vDownstreamStackBusLane[0][0].cb_test                                      ;
                vDownstreamStackBusLane [0][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][1].cb_test                                      ;
                vDownstreamStackBusLane [0][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][2].cb_test                                      ;
                vDownstreamStackBusLane [0][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][3].cb_test                                      ;
                vDownstreamStackBusLane [0][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][4].cb_test                                      ;
                vDownstreamStackBusLane [0][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][5].cb_test                                      ;
                vDownstreamStackBusLane [0][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][6].cb_test                                      ;
                vDownstreamStackBusLane [0][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][7].cb_test                                      ;
                vDownstreamStackBusLane [0][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][8].cb_test                                      ;
                vDownstreamStackBusLane [0][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][9].cb_test                                      ;
                vDownstreamStackBusLane [0][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][10].cb_test                                      ;
                vDownstreamStackBusLane [0][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][11].cb_test                                      ;
                vDownstreamStackBusLane [0][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][12].cb_test                                      ;
                vDownstreamStackBusLane [0][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][13].cb_test                                      ;
                vDownstreamStackBusLane [0][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][14].cb_test                                      ;
                vDownstreamStackBusLane [0][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][15].cb_test                                      ;
                vDownstreamStackBusLane [0][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][16].cb_test                                      ;
                vDownstreamStackBusLane [0][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][17].cb_test                                      ;
                vDownstreamStackBusLane [0][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][18].cb_test                                      ;
                vDownstreamStackBusLane [0][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][19].cb_test                                      ;
                vDownstreamStackBusLane [0][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][20].cb_test                                      ;
                vDownstreamStackBusLane [0][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][21].cb_test                                      ;
                vDownstreamStackBusLane [0][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][22].cb_test                                      ;
                vDownstreamStackBusLane [0][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][23].cb_test                                      ;
                vDownstreamStackBusLane [0][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][24].cb_test                                      ;
                vDownstreamStackBusLane [0][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][25].cb_test                                      ;
                vDownstreamStackBusLane [0][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][26].cb_test                                      ;
                vDownstreamStackBusLane [0][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][27].cb_test                                      ;
                vDownstreamStackBusLane [0][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][28].cb_test                                      ;
                vDownstreamStackBusLane [0][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][29].cb_test                                      ;
                vDownstreamStackBusLane [0][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][30].cb_test                                      ;
                vDownstreamStackBusLane [0][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[0][31].cb_test                                      ;
                vDownstreamStackBusLane [0][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [0][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[1][0].cb_test                                      ;
                vDownstreamStackBusLane [1][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][1].cb_test                                      ;
                vDownstreamStackBusLane [1][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][2].cb_test                                      ;
                vDownstreamStackBusLane [1][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][3].cb_test                                      ;
                vDownstreamStackBusLane [1][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][4].cb_test                                      ;
                vDownstreamStackBusLane [1][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][5].cb_test                                      ;
                vDownstreamStackBusLane [1][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][6].cb_test                                      ;
                vDownstreamStackBusLane [1][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][7].cb_test                                      ;
                vDownstreamStackBusLane [1][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][8].cb_test                                      ;
                vDownstreamStackBusLane [1][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][9].cb_test                                      ;
                vDownstreamStackBusLane [1][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][10].cb_test                                      ;
                vDownstreamStackBusLane [1][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][11].cb_test                                      ;
                vDownstreamStackBusLane [1][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][12].cb_test                                      ;
                vDownstreamStackBusLane [1][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][13].cb_test                                      ;
                vDownstreamStackBusLane [1][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][14].cb_test                                      ;
                vDownstreamStackBusLane [1][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][15].cb_test                                      ;
                vDownstreamStackBusLane [1][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][16].cb_test                                      ;
                vDownstreamStackBusLane [1][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][17].cb_test                                      ;
                vDownstreamStackBusLane [1][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][18].cb_test                                      ;
                vDownstreamStackBusLane [1][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][19].cb_test                                      ;
                vDownstreamStackBusLane [1][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][20].cb_test                                      ;
                vDownstreamStackBusLane [1][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][21].cb_test                                      ;
                vDownstreamStackBusLane [1][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][22].cb_test                                      ;
                vDownstreamStackBusLane [1][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][23].cb_test                                      ;
                vDownstreamStackBusLane [1][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][24].cb_test                                      ;
                vDownstreamStackBusLane [1][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][25].cb_test                                      ;
                vDownstreamStackBusLane [1][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][26].cb_test                                      ;
                vDownstreamStackBusLane [1][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][27].cb_test                                      ;
                vDownstreamStackBusLane [1][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][28].cb_test                                      ;
                vDownstreamStackBusLane [1][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][29].cb_test                                      ;
                vDownstreamStackBusLane [1][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][30].cb_test                                      ;
                vDownstreamStackBusLane [1][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[1][31].cb_test                                      ;
                vDownstreamStackBusLane [1][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [1][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[2][0].cb_test                                      ;
                vDownstreamStackBusLane [2][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][1].cb_test                                      ;
                vDownstreamStackBusLane [2][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][2].cb_test                                      ;
                vDownstreamStackBusLane [2][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][3].cb_test                                      ;
                vDownstreamStackBusLane [2][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][4].cb_test                                      ;
                vDownstreamStackBusLane [2][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][5].cb_test                                      ;
                vDownstreamStackBusLane [2][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][6].cb_test                                      ;
                vDownstreamStackBusLane [2][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][7].cb_test                                      ;
                vDownstreamStackBusLane [2][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][8].cb_test                                      ;
                vDownstreamStackBusLane [2][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][9].cb_test                                      ;
                vDownstreamStackBusLane [2][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][10].cb_test                                      ;
                vDownstreamStackBusLane [2][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][11].cb_test                                      ;
                vDownstreamStackBusLane [2][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][12].cb_test                                      ;
                vDownstreamStackBusLane [2][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][13].cb_test                                      ;
                vDownstreamStackBusLane [2][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][14].cb_test                                      ;
                vDownstreamStackBusLane [2][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][15].cb_test                                      ;
                vDownstreamStackBusLane [2][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][16].cb_test                                      ;
                vDownstreamStackBusLane [2][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][17].cb_test                                      ;
                vDownstreamStackBusLane [2][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][18].cb_test                                      ;
                vDownstreamStackBusLane [2][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][19].cb_test                                      ;
                vDownstreamStackBusLane [2][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][20].cb_test                                      ;
                vDownstreamStackBusLane [2][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][21].cb_test                                      ;
                vDownstreamStackBusLane [2][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][22].cb_test                                      ;
                vDownstreamStackBusLane [2][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][23].cb_test                                      ;
                vDownstreamStackBusLane [2][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][24].cb_test                                      ;
                vDownstreamStackBusLane [2][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][25].cb_test                                      ;
                vDownstreamStackBusLane [2][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][26].cb_test                                      ;
                vDownstreamStackBusLane [2][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][27].cb_test                                      ;
                vDownstreamStackBusLane [2][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][28].cb_test                                      ;
                vDownstreamStackBusLane [2][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][29].cb_test                                      ;
                vDownstreamStackBusLane [2][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][30].cb_test                                      ;
                vDownstreamStackBusLane [2][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[2][31].cb_test                                      ;
                vDownstreamStackBusLane [2][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [2][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[3][0].cb_test                                      ;
                vDownstreamStackBusLane [3][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][1].cb_test                                      ;
                vDownstreamStackBusLane [3][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][2].cb_test                                      ;
                vDownstreamStackBusLane [3][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][3].cb_test                                      ;
                vDownstreamStackBusLane [3][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][4].cb_test                                      ;
                vDownstreamStackBusLane [3][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][5].cb_test                                      ;
                vDownstreamStackBusLane [3][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][6].cb_test                                      ;
                vDownstreamStackBusLane [3][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][7].cb_test                                      ;
                vDownstreamStackBusLane [3][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][8].cb_test                                      ;
                vDownstreamStackBusLane [3][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][9].cb_test                                      ;
                vDownstreamStackBusLane [3][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][10].cb_test                                      ;
                vDownstreamStackBusLane [3][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][11].cb_test                                      ;
                vDownstreamStackBusLane [3][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][12].cb_test                                      ;
                vDownstreamStackBusLane [3][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][13].cb_test                                      ;
                vDownstreamStackBusLane [3][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][14].cb_test                                      ;
                vDownstreamStackBusLane [3][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][15].cb_test                                      ;
                vDownstreamStackBusLane [3][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][16].cb_test                                      ;
                vDownstreamStackBusLane [3][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][17].cb_test                                      ;
                vDownstreamStackBusLane [3][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][18].cb_test                                      ;
                vDownstreamStackBusLane [3][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][19].cb_test                                      ;
                vDownstreamStackBusLane [3][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][20].cb_test                                      ;
                vDownstreamStackBusLane [3][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][21].cb_test                                      ;
                vDownstreamStackBusLane [3][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][22].cb_test                                      ;
                vDownstreamStackBusLane [3][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][23].cb_test                                      ;
                vDownstreamStackBusLane [3][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][24].cb_test                                      ;
                vDownstreamStackBusLane [3][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][25].cb_test                                      ;
                vDownstreamStackBusLane [3][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][26].cb_test                                      ;
                vDownstreamStackBusLane [3][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][27].cb_test                                      ;
                vDownstreamStackBusLane [3][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][28].cb_test                                      ;
                vDownstreamStackBusLane [3][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][29].cb_test                                      ;
                vDownstreamStackBusLane [3][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][30].cb_test                                      ;
                vDownstreamStackBusLane [3][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[3][31].cb_test                                      ;
                vDownstreamStackBusLane [3][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [3][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[4][0].cb_test                                      ;
                vDownstreamStackBusLane [4][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][1].cb_test                                      ;
                vDownstreamStackBusLane [4][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][2].cb_test                                      ;
                vDownstreamStackBusLane [4][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][3].cb_test                                      ;
                vDownstreamStackBusLane [4][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][4].cb_test                                      ;
                vDownstreamStackBusLane [4][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][5].cb_test                                      ;
                vDownstreamStackBusLane [4][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][6].cb_test                                      ;
                vDownstreamStackBusLane [4][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][7].cb_test                                      ;
                vDownstreamStackBusLane [4][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][8].cb_test                                      ;
                vDownstreamStackBusLane [4][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][9].cb_test                                      ;
                vDownstreamStackBusLane [4][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][10].cb_test                                      ;
                vDownstreamStackBusLane [4][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][11].cb_test                                      ;
                vDownstreamStackBusLane [4][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][12].cb_test                                      ;
                vDownstreamStackBusLane [4][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][13].cb_test                                      ;
                vDownstreamStackBusLane [4][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][14].cb_test                                      ;
                vDownstreamStackBusLane [4][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][15].cb_test                                      ;
                vDownstreamStackBusLane [4][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][16].cb_test                                      ;
                vDownstreamStackBusLane [4][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][17].cb_test                                      ;
                vDownstreamStackBusLane [4][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][18].cb_test                                      ;
                vDownstreamStackBusLane [4][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][19].cb_test                                      ;
                vDownstreamStackBusLane [4][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][20].cb_test                                      ;
                vDownstreamStackBusLane [4][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][21].cb_test                                      ;
                vDownstreamStackBusLane [4][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][22].cb_test                                      ;
                vDownstreamStackBusLane [4][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][23].cb_test                                      ;
                vDownstreamStackBusLane [4][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][24].cb_test                                      ;
                vDownstreamStackBusLane [4][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][25].cb_test                                      ;
                vDownstreamStackBusLane [4][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][26].cb_test                                      ;
                vDownstreamStackBusLane [4][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][27].cb_test                                      ;
                vDownstreamStackBusLane [4][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][28].cb_test                                      ;
                vDownstreamStackBusLane [4][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][29].cb_test                                      ;
                vDownstreamStackBusLane [4][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][30].cb_test                                      ;
                vDownstreamStackBusLane [4][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[4][31].cb_test                                      ;
                vDownstreamStackBusLane [4][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [4][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[5][0].cb_test                                      ;
                vDownstreamStackBusLane [5][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][1].cb_test                                      ;
                vDownstreamStackBusLane [5][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][2].cb_test                                      ;
                vDownstreamStackBusLane [5][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][3].cb_test                                      ;
                vDownstreamStackBusLane [5][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][4].cb_test                                      ;
                vDownstreamStackBusLane [5][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][5].cb_test                                      ;
                vDownstreamStackBusLane [5][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][6].cb_test                                      ;
                vDownstreamStackBusLane [5][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][7].cb_test                                      ;
                vDownstreamStackBusLane [5][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][8].cb_test                                      ;
                vDownstreamStackBusLane [5][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][9].cb_test                                      ;
                vDownstreamStackBusLane [5][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][10].cb_test                                      ;
                vDownstreamStackBusLane [5][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][11].cb_test                                      ;
                vDownstreamStackBusLane [5][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][12].cb_test                                      ;
                vDownstreamStackBusLane [5][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][13].cb_test                                      ;
                vDownstreamStackBusLane [5][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][14].cb_test                                      ;
                vDownstreamStackBusLane [5][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][15].cb_test                                      ;
                vDownstreamStackBusLane [5][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][16].cb_test                                      ;
                vDownstreamStackBusLane [5][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][17].cb_test                                      ;
                vDownstreamStackBusLane [5][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][18].cb_test                                      ;
                vDownstreamStackBusLane [5][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][19].cb_test                                      ;
                vDownstreamStackBusLane [5][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][20].cb_test                                      ;
                vDownstreamStackBusLane [5][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][21].cb_test                                      ;
                vDownstreamStackBusLane [5][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][22].cb_test                                      ;
                vDownstreamStackBusLane [5][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][23].cb_test                                      ;
                vDownstreamStackBusLane [5][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][24].cb_test                                      ;
                vDownstreamStackBusLane [5][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][25].cb_test                                      ;
                vDownstreamStackBusLane [5][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][26].cb_test                                      ;
                vDownstreamStackBusLane [5][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][27].cb_test                                      ;
                vDownstreamStackBusLane [5][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][28].cb_test                                      ;
                vDownstreamStackBusLane [5][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][29].cb_test                                      ;
                vDownstreamStackBusLane [5][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][30].cb_test                                      ;
                vDownstreamStackBusLane [5][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[5][31].cb_test                                      ;
                vDownstreamStackBusLane [5][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [5][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[6][0].cb_test                                      ;
                vDownstreamStackBusLane [6][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][1].cb_test                                      ;
                vDownstreamStackBusLane [6][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][2].cb_test                                      ;
                vDownstreamStackBusLane [6][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][3].cb_test                                      ;
                vDownstreamStackBusLane [6][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][4].cb_test                                      ;
                vDownstreamStackBusLane [6][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][5].cb_test                                      ;
                vDownstreamStackBusLane [6][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][6].cb_test                                      ;
                vDownstreamStackBusLane [6][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][7].cb_test                                      ;
                vDownstreamStackBusLane [6][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][8].cb_test                                      ;
                vDownstreamStackBusLane [6][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][9].cb_test                                      ;
                vDownstreamStackBusLane [6][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][10].cb_test                                      ;
                vDownstreamStackBusLane [6][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][11].cb_test                                      ;
                vDownstreamStackBusLane [6][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][12].cb_test                                      ;
                vDownstreamStackBusLane [6][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][13].cb_test                                      ;
                vDownstreamStackBusLane [6][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][14].cb_test                                      ;
                vDownstreamStackBusLane [6][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][15].cb_test                                      ;
                vDownstreamStackBusLane [6][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][16].cb_test                                      ;
                vDownstreamStackBusLane [6][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][17].cb_test                                      ;
                vDownstreamStackBusLane [6][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][18].cb_test                                      ;
                vDownstreamStackBusLane [6][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][19].cb_test                                      ;
                vDownstreamStackBusLane [6][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][20].cb_test                                      ;
                vDownstreamStackBusLane [6][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][21].cb_test                                      ;
                vDownstreamStackBusLane [6][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][22].cb_test                                      ;
                vDownstreamStackBusLane [6][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][23].cb_test                                      ;
                vDownstreamStackBusLane [6][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][24].cb_test                                      ;
                vDownstreamStackBusLane [6][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][25].cb_test                                      ;
                vDownstreamStackBusLane [6][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][26].cb_test                                      ;
                vDownstreamStackBusLane [6][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][27].cb_test                                      ;
                vDownstreamStackBusLane [6][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][28].cb_test                                      ;
                vDownstreamStackBusLane [6][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][29].cb_test                                      ;
                vDownstreamStackBusLane [6][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][30].cb_test                                      ;
                vDownstreamStackBusLane [6][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[6][31].cb_test                                      ;
                vDownstreamStackBusLane [6][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [6][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[7][0].cb_test                                      ;
                vDownstreamStackBusLane [7][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][1].cb_test                                      ;
                vDownstreamStackBusLane [7][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][2].cb_test                                      ;
                vDownstreamStackBusLane [7][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][3].cb_test                                      ;
                vDownstreamStackBusLane [7][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][4].cb_test                                      ;
                vDownstreamStackBusLane [7][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][5].cb_test                                      ;
                vDownstreamStackBusLane [7][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][6].cb_test                                      ;
                vDownstreamStackBusLane [7][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][7].cb_test                                      ;
                vDownstreamStackBusLane [7][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][8].cb_test                                      ;
                vDownstreamStackBusLane [7][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][9].cb_test                                      ;
                vDownstreamStackBusLane [7][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][10].cb_test                                      ;
                vDownstreamStackBusLane [7][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][11].cb_test                                      ;
                vDownstreamStackBusLane [7][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][12].cb_test                                      ;
                vDownstreamStackBusLane [7][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][13].cb_test                                      ;
                vDownstreamStackBusLane [7][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][14].cb_test                                      ;
                vDownstreamStackBusLane [7][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][15].cb_test                                      ;
                vDownstreamStackBusLane [7][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][16].cb_test                                      ;
                vDownstreamStackBusLane [7][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][17].cb_test                                      ;
                vDownstreamStackBusLane [7][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][18].cb_test                                      ;
                vDownstreamStackBusLane [7][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][19].cb_test                                      ;
                vDownstreamStackBusLane [7][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][20].cb_test                                      ;
                vDownstreamStackBusLane [7][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][21].cb_test                                      ;
                vDownstreamStackBusLane [7][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][22].cb_test                                      ;
                vDownstreamStackBusLane [7][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][23].cb_test                                      ;
                vDownstreamStackBusLane [7][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][24].cb_test                                      ;
                vDownstreamStackBusLane [7][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][25].cb_test                                      ;
                vDownstreamStackBusLane [7][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][26].cb_test                                      ;
                vDownstreamStackBusLane [7][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][27].cb_test                                      ;
                vDownstreamStackBusLane [7][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][28].cb_test                                      ;
                vDownstreamStackBusLane [7][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][29].cb_test                                      ;
                vDownstreamStackBusLane [7][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][30].cb_test                                      ;
                vDownstreamStackBusLane [7][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[7][31].cb_test                                      ;
                vDownstreamStackBusLane [7][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [7][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[8][0].cb_test                                      ;
                vDownstreamStackBusLane [8][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][1].cb_test                                      ;
                vDownstreamStackBusLane [8][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][2].cb_test                                      ;
                vDownstreamStackBusLane [8][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][3].cb_test                                      ;
                vDownstreamStackBusLane [8][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][4].cb_test                                      ;
                vDownstreamStackBusLane [8][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][5].cb_test                                      ;
                vDownstreamStackBusLane [8][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][6].cb_test                                      ;
                vDownstreamStackBusLane [8][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][7].cb_test                                      ;
                vDownstreamStackBusLane [8][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][8].cb_test                                      ;
                vDownstreamStackBusLane [8][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][9].cb_test                                      ;
                vDownstreamStackBusLane [8][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][10].cb_test                                      ;
                vDownstreamStackBusLane [8][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][11].cb_test                                      ;
                vDownstreamStackBusLane [8][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][12].cb_test                                      ;
                vDownstreamStackBusLane [8][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][13].cb_test                                      ;
                vDownstreamStackBusLane [8][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][14].cb_test                                      ;
                vDownstreamStackBusLane [8][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][15].cb_test                                      ;
                vDownstreamStackBusLane [8][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][16].cb_test                                      ;
                vDownstreamStackBusLane [8][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][17].cb_test                                      ;
                vDownstreamStackBusLane [8][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][18].cb_test                                      ;
                vDownstreamStackBusLane [8][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][19].cb_test                                      ;
                vDownstreamStackBusLane [8][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][20].cb_test                                      ;
                vDownstreamStackBusLane [8][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][21].cb_test                                      ;
                vDownstreamStackBusLane [8][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][22].cb_test                                      ;
                vDownstreamStackBusLane [8][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][23].cb_test                                      ;
                vDownstreamStackBusLane [8][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][24].cb_test                                      ;
                vDownstreamStackBusLane [8][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][25].cb_test                                      ;
                vDownstreamStackBusLane [8][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][26].cb_test                                      ;
                vDownstreamStackBusLane [8][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][27].cb_test                                      ;
                vDownstreamStackBusLane [8][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][28].cb_test                                      ;
                vDownstreamStackBusLane [8][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][29].cb_test                                      ;
                vDownstreamStackBusLane [8][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][30].cb_test                                      ;
                vDownstreamStackBusLane [8][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[8][31].cb_test                                      ;
                vDownstreamStackBusLane [8][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [8][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[9][0].cb_test                                      ;
                vDownstreamStackBusLane [9][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][1].cb_test                                      ;
                vDownstreamStackBusLane [9][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][2].cb_test                                      ;
                vDownstreamStackBusLane [9][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][3].cb_test                                      ;
                vDownstreamStackBusLane [9][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][4].cb_test                                      ;
                vDownstreamStackBusLane [9][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][5].cb_test                                      ;
                vDownstreamStackBusLane [9][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][6].cb_test                                      ;
                vDownstreamStackBusLane [9][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][7].cb_test                                      ;
                vDownstreamStackBusLane [9][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][8].cb_test                                      ;
                vDownstreamStackBusLane [9][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][9].cb_test                                      ;
                vDownstreamStackBusLane [9][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][10].cb_test                                      ;
                vDownstreamStackBusLane [9][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][11].cb_test                                      ;
                vDownstreamStackBusLane [9][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][12].cb_test                                      ;
                vDownstreamStackBusLane [9][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][13].cb_test                                      ;
                vDownstreamStackBusLane [9][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][14].cb_test                                      ;
                vDownstreamStackBusLane [9][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][15].cb_test                                      ;
                vDownstreamStackBusLane [9][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][16].cb_test                                      ;
                vDownstreamStackBusLane [9][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][17].cb_test                                      ;
                vDownstreamStackBusLane [9][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][18].cb_test                                      ;
                vDownstreamStackBusLane [9][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][19].cb_test                                      ;
                vDownstreamStackBusLane [9][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][20].cb_test                                      ;
                vDownstreamStackBusLane [9][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][21].cb_test                                      ;
                vDownstreamStackBusLane [9][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][22].cb_test                                      ;
                vDownstreamStackBusLane [9][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][23].cb_test                                      ;
                vDownstreamStackBusLane [9][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][24].cb_test                                      ;
                vDownstreamStackBusLane [9][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][25].cb_test                                      ;
                vDownstreamStackBusLane [9][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][26].cb_test                                      ;
                vDownstreamStackBusLane [9][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][27].cb_test                                      ;
                vDownstreamStackBusLane [9][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][28].cb_test                                      ;
                vDownstreamStackBusLane [9][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][29].cb_test                                      ;
                vDownstreamStackBusLane [9][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][30].cb_test                                      ;
                vDownstreamStackBusLane [9][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[9][31].cb_test                                      ;
                vDownstreamStackBusLane [9][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [9][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[10][0].cb_test                                      ;
                vDownstreamStackBusLane [10][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][1].cb_test                                      ;
                vDownstreamStackBusLane [10][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][2].cb_test                                      ;
                vDownstreamStackBusLane [10][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][3].cb_test                                      ;
                vDownstreamStackBusLane [10][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][4].cb_test                                      ;
                vDownstreamStackBusLane [10][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][5].cb_test                                      ;
                vDownstreamStackBusLane [10][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][6].cb_test                                      ;
                vDownstreamStackBusLane [10][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][7].cb_test                                      ;
                vDownstreamStackBusLane [10][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][8].cb_test                                      ;
                vDownstreamStackBusLane [10][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][9].cb_test                                      ;
                vDownstreamStackBusLane [10][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][10].cb_test                                      ;
                vDownstreamStackBusLane [10][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][11].cb_test                                      ;
                vDownstreamStackBusLane [10][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][12].cb_test                                      ;
                vDownstreamStackBusLane [10][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][13].cb_test                                      ;
                vDownstreamStackBusLane [10][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][14].cb_test                                      ;
                vDownstreamStackBusLane [10][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][15].cb_test                                      ;
                vDownstreamStackBusLane [10][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][16].cb_test                                      ;
                vDownstreamStackBusLane [10][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][17].cb_test                                      ;
                vDownstreamStackBusLane [10][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][18].cb_test                                      ;
                vDownstreamStackBusLane [10][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][19].cb_test                                      ;
                vDownstreamStackBusLane [10][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][20].cb_test                                      ;
                vDownstreamStackBusLane [10][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][21].cb_test                                      ;
                vDownstreamStackBusLane [10][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][22].cb_test                                      ;
                vDownstreamStackBusLane [10][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][23].cb_test                                      ;
                vDownstreamStackBusLane [10][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][24].cb_test                                      ;
                vDownstreamStackBusLane [10][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][25].cb_test                                      ;
                vDownstreamStackBusLane [10][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][26].cb_test                                      ;
                vDownstreamStackBusLane [10][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][27].cb_test                                      ;
                vDownstreamStackBusLane [10][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][28].cb_test                                      ;
                vDownstreamStackBusLane [10][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][29].cb_test                                      ;
                vDownstreamStackBusLane [10][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][30].cb_test                                      ;
                vDownstreamStackBusLane [10][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[10][31].cb_test                                      ;
                vDownstreamStackBusLane [10][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [10][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[11][0].cb_test                                      ;
                vDownstreamStackBusLane [11][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][1].cb_test                                      ;
                vDownstreamStackBusLane [11][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][2].cb_test                                      ;
                vDownstreamStackBusLane [11][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][3].cb_test                                      ;
                vDownstreamStackBusLane [11][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][4].cb_test                                      ;
                vDownstreamStackBusLane [11][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][5].cb_test                                      ;
                vDownstreamStackBusLane [11][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][6].cb_test                                      ;
                vDownstreamStackBusLane [11][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][7].cb_test                                      ;
                vDownstreamStackBusLane [11][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][8].cb_test                                      ;
                vDownstreamStackBusLane [11][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][9].cb_test                                      ;
                vDownstreamStackBusLane [11][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][10].cb_test                                      ;
                vDownstreamStackBusLane [11][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][11].cb_test                                      ;
                vDownstreamStackBusLane [11][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][12].cb_test                                      ;
                vDownstreamStackBusLane [11][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][13].cb_test                                      ;
                vDownstreamStackBusLane [11][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][14].cb_test                                      ;
                vDownstreamStackBusLane [11][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][15].cb_test                                      ;
                vDownstreamStackBusLane [11][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][16].cb_test                                      ;
                vDownstreamStackBusLane [11][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][17].cb_test                                      ;
                vDownstreamStackBusLane [11][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][18].cb_test                                      ;
                vDownstreamStackBusLane [11][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][19].cb_test                                      ;
                vDownstreamStackBusLane [11][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][20].cb_test                                      ;
                vDownstreamStackBusLane [11][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][21].cb_test                                      ;
                vDownstreamStackBusLane [11][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][22].cb_test                                      ;
                vDownstreamStackBusLane [11][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][23].cb_test                                      ;
                vDownstreamStackBusLane [11][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][24].cb_test                                      ;
                vDownstreamStackBusLane [11][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][25].cb_test                                      ;
                vDownstreamStackBusLane [11][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][26].cb_test                                      ;
                vDownstreamStackBusLane [11][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][27].cb_test                                      ;
                vDownstreamStackBusLane [11][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][28].cb_test                                      ;
                vDownstreamStackBusLane [11][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][29].cb_test                                      ;
                vDownstreamStackBusLane [11][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][30].cb_test                                      ;
                vDownstreamStackBusLane [11][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[11][31].cb_test                                      ;
                vDownstreamStackBusLane [11][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [11][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[12][0].cb_test                                      ;
                vDownstreamStackBusLane [12][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][1].cb_test                                      ;
                vDownstreamStackBusLane [12][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][2].cb_test                                      ;
                vDownstreamStackBusLane [12][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][3].cb_test                                      ;
                vDownstreamStackBusLane [12][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][4].cb_test                                      ;
                vDownstreamStackBusLane [12][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][5].cb_test                                      ;
                vDownstreamStackBusLane [12][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][6].cb_test                                      ;
                vDownstreamStackBusLane [12][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][7].cb_test                                      ;
                vDownstreamStackBusLane [12][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][8].cb_test                                      ;
                vDownstreamStackBusLane [12][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][9].cb_test                                      ;
                vDownstreamStackBusLane [12][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][10].cb_test                                      ;
                vDownstreamStackBusLane [12][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][11].cb_test                                      ;
                vDownstreamStackBusLane [12][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][12].cb_test                                      ;
                vDownstreamStackBusLane [12][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][13].cb_test                                      ;
                vDownstreamStackBusLane [12][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][14].cb_test                                      ;
                vDownstreamStackBusLane [12][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][15].cb_test                                      ;
                vDownstreamStackBusLane [12][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][16].cb_test                                      ;
                vDownstreamStackBusLane [12][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][17].cb_test                                      ;
                vDownstreamStackBusLane [12][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][18].cb_test                                      ;
                vDownstreamStackBusLane [12][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][19].cb_test                                      ;
                vDownstreamStackBusLane [12][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][20].cb_test                                      ;
                vDownstreamStackBusLane [12][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][21].cb_test                                      ;
                vDownstreamStackBusLane [12][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][22].cb_test                                      ;
                vDownstreamStackBusLane [12][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][23].cb_test                                      ;
                vDownstreamStackBusLane [12][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][24].cb_test                                      ;
                vDownstreamStackBusLane [12][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][25].cb_test                                      ;
                vDownstreamStackBusLane [12][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][26].cb_test                                      ;
                vDownstreamStackBusLane [12][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][27].cb_test                                      ;
                vDownstreamStackBusLane [12][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][28].cb_test                                      ;
                vDownstreamStackBusLane [12][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][29].cb_test                                      ;
                vDownstreamStackBusLane [12][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][30].cb_test                                      ;
                vDownstreamStackBusLane [12][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[12][31].cb_test                                      ;
                vDownstreamStackBusLane [12][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [12][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[13][0].cb_test                                      ;
                vDownstreamStackBusLane [13][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][1].cb_test                                      ;
                vDownstreamStackBusLane [13][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][2].cb_test                                      ;
                vDownstreamStackBusLane [13][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][3].cb_test                                      ;
                vDownstreamStackBusLane [13][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][4].cb_test                                      ;
                vDownstreamStackBusLane [13][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][5].cb_test                                      ;
                vDownstreamStackBusLane [13][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][6].cb_test                                      ;
                vDownstreamStackBusLane [13][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][7].cb_test                                      ;
                vDownstreamStackBusLane [13][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][8].cb_test                                      ;
                vDownstreamStackBusLane [13][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][9].cb_test                                      ;
                vDownstreamStackBusLane [13][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][10].cb_test                                      ;
                vDownstreamStackBusLane [13][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][11].cb_test                                      ;
                vDownstreamStackBusLane [13][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][12].cb_test                                      ;
                vDownstreamStackBusLane [13][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][13].cb_test                                      ;
                vDownstreamStackBusLane [13][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][14].cb_test                                      ;
                vDownstreamStackBusLane [13][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][15].cb_test                                      ;
                vDownstreamStackBusLane [13][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][16].cb_test                                      ;
                vDownstreamStackBusLane [13][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][17].cb_test                                      ;
                vDownstreamStackBusLane [13][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][18].cb_test                                      ;
                vDownstreamStackBusLane [13][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][19].cb_test                                      ;
                vDownstreamStackBusLane [13][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][20].cb_test                                      ;
                vDownstreamStackBusLane [13][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][21].cb_test                                      ;
                vDownstreamStackBusLane [13][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][22].cb_test                                      ;
                vDownstreamStackBusLane [13][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][23].cb_test                                      ;
                vDownstreamStackBusLane [13][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][24].cb_test                                      ;
                vDownstreamStackBusLane [13][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][25].cb_test                                      ;
                vDownstreamStackBusLane [13][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][26].cb_test                                      ;
                vDownstreamStackBusLane [13][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][27].cb_test                                      ;
                vDownstreamStackBusLane [13][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][28].cb_test                                      ;
                vDownstreamStackBusLane [13][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][29].cb_test                                      ;
                vDownstreamStackBusLane [13][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][30].cb_test                                      ;
                vDownstreamStackBusLane [13][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[13][31].cb_test                                      ;
                vDownstreamStackBusLane [13][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [13][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[14][0].cb_test                                      ;
                vDownstreamStackBusLane [14][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][1].cb_test                                      ;
                vDownstreamStackBusLane [14][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][2].cb_test                                      ;
                vDownstreamStackBusLane [14][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][3].cb_test                                      ;
                vDownstreamStackBusLane [14][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][4].cb_test                                      ;
                vDownstreamStackBusLane [14][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][5].cb_test                                      ;
                vDownstreamStackBusLane [14][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][6].cb_test                                      ;
                vDownstreamStackBusLane [14][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][7].cb_test                                      ;
                vDownstreamStackBusLane [14][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][8].cb_test                                      ;
                vDownstreamStackBusLane [14][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][9].cb_test                                      ;
                vDownstreamStackBusLane [14][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][10].cb_test                                      ;
                vDownstreamStackBusLane [14][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][11].cb_test                                      ;
                vDownstreamStackBusLane [14][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][12].cb_test                                      ;
                vDownstreamStackBusLane [14][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][13].cb_test                                      ;
                vDownstreamStackBusLane [14][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][14].cb_test                                      ;
                vDownstreamStackBusLane [14][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][15].cb_test                                      ;
                vDownstreamStackBusLane [14][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][16].cb_test                                      ;
                vDownstreamStackBusLane [14][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][17].cb_test                                      ;
                vDownstreamStackBusLane [14][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][18].cb_test                                      ;
                vDownstreamStackBusLane [14][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][19].cb_test                                      ;
                vDownstreamStackBusLane [14][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][20].cb_test                                      ;
                vDownstreamStackBusLane [14][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][21].cb_test                                      ;
                vDownstreamStackBusLane [14][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][22].cb_test                                      ;
                vDownstreamStackBusLane [14][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][23].cb_test                                      ;
                vDownstreamStackBusLane [14][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][24].cb_test                                      ;
                vDownstreamStackBusLane [14][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][25].cb_test                                      ;
                vDownstreamStackBusLane [14][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][26].cb_test                                      ;
                vDownstreamStackBusLane [14][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][27].cb_test                                      ;
                vDownstreamStackBusLane [14][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][28].cb_test                                      ;
                vDownstreamStackBusLane [14][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][29].cb_test                                      ;
                vDownstreamStackBusLane [14][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][30].cb_test                                      ;
                vDownstreamStackBusLane [14][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[14][31].cb_test                                      ;
                vDownstreamStackBusLane [14][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [14][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[15][0].cb_test                                      ;
                vDownstreamStackBusLane [15][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][1].cb_test                                      ;
                vDownstreamStackBusLane [15][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][2].cb_test                                      ;
                vDownstreamStackBusLane [15][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][3].cb_test                                      ;
                vDownstreamStackBusLane [15][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][4].cb_test                                      ;
                vDownstreamStackBusLane [15][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][5].cb_test                                      ;
                vDownstreamStackBusLane [15][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][6].cb_test                                      ;
                vDownstreamStackBusLane [15][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][7].cb_test                                      ;
                vDownstreamStackBusLane [15][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][8].cb_test                                      ;
                vDownstreamStackBusLane [15][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][9].cb_test                                      ;
                vDownstreamStackBusLane [15][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][10].cb_test                                      ;
                vDownstreamStackBusLane [15][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][11].cb_test                                      ;
                vDownstreamStackBusLane [15][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][12].cb_test                                      ;
                vDownstreamStackBusLane [15][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][13].cb_test                                      ;
                vDownstreamStackBusLane [15][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][14].cb_test                                      ;
                vDownstreamStackBusLane [15][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][15].cb_test                                      ;
                vDownstreamStackBusLane [15][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][16].cb_test                                      ;
                vDownstreamStackBusLane [15][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][17].cb_test                                      ;
                vDownstreamStackBusLane [15][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][18].cb_test                                      ;
                vDownstreamStackBusLane [15][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][19].cb_test                                      ;
                vDownstreamStackBusLane [15][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][20].cb_test                                      ;
                vDownstreamStackBusLane [15][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][21].cb_test                                      ;
                vDownstreamStackBusLane [15][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][22].cb_test                                      ;
                vDownstreamStackBusLane [15][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][23].cb_test                                      ;
                vDownstreamStackBusLane [15][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][24].cb_test                                      ;
                vDownstreamStackBusLane [15][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][25].cb_test                                      ;
                vDownstreamStackBusLane [15][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][26].cb_test                                      ;
                vDownstreamStackBusLane [15][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][27].cb_test                                      ;
                vDownstreamStackBusLane [15][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][28].cb_test                                      ;
                vDownstreamStackBusLane [15][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][29].cb_test                                      ;
                vDownstreamStackBusLane [15][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][30].cb_test                                      ;
                vDownstreamStackBusLane [15][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[15][31].cb_test                                      ;
                vDownstreamStackBusLane [15][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [15][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[16][0].cb_test                                      ;
                vDownstreamStackBusLane [16][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][1].cb_test                                      ;
                vDownstreamStackBusLane [16][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][2].cb_test                                      ;
                vDownstreamStackBusLane [16][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][3].cb_test                                      ;
                vDownstreamStackBusLane [16][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][4].cb_test                                      ;
                vDownstreamStackBusLane [16][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][5].cb_test                                      ;
                vDownstreamStackBusLane [16][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][6].cb_test                                      ;
                vDownstreamStackBusLane [16][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][7].cb_test                                      ;
                vDownstreamStackBusLane [16][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][8].cb_test                                      ;
                vDownstreamStackBusLane [16][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][9].cb_test                                      ;
                vDownstreamStackBusLane [16][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][10].cb_test                                      ;
                vDownstreamStackBusLane [16][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][11].cb_test                                      ;
                vDownstreamStackBusLane [16][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][12].cb_test                                      ;
                vDownstreamStackBusLane [16][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][13].cb_test                                      ;
                vDownstreamStackBusLane [16][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][14].cb_test                                      ;
                vDownstreamStackBusLane [16][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][15].cb_test                                      ;
                vDownstreamStackBusLane [16][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][16].cb_test                                      ;
                vDownstreamStackBusLane [16][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][17].cb_test                                      ;
                vDownstreamStackBusLane [16][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][18].cb_test                                      ;
                vDownstreamStackBusLane [16][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][19].cb_test                                      ;
                vDownstreamStackBusLane [16][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][20].cb_test                                      ;
                vDownstreamStackBusLane [16][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][21].cb_test                                      ;
                vDownstreamStackBusLane [16][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][22].cb_test                                      ;
                vDownstreamStackBusLane [16][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][23].cb_test                                      ;
                vDownstreamStackBusLane [16][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][24].cb_test                                      ;
                vDownstreamStackBusLane [16][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][25].cb_test                                      ;
                vDownstreamStackBusLane [16][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][26].cb_test                                      ;
                vDownstreamStackBusLane [16][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][27].cb_test                                      ;
                vDownstreamStackBusLane [16][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][28].cb_test                                      ;
                vDownstreamStackBusLane [16][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][29].cb_test                                      ;
                vDownstreamStackBusLane [16][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][30].cb_test                                      ;
                vDownstreamStackBusLane [16][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[16][31].cb_test                                      ;
                vDownstreamStackBusLane [16][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [16][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[17][0].cb_test                                      ;
                vDownstreamStackBusLane [17][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][1].cb_test                                      ;
                vDownstreamStackBusLane [17][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][2].cb_test                                      ;
                vDownstreamStackBusLane [17][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][3].cb_test                                      ;
                vDownstreamStackBusLane [17][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][4].cb_test                                      ;
                vDownstreamStackBusLane [17][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][5].cb_test                                      ;
                vDownstreamStackBusLane [17][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][6].cb_test                                      ;
                vDownstreamStackBusLane [17][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][7].cb_test                                      ;
                vDownstreamStackBusLane [17][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][8].cb_test                                      ;
                vDownstreamStackBusLane [17][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][9].cb_test                                      ;
                vDownstreamStackBusLane [17][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][10].cb_test                                      ;
                vDownstreamStackBusLane [17][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][11].cb_test                                      ;
                vDownstreamStackBusLane [17][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][12].cb_test                                      ;
                vDownstreamStackBusLane [17][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][13].cb_test                                      ;
                vDownstreamStackBusLane [17][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][14].cb_test                                      ;
                vDownstreamStackBusLane [17][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][15].cb_test                                      ;
                vDownstreamStackBusLane [17][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][16].cb_test                                      ;
                vDownstreamStackBusLane [17][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][17].cb_test                                      ;
                vDownstreamStackBusLane [17][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][18].cb_test                                      ;
                vDownstreamStackBusLane [17][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][19].cb_test                                      ;
                vDownstreamStackBusLane [17][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][20].cb_test                                      ;
                vDownstreamStackBusLane [17][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][21].cb_test                                      ;
                vDownstreamStackBusLane [17][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][22].cb_test                                      ;
                vDownstreamStackBusLane [17][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][23].cb_test                                      ;
                vDownstreamStackBusLane [17][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][24].cb_test                                      ;
                vDownstreamStackBusLane [17][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][25].cb_test                                      ;
                vDownstreamStackBusLane [17][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][26].cb_test                                      ;
                vDownstreamStackBusLane [17][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][27].cb_test                                      ;
                vDownstreamStackBusLane [17][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][28].cb_test                                      ;
                vDownstreamStackBusLane [17][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][29].cb_test                                      ;
                vDownstreamStackBusLane [17][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][30].cb_test                                      ;
                vDownstreamStackBusLane [17][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[17][31].cb_test                                      ;
                vDownstreamStackBusLane [17][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [17][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[18][0].cb_test                                      ;
                vDownstreamStackBusLane [18][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][1].cb_test                                      ;
                vDownstreamStackBusLane [18][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][2].cb_test                                      ;
                vDownstreamStackBusLane [18][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][3].cb_test                                      ;
                vDownstreamStackBusLane [18][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][4].cb_test                                      ;
                vDownstreamStackBusLane [18][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][5].cb_test                                      ;
                vDownstreamStackBusLane [18][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][6].cb_test                                      ;
                vDownstreamStackBusLane [18][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][7].cb_test                                      ;
                vDownstreamStackBusLane [18][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][8].cb_test                                      ;
                vDownstreamStackBusLane [18][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][9].cb_test                                      ;
                vDownstreamStackBusLane [18][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][10].cb_test                                      ;
                vDownstreamStackBusLane [18][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][11].cb_test                                      ;
                vDownstreamStackBusLane [18][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][12].cb_test                                      ;
                vDownstreamStackBusLane [18][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][13].cb_test                                      ;
                vDownstreamStackBusLane [18][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][14].cb_test                                      ;
                vDownstreamStackBusLane [18][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][15].cb_test                                      ;
                vDownstreamStackBusLane [18][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][16].cb_test                                      ;
                vDownstreamStackBusLane [18][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][17].cb_test                                      ;
                vDownstreamStackBusLane [18][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][18].cb_test                                      ;
                vDownstreamStackBusLane [18][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][19].cb_test                                      ;
                vDownstreamStackBusLane [18][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][20].cb_test                                      ;
                vDownstreamStackBusLane [18][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][21].cb_test                                      ;
                vDownstreamStackBusLane [18][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][22].cb_test                                      ;
                vDownstreamStackBusLane [18][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][23].cb_test                                      ;
                vDownstreamStackBusLane [18][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][24].cb_test                                      ;
                vDownstreamStackBusLane [18][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][25].cb_test                                      ;
                vDownstreamStackBusLane [18][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][26].cb_test                                      ;
                vDownstreamStackBusLane [18][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][27].cb_test                                      ;
                vDownstreamStackBusLane [18][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][28].cb_test                                      ;
                vDownstreamStackBusLane [18][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][29].cb_test                                      ;
                vDownstreamStackBusLane [18][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][30].cb_test                                      ;
                vDownstreamStackBusLane [18][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[18][31].cb_test                                      ;
                vDownstreamStackBusLane [18][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [18][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[19][0].cb_test                                      ;
                vDownstreamStackBusLane [19][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][1].cb_test                                      ;
                vDownstreamStackBusLane [19][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][2].cb_test                                      ;
                vDownstreamStackBusLane [19][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][3].cb_test                                      ;
                vDownstreamStackBusLane [19][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][4].cb_test                                      ;
                vDownstreamStackBusLane [19][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][5].cb_test                                      ;
                vDownstreamStackBusLane [19][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][6].cb_test                                      ;
                vDownstreamStackBusLane [19][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][7].cb_test                                      ;
                vDownstreamStackBusLane [19][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][8].cb_test                                      ;
                vDownstreamStackBusLane [19][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][9].cb_test                                      ;
                vDownstreamStackBusLane [19][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][10].cb_test                                      ;
                vDownstreamStackBusLane [19][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][11].cb_test                                      ;
                vDownstreamStackBusLane [19][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][12].cb_test                                      ;
                vDownstreamStackBusLane [19][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][13].cb_test                                      ;
                vDownstreamStackBusLane [19][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][14].cb_test                                      ;
                vDownstreamStackBusLane [19][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][15].cb_test                                      ;
                vDownstreamStackBusLane [19][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][16].cb_test                                      ;
                vDownstreamStackBusLane [19][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][17].cb_test                                      ;
                vDownstreamStackBusLane [19][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][18].cb_test                                      ;
                vDownstreamStackBusLane [19][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][19].cb_test                                      ;
                vDownstreamStackBusLane [19][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][20].cb_test                                      ;
                vDownstreamStackBusLane [19][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][21].cb_test                                      ;
                vDownstreamStackBusLane [19][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][22].cb_test                                      ;
                vDownstreamStackBusLane [19][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][23].cb_test                                      ;
                vDownstreamStackBusLane [19][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][24].cb_test                                      ;
                vDownstreamStackBusLane [19][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][25].cb_test                                      ;
                vDownstreamStackBusLane [19][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][26].cb_test                                      ;
                vDownstreamStackBusLane [19][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][27].cb_test                                      ;
                vDownstreamStackBusLane [19][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][28].cb_test                                      ;
                vDownstreamStackBusLane [19][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][29].cb_test                                      ;
                vDownstreamStackBusLane [19][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][30].cb_test                                      ;
                vDownstreamStackBusLane [19][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[19][31].cb_test                                      ;
                vDownstreamStackBusLane [19][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [19][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[20][0].cb_test                                      ;
                vDownstreamStackBusLane [20][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][1].cb_test                                      ;
                vDownstreamStackBusLane [20][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][2].cb_test                                      ;
                vDownstreamStackBusLane [20][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][3].cb_test                                      ;
                vDownstreamStackBusLane [20][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][4].cb_test                                      ;
                vDownstreamStackBusLane [20][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][5].cb_test                                      ;
                vDownstreamStackBusLane [20][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][6].cb_test                                      ;
                vDownstreamStackBusLane [20][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][7].cb_test                                      ;
                vDownstreamStackBusLane [20][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][8].cb_test                                      ;
                vDownstreamStackBusLane [20][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][9].cb_test                                      ;
                vDownstreamStackBusLane [20][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][10].cb_test                                      ;
                vDownstreamStackBusLane [20][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][11].cb_test                                      ;
                vDownstreamStackBusLane [20][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][12].cb_test                                      ;
                vDownstreamStackBusLane [20][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][13].cb_test                                      ;
                vDownstreamStackBusLane [20][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][14].cb_test                                      ;
                vDownstreamStackBusLane [20][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][15].cb_test                                      ;
                vDownstreamStackBusLane [20][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][16].cb_test                                      ;
                vDownstreamStackBusLane [20][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][17].cb_test                                      ;
                vDownstreamStackBusLane [20][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][18].cb_test                                      ;
                vDownstreamStackBusLane [20][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][19].cb_test                                      ;
                vDownstreamStackBusLane [20][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][20].cb_test                                      ;
                vDownstreamStackBusLane [20][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][21].cb_test                                      ;
                vDownstreamStackBusLane [20][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][22].cb_test                                      ;
                vDownstreamStackBusLane [20][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][23].cb_test                                      ;
                vDownstreamStackBusLane [20][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][24].cb_test                                      ;
                vDownstreamStackBusLane [20][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][25].cb_test                                      ;
                vDownstreamStackBusLane [20][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][26].cb_test                                      ;
                vDownstreamStackBusLane [20][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][27].cb_test                                      ;
                vDownstreamStackBusLane [20][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][28].cb_test                                      ;
                vDownstreamStackBusLane [20][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][29].cb_test                                      ;
                vDownstreamStackBusLane [20][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][30].cb_test                                      ;
                vDownstreamStackBusLane [20][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[20][31].cb_test                                      ;
                vDownstreamStackBusLane [20][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [20][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[21][0].cb_test                                      ;
                vDownstreamStackBusLane [21][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][1].cb_test                                      ;
                vDownstreamStackBusLane [21][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][2].cb_test                                      ;
                vDownstreamStackBusLane [21][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][3].cb_test                                      ;
                vDownstreamStackBusLane [21][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][4].cb_test                                      ;
                vDownstreamStackBusLane [21][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][5].cb_test                                      ;
                vDownstreamStackBusLane [21][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][6].cb_test                                      ;
                vDownstreamStackBusLane [21][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][7].cb_test                                      ;
                vDownstreamStackBusLane [21][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][8].cb_test                                      ;
                vDownstreamStackBusLane [21][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][9].cb_test                                      ;
                vDownstreamStackBusLane [21][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][10].cb_test                                      ;
                vDownstreamStackBusLane [21][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][11].cb_test                                      ;
                vDownstreamStackBusLane [21][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][12].cb_test                                      ;
                vDownstreamStackBusLane [21][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][13].cb_test                                      ;
                vDownstreamStackBusLane [21][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][14].cb_test                                      ;
                vDownstreamStackBusLane [21][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][15].cb_test                                      ;
                vDownstreamStackBusLane [21][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][16].cb_test                                      ;
                vDownstreamStackBusLane [21][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][17].cb_test                                      ;
                vDownstreamStackBusLane [21][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][18].cb_test                                      ;
                vDownstreamStackBusLane [21][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][19].cb_test                                      ;
                vDownstreamStackBusLane [21][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][20].cb_test                                      ;
                vDownstreamStackBusLane [21][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][21].cb_test                                      ;
                vDownstreamStackBusLane [21][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][22].cb_test                                      ;
                vDownstreamStackBusLane [21][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][23].cb_test                                      ;
                vDownstreamStackBusLane [21][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][24].cb_test                                      ;
                vDownstreamStackBusLane [21][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][25].cb_test                                      ;
                vDownstreamStackBusLane [21][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][26].cb_test                                      ;
                vDownstreamStackBusLane [21][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][27].cb_test                                      ;
                vDownstreamStackBusLane [21][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][28].cb_test                                      ;
                vDownstreamStackBusLane [21][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][29].cb_test                                      ;
                vDownstreamStackBusLane [21][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][30].cb_test                                      ;
                vDownstreamStackBusLane [21][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[21][31].cb_test                                      ;
                vDownstreamStackBusLane [21][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [21][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[22][0].cb_test                                      ;
                vDownstreamStackBusLane [22][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][1].cb_test                                      ;
                vDownstreamStackBusLane [22][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][2].cb_test                                      ;
                vDownstreamStackBusLane [22][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][3].cb_test                                      ;
                vDownstreamStackBusLane [22][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][4].cb_test                                      ;
                vDownstreamStackBusLane [22][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][5].cb_test                                      ;
                vDownstreamStackBusLane [22][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][6].cb_test                                      ;
                vDownstreamStackBusLane [22][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][7].cb_test                                      ;
                vDownstreamStackBusLane [22][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][8].cb_test                                      ;
                vDownstreamStackBusLane [22][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][9].cb_test                                      ;
                vDownstreamStackBusLane [22][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][10].cb_test                                      ;
                vDownstreamStackBusLane [22][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][11].cb_test                                      ;
                vDownstreamStackBusLane [22][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][12].cb_test                                      ;
                vDownstreamStackBusLane [22][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][13].cb_test                                      ;
                vDownstreamStackBusLane [22][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][14].cb_test                                      ;
                vDownstreamStackBusLane [22][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][15].cb_test                                      ;
                vDownstreamStackBusLane [22][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][16].cb_test                                      ;
                vDownstreamStackBusLane [22][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][17].cb_test                                      ;
                vDownstreamStackBusLane [22][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][18].cb_test                                      ;
                vDownstreamStackBusLane [22][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][19].cb_test                                      ;
                vDownstreamStackBusLane [22][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][20].cb_test                                      ;
                vDownstreamStackBusLane [22][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][21].cb_test                                      ;
                vDownstreamStackBusLane [22][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][22].cb_test                                      ;
                vDownstreamStackBusLane [22][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][23].cb_test                                      ;
                vDownstreamStackBusLane [22][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][24].cb_test                                      ;
                vDownstreamStackBusLane [22][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][25].cb_test                                      ;
                vDownstreamStackBusLane [22][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][26].cb_test                                      ;
                vDownstreamStackBusLane [22][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][27].cb_test                                      ;
                vDownstreamStackBusLane [22][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][28].cb_test                                      ;
                vDownstreamStackBusLane [22][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][29].cb_test                                      ;
                vDownstreamStackBusLane [22][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][30].cb_test                                      ;
                vDownstreamStackBusLane [22][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[22][31].cb_test                                      ;
                vDownstreamStackBusLane [22][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [22][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[23][0].cb_test                                      ;
                vDownstreamStackBusLane [23][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][1].cb_test                                      ;
                vDownstreamStackBusLane [23][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][2].cb_test                                      ;
                vDownstreamStackBusLane [23][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][3].cb_test                                      ;
                vDownstreamStackBusLane [23][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][4].cb_test                                      ;
                vDownstreamStackBusLane [23][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][5].cb_test                                      ;
                vDownstreamStackBusLane [23][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][6].cb_test                                      ;
                vDownstreamStackBusLane [23][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][7].cb_test                                      ;
                vDownstreamStackBusLane [23][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][8].cb_test                                      ;
                vDownstreamStackBusLane [23][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][9].cb_test                                      ;
                vDownstreamStackBusLane [23][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][10].cb_test                                      ;
                vDownstreamStackBusLane [23][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][11].cb_test                                      ;
                vDownstreamStackBusLane [23][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][12].cb_test                                      ;
                vDownstreamStackBusLane [23][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][13].cb_test                                      ;
                vDownstreamStackBusLane [23][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][14].cb_test                                      ;
                vDownstreamStackBusLane [23][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][15].cb_test                                      ;
                vDownstreamStackBusLane [23][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][16].cb_test                                      ;
                vDownstreamStackBusLane [23][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][17].cb_test                                      ;
                vDownstreamStackBusLane [23][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][18].cb_test                                      ;
                vDownstreamStackBusLane [23][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][19].cb_test                                      ;
                vDownstreamStackBusLane [23][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][20].cb_test                                      ;
                vDownstreamStackBusLane [23][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][21].cb_test                                      ;
                vDownstreamStackBusLane [23][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][22].cb_test                                      ;
                vDownstreamStackBusLane [23][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][23].cb_test                                      ;
                vDownstreamStackBusLane [23][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][24].cb_test                                      ;
                vDownstreamStackBusLane [23][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][25].cb_test                                      ;
                vDownstreamStackBusLane [23][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][26].cb_test                                      ;
                vDownstreamStackBusLane [23][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][27].cb_test                                      ;
                vDownstreamStackBusLane [23][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][28].cb_test                                      ;
                vDownstreamStackBusLane [23][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][29].cb_test                                      ;
                vDownstreamStackBusLane [23][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][30].cb_test                                      ;
                vDownstreamStackBusLane [23][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[23][31].cb_test                                      ;
                vDownstreamStackBusLane [23][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [23][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[24][0].cb_test                                      ;
                vDownstreamStackBusLane [24][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][1].cb_test                                      ;
                vDownstreamStackBusLane [24][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][2].cb_test                                      ;
                vDownstreamStackBusLane [24][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][3].cb_test                                      ;
                vDownstreamStackBusLane [24][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][4].cb_test                                      ;
                vDownstreamStackBusLane [24][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][5].cb_test                                      ;
                vDownstreamStackBusLane [24][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][6].cb_test                                      ;
                vDownstreamStackBusLane [24][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][7].cb_test                                      ;
                vDownstreamStackBusLane [24][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][8].cb_test                                      ;
                vDownstreamStackBusLane [24][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][9].cb_test                                      ;
                vDownstreamStackBusLane [24][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][10].cb_test                                      ;
                vDownstreamStackBusLane [24][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][11].cb_test                                      ;
                vDownstreamStackBusLane [24][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][12].cb_test                                      ;
                vDownstreamStackBusLane [24][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][13].cb_test                                      ;
                vDownstreamStackBusLane [24][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][14].cb_test                                      ;
                vDownstreamStackBusLane [24][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][15].cb_test                                      ;
                vDownstreamStackBusLane [24][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][16].cb_test                                      ;
                vDownstreamStackBusLane [24][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][17].cb_test                                      ;
                vDownstreamStackBusLane [24][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][18].cb_test                                      ;
                vDownstreamStackBusLane [24][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][19].cb_test                                      ;
                vDownstreamStackBusLane [24][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][20].cb_test                                      ;
                vDownstreamStackBusLane [24][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][21].cb_test                                      ;
                vDownstreamStackBusLane [24][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][22].cb_test                                      ;
                vDownstreamStackBusLane [24][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][23].cb_test                                      ;
                vDownstreamStackBusLane [24][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][24].cb_test                                      ;
                vDownstreamStackBusLane [24][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][25].cb_test                                      ;
                vDownstreamStackBusLane [24][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][26].cb_test                                      ;
                vDownstreamStackBusLane [24][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][27].cb_test                                      ;
                vDownstreamStackBusLane [24][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][28].cb_test                                      ;
                vDownstreamStackBusLane [24][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][29].cb_test                                      ;
                vDownstreamStackBusLane [24][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][30].cb_test                                      ;
                vDownstreamStackBusLane [24][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[24][31].cb_test                                      ;
                vDownstreamStackBusLane [24][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [24][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[25][0].cb_test                                      ;
                vDownstreamStackBusLane [25][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][1].cb_test                                      ;
                vDownstreamStackBusLane [25][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][2].cb_test                                      ;
                vDownstreamStackBusLane [25][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][3].cb_test                                      ;
                vDownstreamStackBusLane [25][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][4].cb_test                                      ;
                vDownstreamStackBusLane [25][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][5].cb_test                                      ;
                vDownstreamStackBusLane [25][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][6].cb_test                                      ;
                vDownstreamStackBusLane [25][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][7].cb_test                                      ;
                vDownstreamStackBusLane [25][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][8].cb_test                                      ;
                vDownstreamStackBusLane [25][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][9].cb_test                                      ;
                vDownstreamStackBusLane [25][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][10].cb_test                                      ;
                vDownstreamStackBusLane [25][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][11].cb_test                                      ;
                vDownstreamStackBusLane [25][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][12].cb_test                                      ;
                vDownstreamStackBusLane [25][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][13].cb_test                                      ;
                vDownstreamStackBusLane [25][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][14].cb_test                                      ;
                vDownstreamStackBusLane [25][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][15].cb_test                                      ;
                vDownstreamStackBusLane [25][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][16].cb_test                                      ;
                vDownstreamStackBusLane [25][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][17].cb_test                                      ;
                vDownstreamStackBusLane [25][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][18].cb_test                                      ;
                vDownstreamStackBusLane [25][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][19].cb_test                                      ;
                vDownstreamStackBusLane [25][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][20].cb_test                                      ;
                vDownstreamStackBusLane [25][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][21].cb_test                                      ;
                vDownstreamStackBusLane [25][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][22].cb_test                                      ;
                vDownstreamStackBusLane [25][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][23].cb_test                                      ;
                vDownstreamStackBusLane [25][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][24].cb_test                                      ;
                vDownstreamStackBusLane [25][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][25].cb_test                                      ;
                vDownstreamStackBusLane [25][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][26].cb_test                                      ;
                vDownstreamStackBusLane [25][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][27].cb_test                                      ;
                vDownstreamStackBusLane [25][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][28].cb_test                                      ;
                vDownstreamStackBusLane [25][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][29].cb_test                                      ;
                vDownstreamStackBusLane [25][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][30].cb_test                                      ;
                vDownstreamStackBusLane [25][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[25][31].cb_test                                      ;
                vDownstreamStackBusLane [25][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [25][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[26][0].cb_test                                      ;
                vDownstreamStackBusLane [26][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][1].cb_test                                      ;
                vDownstreamStackBusLane [26][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][2].cb_test                                      ;
                vDownstreamStackBusLane [26][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][3].cb_test                                      ;
                vDownstreamStackBusLane [26][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][4].cb_test                                      ;
                vDownstreamStackBusLane [26][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][5].cb_test                                      ;
                vDownstreamStackBusLane [26][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][6].cb_test                                      ;
                vDownstreamStackBusLane [26][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][7].cb_test                                      ;
                vDownstreamStackBusLane [26][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][8].cb_test                                      ;
                vDownstreamStackBusLane [26][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][9].cb_test                                      ;
                vDownstreamStackBusLane [26][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][10].cb_test                                      ;
                vDownstreamStackBusLane [26][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][11].cb_test                                      ;
                vDownstreamStackBusLane [26][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][12].cb_test                                      ;
                vDownstreamStackBusLane [26][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][13].cb_test                                      ;
                vDownstreamStackBusLane [26][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][14].cb_test                                      ;
                vDownstreamStackBusLane [26][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][15].cb_test                                      ;
                vDownstreamStackBusLane [26][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][16].cb_test                                      ;
                vDownstreamStackBusLane [26][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][17].cb_test                                      ;
                vDownstreamStackBusLane [26][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][18].cb_test                                      ;
                vDownstreamStackBusLane [26][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][19].cb_test                                      ;
                vDownstreamStackBusLane [26][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][20].cb_test                                      ;
                vDownstreamStackBusLane [26][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][21].cb_test                                      ;
                vDownstreamStackBusLane [26][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][22].cb_test                                      ;
                vDownstreamStackBusLane [26][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][23].cb_test                                      ;
                vDownstreamStackBusLane [26][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][24].cb_test                                      ;
                vDownstreamStackBusLane [26][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][25].cb_test                                      ;
                vDownstreamStackBusLane [26][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][26].cb_test                                      ;
                vDownstreamStackBusLane [26][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][27].cb_test                                      ;
                vDownstreamStackBusLane [26][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][28].cb_test                                      ;
                vDownstreamStackBusLane [26][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][29].cb_test                                      ;
                vDownstreamStackBusLane [26][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][30].cb_test                                      ;
                vDownstreamStackBusLane [26][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[26][31].cb_test                                      ;
                vDownstreamStackBusLane [26][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [26][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[27][0].cb_test                                      ;
                vDownstreamStackBusLane [27][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][1].cb_test                                      ;
                vDownstreamStackBusLane [27][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][2].cb_test                                      ;
                vDownstreamStackBusLane [27][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][3].cb_test                                      ;
                vDownstreamStackBusLane [27][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][4].cb_test                                      ;
                vDownstreamStackBusLane [27][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][5].cb_test                                      ;
                vDownstreamStackBusLane [27][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][6].cb_test                                      ;
                vDownstreamStackBusLane [27][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][7].cb_test                                      ;
                vDownstreamStackBusLane [27][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][8].cb_test                                      ;
                vDownstreamStackBusLane [27][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][9].cb_test                                      ;
                vDownstreamStackBusLane [27][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][10].cb_test                                      ;
                vDownstreamStackBusLane [27][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][11].cb_test                                      ;
                vDownstreamStackBusLane [27][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][12].cb_test                                      ;
                vDownstreamStackBusLane [27][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][13].cb_test                                      ;
                vDownstreamStackBusLane [27][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][14].cb_test                                      ;
                vDownstreamStackBusLane [27][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][15].cb_test                                      ;
                vDownstreamStackBusLane [27][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][16].cb_test                                      ;
                vDownstreamStackBusLane [27][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][17].cb_test                                      ;
                vDownstreamStackBusLane [27][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][18].cb_test                                      ;
                vDownstreamStackBusLane [27][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][19].cb_test                                      ;
                vDownstreamStackBusLane [27][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][20].cb_test                                      ;
                vDownstreamStackBusLane [27][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][21].cb_test                                      ;
                vDownstreamStackBusLane [27][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][22].cb_test                                      ;
                vDownstreamStackBusLane [27][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][23].cb_test                                      ;
                vDownstreamStackBusLane [27][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][24].cb_test                                      ;
                vDownstreamStackBusLane [27][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][25].cb_test                                      ;
                vDownstreamStackBusLane [27][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][26].cb_test                                      ;
                vDownstreamStackBusLane [27][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][27].cb_test                                      ;
                vDownstreamStackBusLane [27][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][28].cb_test                                      ;
                vDownstreamStackBusLane [27][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][29].cb_test                                      ;
                vDownstreamStackBusLane [27][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][30].cb_test                                      ;
                vDownstreamStackBusLane [27][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[27][31].cb_test                                      ;
                vDownstreamStackBusLane [27][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [27][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[28][0].cb_test                                      ;
                vDownstreamStackBusLane [28][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][1].cb_test                                      ;
                vDownstreamStackBusLane [28][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][2].cb_test                                      ;
                vDownstreamStackBusLane [28][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][3].cb_test                                      ;
                vDownstreamStackBusLane [28][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][4].cb_test                                      ;
                vDownstreamStackBusLane [28][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][5].cb_test                                      ;
                vDownstreamStackBusLane [28][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][6].cb_test                                      ;
                vDownstreamStackBusLane [28][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][7].cb_test                                      ;
                vDownstreamStackBusLane [28][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][8].cb_test                                      ;
                vDownstreamStackBusLane [28][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][9].cb_test                                      ;
                vDownstreamStackBusLane [28][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][10].cb_test                                      ;
                vDownstreamStackBusLane [28][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][11].cb_test                                      ;
                vDownstreamStackBusLane [28][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][12].cb_test                                      ;
                vDownstreamStackBusLane [28][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][13].cb_test                                      ;
                vDownstreamStackBusLane [28][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][14].cb_test                                      ;
                vDownstreamStackBusLane [28][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][15].cb_test                                      ;
                vDownstreamStackBusLane [28][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][16].cb_test                                      ;
                vDownstreamStackBusLane [28][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][17].cb_test                                      ;
                vDownstreamStackBusLane [28][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][18].cb_test                                      ;
                vDownstreamStackBusLane [28][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][19].cb_test                                      ;
                vDownstreamStackBusLane [28][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][20].cb_test                                      ;
                vDownstreamStackBusLane [28][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][21].cb_test                                      ;
                vDownstreamStackBusLane [28][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][22].cb_test                                      ;
                vDownstreamStackBusLane [28][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][23].cb_test                                      ;
                vDownstreamStackBusLane [28][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][24].cb_test                                      ;
                vDownstreamStackBusLane [28][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][25].cb_test                                      ;
                vDownstreamStackBusLane [28][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][26].cb_test                                      ;
                vDownstreamStackBusLane [28][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][27].cb_test                                      ;
                vDownstreamStackBusLane [28][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][28].cb_test                                      ;
                vDownstreamStackBusLane [28][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][29].cb_test                                      ;
                vDownstreamStackBusLane [28][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][30].cb_test                                      ;
                vDownstreamStackBusLane [28][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[28][31].cb_test                                      ;
                vDownstreamStackBusLane [28][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [28][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[29][0].cb_test                                      ;
                vDownstreamStackBusLane [29][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][1].cb_test                                      ;
                vDownstreamStackBusLane [29][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][2].cb_test                                      ;
                vDownstreamStackBusLane [29][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][3].cb_test                                      ;
                vDownstreamStackBusLane [29][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][4].cb_test                                      ;
                vDownstreamStackBusLane [29][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][5].cb_test                                      ;
                vDownstreamStackBusLane [29][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][6].cb_test                                      ;
                vDownstreamStackBusLane [29][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][7].cb_test                                      ;
                vDownstreamStackBusLane [29][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][8].cb_test                                      ;
                vDownstreamStackBusLane [29][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][9].cb_test                                      ;
                vDownstreamStackBusLane [29][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][10].cb_test                                      ;
                vDownstreamStackBusLane [29][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][11].cb_test                                      ;
                vDownstreamStackBusLane [29][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][12].cb_test                                      ;
                vDownstreamStackBusLane [29][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][13].cb_test                                      ;
                vDownstreamStackBusLane [29][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][14].cb_test                                      ;
                vDownstreamStackBusLane [29][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][15].cb_test                                      ;
                vDownstreamStackBusLane [29][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][16].cb_test                                      ;
                vDownstreamStackBusLane [29][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][17].cb_test                                      ;
                vDownstreamStackBusLane [29][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][18].cb_test                                      ;
                vDownstreamStackBusLane [29][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][19].cb_test                                      ;
                vDownstreamStackBusLane [29][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][20].cb_test                                      ;
                vDownstreamStackBusLane [29][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][21].cb_test                                      ;
                vDownstreamStackBusLane [29][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][22].cb_test                                      ;
                vDownstreamStackBusLane [29][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][23].cb_test                                      ;
                vDownstreamStackBusLane [29][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][24].cb_test                                      ;
                vDownstreamStackBusLane [29][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][25].cb_test                                      ;
                vDownstreamStackBusLane [29][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][26].cb_test                                      ;
                vDownstreamStackBusLane [29][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][27].cb_test                                      ;
                vDownstreamStackBusLane [29][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][28].cb_test                                      ;
                vDownstreamStackBusLane [29][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][29].cb_test                                      ;
                vDownstreamStackBusLane [29][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][30].cb_test                                      ;
                vDownstreamStackBusLane [29][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[29][31].cb_test                                      ;
                vDownstreamStackBusLane [29][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [29][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[30][0].cb_test                                      ;
                vDownstreamStackBusLane [30][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][1].cb_test                                      ;
                vDownstreamStackBusLane [30][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][2].cb_test                                      ;
                vDownstreamStackBusLane [30][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][3].cb_test                                      ;
                vDownstreamStackBusLane [30][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][4].cb_test                                      ;
                vDownstreamStackBusLane [30][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][5].cb_test                                      ;
                vDownstreamStackBusLane [30][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][6].cb_test                                      ;
                vDownstreamStackBusLane [30][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][7].cb_test                                      ;
                vDownstreamStackBusLane [30][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][8].cb_test                                      ;
                vDownstreamStackBusLane [30][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][9].cb_test                                      ;
                vDownstreamStackBusLane [30][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][10].cb_test                                      ;
                vDownstreamStackBusLane [30][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][11].cb_test                                      ;
                vDownstreamStackBusLane [30][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][12].cb_test                                      ;
                vDownstreamStackBusLane [30][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][13].cb_test                                      ;
                vDownstreamStackBusLane [30][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][14].cb_test                                      ;
                vDownstreamStackBusLane [30][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][15].cb_test                                      ;
                vDownstreamStackBusLane [30][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][16].cb_test                                      ;
                vDownstreamStackBusLane [30][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][17].cb_test                                      ;
                vDownstreamStackBusLane [30][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][18].cb_test                                      ;
                vDownstreamStackBusLane [30][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][19].cb_test                                      ;
                vDownstreamStackBusLane [30][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][20].cb_test                                      ;
                vDownstreamStackBusLane [30][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][21].cb_test                                      ;
                vDownstreamStackBusLane [30][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][22].cb_test                                      ;
                vDownstreamStackBusLane [30][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][23].cb_test                                      ;
                vDownstreamStackBusLane [30][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][24].cb_test                                      ;
                vDownstreamStackBusLane [30][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][25].cb_test                                      ;
                vDownstreamStackBusLane [30][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][26].cb_test                                      ;
                vDownstreamStackBusLane [30][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][27].cb_test                                      ;
                vDownstreamStackBusLane [30][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][28].cb_test                                      ;
                vDownstreamStackBusLane [30][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][29].cb_test                                      ;
                vDownstreamStackBusLane [30][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][30].cb_test                                      ;
                vDownstreamStackBusLane [30][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[30][31].cb_test                                      ;
                vDownstreamStackBusLane [30][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [30][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[31][0].cb_test                                      ;
                vDownstreamStackBusLane [31][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][1].cb_test                                      ;
                vDownstreamStackBusLane [31][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][2].cb_test                                      ;
                vDownstreamStackBusLane [31][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][3].cb_test                                      ;
                vDownstreamStackBusLane [31][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][4].cb_test                                      ;
                vDownstreamStackBusLane [31][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][5].cb_test                                      ;
                vDownstreamStackBusLane [31][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][6].cb_test                                      ;
                vDownstreamStackBusLane [31][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][7].cb_test                                      ;
                vDownstreamStackBusLane [31][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][8].cb_test                                      ;
                vDownstreamStackBusLane [31][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][9].cb_test                                      ;
                vDownstreamStackBusLane [31][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][10].cb_test                                      ;
                vDownstreamStackBusLane [31][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][11].cb_test                                      ;
                vDownstreamStackBusLane [31][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][12].cb_test                                      ;
                vDownstreamStackBusLane [31][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][13].cb_test                                      ;
                vDownstreamStackBusLane [31][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][14].cb_test                                      ;
                vDownstreamStackBusLane [31][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][15].cb_test                                      ;
                vDownstreamStackBusLane [31][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][16].cb_test                                      ;
                vDownstreamStackBusLane [31][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][17].cb_test                                      ;
                vDownstreamStackBusLane [31][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][18].cb_test                                      ;
                vDownstreamStackBusLane [31][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][19].cb_test                                      ;
                vDownstreamStackBusLane [31][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][20].cb_test                                      ;
                vDownstreamStackBusLane [31][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][21].cb_test                                      ;
                vDownstreamStackBusLane [31][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][22].cb_test                                      ;
                vDownstreamStackBusLane [31][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][23].cb_test                                      ;
                vDownstreamStackBusLane [31][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][24].cb_test                                      ;
                vDownstreamStackBusLane [31][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][25].cb_test                                      ;
                vDownstreamStackBusLane [31][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][26].cb_test                                      ;
                vDownstreamStackBusLane [31][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][27].cb_test                                      ;
                vDownstreamStackBusLane [31][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][28].cb_test                                      ;
                vDownstreamStackBusLane [31][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][29].cb_test                                      ;
                vDownstreamStackBusLane [31][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][30].cb_test                                      ;
                vDownstreamStackBusLane [31][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[31][31].cb_test                                      ;
                vDownstreamStackBusLane [31][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [31][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[32][0].cb_test                                      ;
                vDownstreamStackBusLane [32][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][1].cb_test                                      ;
                vDownstreamStackBusLane [32][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][2].cb_test                                      ;
                vDownstreamStackBusLane [32][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][3].cb_test                                      ;
                vDownstreamStackBusLane [32][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][4].cb_test                                      ;
                vDownstreamStackBusLane [32][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][5].cb_test                                      ;
                vDownstreamStackBusLane [32][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][6].cb_test                                      ;
                vDownstreamStackBusLane [32][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][7].cb_test                                      ;
                vDownstreamStackBusLane [32][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][8].cb_test                                      ;
                vDownstreamStackBusLane [32][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][9].cb_test                                      ;
                vDownstreamStackBusLane [32][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][10].cb_test                                      ;
                vDownstreamStackBusLane [32][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][11].cb_test                                      ;
                vDownstreamStackBusLane [32][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][12].cb_test                                      ;
                vDownstreamStackBusLane [32][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][13].cb_test                                      ;
                vDownstreamStackBusLane [32][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][14].cb_test                                      ;
                vDownstreamStackBusLane [32][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][15].cb_test                                      ;
                vDownstreamStackBusLane [32][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][16].cb_test                                      ;
                vDownstreamStackBusLane [32][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][17].cb_test                                      ;
                vDownstreamStackBusLane [32][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][18].cb_test                                      ;
                vDownstreamStackBusLane [32][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][19].cb_test                                      ;
                vDownstreamStackBusLane [32][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][20].cb_test                                      ;
                vDownstreamStackBusLane [32][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][21].cb_test                                      ;
                vDownstreamStackBusLane [32][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][22].cb_test                                      ;
                vDownstreamStackBusLane [32][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][23].cb_test                                      ;
                vDownstreamStackBusLane [32][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][24].cb_test                                      ;
                vDownstreamStackBusLane [32][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][25].cb_test                                      ;
                vDownstreamStackBusLane [32][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][26].cb_test                                      ;
                vDownstreamStackBusLane [32][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][27].cb_test                                      ;
                vDownstreamStackBusLane [32][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][28].cb_test                                      ;
                vDownstreamStackBusLane [32][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][29].cb_test                                      ;
                vDownstreamStackBusLane [32][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][30].cb_test                                      ;
                vDownstreamStackBusLane [32][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[32][31].cb_test                                      ;
                vDownstreamStackBusLane [32][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [32][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[33][0].cb_test                                      ;
                vDownstreamStackBusLane [33][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][1].cb_test                                      ;
                vDownstreamStackBusLane [33][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][2].cb_test                                      ;
                vDownstreamStackBusLane [33][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][3].cb_test                                      ;
                vDownstreamStackBusLane [33][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][4].cb_test                                      ;
                vDownstreamStackBusLane [33][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][5].cb_test                                      ;
                vDownstreamStackBusLane [33][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][6].cb_test                                      ;
                vDownstreamStackBusLane [33][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][7].cb_test                                      ;
                vDownstreamStackBusLane [33][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][8].cb_test                                      ;
                vDownstreamStackBusLane [33][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][9].cb_test                                      ;
                vDownstreamStackBusLane [33][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][10].cb_test                                      ;
                vDownstreamStackBusLane [33][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][11].cb_test                                      ;
                vDownstreamStackBusLane [33][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][12].cb_test                                      ;
                vDownstreamStackBusLane [33][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][13].cb_test                                      ;
                vDownstreamStackBusLane [33][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][14].cb_test                                      ;
                vDownstreamStackBusLane [33][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][15].cb_test                                      ;
                vDownstreamStackBusLane [33][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][16].cb_test                                      ;
                vDownstreamStackBusLane [33][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][17].cb_test                                      ;
                vDownstreamStackBusLane [33][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][18].cb_test                                      ;
                vDownstreamStackBusLane [33][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][19].cb_test                                      ;
                vDownstreamStackBusLane [33][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][20].cb_test                                      ;
                vDownstreamStackBusLane [33][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][21].cb_test                                      ;
                vDownstreamStackBusLane [33][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][22].cb_test                                      ;
                vDownstreamStackBusLane [33][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][23].cb_test                                      ;
                vDownstreamStackBusLane [33][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][24].cb_test                                      ;
                vDownstreamStackBusLane [33][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][25].cb_test                                      ;
                vDownstreamStackBusLane [33][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][26].cb_test                                      ;
                vDownstreamStackBusLane [33][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][27].cb_test                                      ;
                vDownstreamStackBusLane [33][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][28].cb_test                                      ;
                vDownstreamStackBusLane [33][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][29].cb_test                                      ;
                vDownstreamStackBusLane [33][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][30].cb_test                                      ;
                vDownstreamStackBusLane [33][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[33][31].cb_test                                      ;
                vDownstreamStackBusLane [33][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [33][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[34][0].cb_test                                      ;
                vDownstreamStackBusLane [34][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][1].cb_test                                      ;
                vDownstreamStackBusLane [34][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][2].cb_test                                      ;
                vDownstreamStackBusLane [34][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][3].cb_test                                      ;
                vDownstreamStackBusLane [34][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][4].cb_test                                      ;
                vDownstreamStackBusLane [34][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][5].cb_test                                      ;
                vDownstreamStackBusLane [34][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][6].cb_test                                      ;
                vDownstreamStackBusLane [34][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][7].cb_test                                      ;
                vDownstreamStackBusLane [34][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][8].cb_test                                      ;
                vDownstreamStackBusLane [34][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][9].cb_test                                      ;
                vDownstreamStackBusLane [34][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][10].cb_test                                      ;
                vDownstreamStackBusLane [34][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][11].cb_test                                      ;
                vDownstreamStackBusLane [34][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][12].cb_test                                      ;
                vDownstreamStackBusLane [34][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][13].cb_test                                      ;
                vDownstreamStackBusLane [34][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][14].cb_test                                      ;
                vDownstreamStackBusLane [34][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][15].cb_test                                      ;
                vDownstreamStackBusLane [34][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][16].cb_test                                      ;
                vDownstreamStackBusLane [34][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][17].cb_test                                      ;
                vDownstreamStackBusLane [34][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][18].cb_test                                      ;
                vDownstreamStackBusLane [34][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][19].cb_test                                      ;
                vDownstreamStackBusLane [34][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][20].cb_test                                      ;
                vDownstreamStackBusLane [34][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][21].cb_test                                      ;
                vDownstreamStackBusLane [34][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][22].cb_test                                      ;
                vDownstreamStackBusLane [34][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][23].cb_test                                      ;
                vDownstreamStackBusLane [34][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][24].cb_test                                      ;
                vDownstreamStackBusLane [34][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][25].cb_test                                      ;
                vDownstreamStackBusLane [34][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][26].cb_test                                      ;
                vDownstreamStackBusLane [34][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][27].cb_test                                      ;
                vDownstreamStackBusLane [34][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][28].cb_test                                      ;
                vDownstreamStackBusLane [34][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][29].cb_test                                      ;
                vDownstreamStackBusLane [34][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][30].cb_test                                      ;
                vDownstreamStackBusLane [34][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[34][31].cb_test                                      ;
                vDownstreamStackBusLane [34][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [34][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[35][0].cb_test                                      ;
                vDownstreamStackBusLane [35][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][1].cb_test                                      ;
                vDownstreamStackBusLane [35][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][2].cb_test                                      ;
                vDownstreamStackBusLane [35][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][3].cb_test                                      ;
                vDownstreamStackBusLane [35][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][4].cb_test                                      ;
                vDownstreamStackBusLane [35][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][5].cb_test                                      ;
                vDownstreamStackBusLane [35][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][6].cb_test                                      ;
                vDownstreamStackBusLane [35][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][7].cb_test                                      ;
                vDownstreamStackBusLane [35][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][8].cb_test                                      ;
                vDownstreamStackBusLane [35][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][9].cb_test                                      ;
                vDownstreamStackBusLane [35][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][10].cb_test                                      ;
                vDownstreamStackBusLane [35][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][11].cb_test                                      ;
                vDownstreamStackBusLane [35][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][12].cb_test                                      ;
                vDownstreamStackBusLane [35][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][13].cb_test                                      ;
                vDownstreamStackBusLane [35][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][14].cb_test                                      ;
                vDownstreamStackBusLane [35][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][15].cb_test                                      ;
                vDownstreamStackBusLane [35][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][16].cb_test                                      ;
                vDownstreamStackBusLane [35][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][17].cb_test                                      ;
                vDownstreamStackBusLane [35][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][18].cb_test                                      ;
                vDownstreamStackBusLane [35][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][19].cb_test                                      ;
                vDownstreamStackBusLane [35][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][20].cb_test                                      ;
                vDownstreamStackBusLane [35][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][21].cb_test                                      ;
                vDownstreamStackBusLane [35][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][22].cb_test                                      ;
                vDownstreamStackBusLane [35][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][23].cb_test                                      ;
                vDownstreamStackBusLane [35][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][24].cb_test                                      ;
                vDownstreamStackBusLane [35][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][25].cb_test                                      ;
                vDownstreamStackBusLane [35][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][26].cb_test                                      ;
                vDownstreamStackBusLane [35][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][27].cb_test                                      ;
                vDownstreamStackBusLane [35][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][28].cb_test                                      ;
                vDownstreamStackBusLane [35][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][29].cb_test                                      ;
                vDownstreamStackBusLane [35][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][30].cb_test                                      ;
                vDownstreamStackBusLane [35][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[35][31].cb_test                                      ;
                vDownstreamStackBusLane [35][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [35][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[36][0].cb_test                                      ;
                vDownstreamStackBusLane [36][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][1].cb_test                                      ;
                vDownstreamStackBusLane [36][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][2].cb_test                                      ;
                vDownstreamStackBusLane [36][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][3].cb_test                                      ;
                vDownstreamStackBusLane [36][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][4].cb_test                                      ;
                vDownstreamStackBusLane [36][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][5].cb_test                                      ;
                vDownstreamStackBusLane [36][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][6].cb_test                                      ;
                vDownstreamStackBusLane [36][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][7].cb_test                                      ;
                vDownstreamStackBusLane [36][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][8].cb_test                                      ;
                vDownstreamStackBusLane [36][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][9].cb_test                                      ;
                vDownstreamStackBusLane [36][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][10].cb_test                                      ;
                vDownstreamStackBusLane [36][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][11].cb_test                                      ;
                vDownstreamStackBusLane [36][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][12].cb_test                                      ;
                vDownstreamStackBusLane [36][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][13].cb_test                                      ;
                vDownstreamStackBusLane [36][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][14].cb_test                                      ;
                vDownstreamStackBusLane [36][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][15].cb_test                                      ;
                vDownstreamStackBusLane [36][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][16].cb_test                                      ;
                vDownstreamStackBusLane [36][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][17].cb_test                                      ;
                vDownstreamStackBusLane [36][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][18].cb_test                                      ;
                vDownstreamStackBusLane [36][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][19].cb_test                                      ;
                vDownstreamStackBusLane [36][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][20].cb_test                                      ;
                vDownstreamStackBusLane [36][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][21].cb_test                                      ;
                vDownstreamStackBusLane [36][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][22].cb_test                                      ;
                vDownstreamStackBusLane [36][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][23].cb_test                                      ;
                vDownstreamStackBusLane [36][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][24].cb_test                                      ;
                vDownstreamStackBusLane [36][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][25].cb_test                                      ;
                vDownstreamStackBusLane [36][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][26].cb_test                                      ;
                vDownstreamStackBusLane [36][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][27].cb_test                                      ;
                vDownstreamStackBusLane [36][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][28].cb_test                                      ;
                vDownstreamStackBusLane [36][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][29].cb_test                                      ;
                vDownstreamStackBusLane [36][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][30].cb_test                                      ;
                vDownstreamStackBusLane [36][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[36][31].cb_test                                      ;
                vDownstreamStackBusLane [36][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [36][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[37][0].cb_test                                      ;
                vDownstreamStackBusLane [37][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][1].cb_test                                      ;
                vDownstreamStackBusLane [37][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][2].cb_test                                      ;
                vDownstreamStackBusLane [37][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][3].cb_test                                      ;
                vDownstreamStackBusLane [37][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][4].cb_test                                      ;
                vDownstreamStackBusLane [37][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][5].cb_test                                      ;
                vDownstreamStackBusLane [37][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][6].cb_test                                      ;
                vDownstreamStackBusLane [37][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][7].cb_test                                      ;
                vDownstreamStackBusLane [37][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][8].cb_test                                      ;
                vDownstreamStackBusLane [37][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][9].cb_test                                      ;
                vDownstreamStackBusLane [37][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][10].cb_test                                      ;
                vDownstreamStackBusLane [37][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][11].cb_test                                      ;
                vDownstreamStackBusLane [37][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][12].cb_test                                      ;
                vDownstreamStackBusLane [37][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][13].cb_test                                      ;
                vDownstreamStackBusLane [37][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][14].cb_test                                      ;
                vDownstreamStackBusLane [37][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][15].cb_test                                      ;
                vDownstreamStackBusLane [37][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][16].cb_test                                      ;
                vDownstreamStackBusLane [37][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][17].cb_test                                      ;
                vDownstreamStackBusLane [37][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][18].cb_test                                      ;
                vDownstreamStackBusLane [37][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][19].cb_test                                      ;
                vDownstreamStackBusLane [37][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][20].cb_test                                      ;
                vDownstreamStackBusLane [37][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][21].cb_test                                      ;
                vDownstreamStackBusLane [37][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][22].cb_test                                      ;
                vDownstreamStackBusLane [37][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][23].cb_test                                      ;
                vDownstreamStackBusLane [37][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][24].cb_test                                      ;
                vDownstreamStackBusLane [37][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][25].cb_test                                      ;
                vDownstreamStackBusLane [37][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][26].cb_test                                      ;
                vDownstreamStackBusLane [37][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][27].cb_test                                      ;
                vDownstreamStackBusLane [37][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][28].cb_test                                      ;
                vDownstreamStackBusLane [37][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][29].cb_test                                      ;
                vDownstreamStackBusLane [37][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][30].cb_test                                      ;
                vDownstreamStackBusLane [37][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[37][31].cb_test                                      ;
                vDownstreamStackBusLane [37][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [37][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[38][0].cb_test                                      ;
                vDownstreamStackBusLane [38][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][1].cb_test                                      ;
                vDownstreamStackBusLane [38][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][2].cb_test                                      ;
                vDownstreamStackBusLane [38][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][3].cb_test                                      ;
                vDownstreamStackBusLane [38][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][4].cb_test                                      ;
                vDownstreamStackBusLane [38][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][5].cb_test                                      ;
                vDownstreamStackBusLane [38][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][6].cb_test                                      ;
                vDownstreamStackBusLane [38][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][7].cb_test                                      ;
                vDownstreamStackBusLane [38][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][8].cb_test                                      ;
                vDownstreamStackBusLane [38][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][9].cb_test                                      ;
                vDownstreamStackBusLane [38][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][10].cb_test                                      ;
                vDownstreamStackBusLane [38][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][11].cb_test                                      ;
                vDownstreamStackBusLane [38][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][12].cb_test                                      ;
                vDownstreamStackBusLane [38][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][13].cb_test                                      ;
                vDownstreamStackBusLane [38][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][14].cb_test                                      ;
                vDownstreamStackBusLane [38][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][15].cb_test                                      ;
                vDownstreamStackBusLane [38][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][16].cb_test                                      ;
                vDownstreamStackBusLane [38][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][17].cb_test                                      ;
                vDownstreamStackBusLane [38][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][18].cb_test                                      ;
                vDownstreamStackBusLane [38][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][19].cb_test                                      ;
                vDownstreamStackBusLane [38][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][20].cb_test                                      ;
                vDownstreamStackBusLane [38][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][21].cb_test                                      ;
                vDownstreamStackBusLane [38][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][22].cb_test                                      ;
                vDownstreamStackBusLane [38][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][23].cb_test                                      ;
                vDownstreamStackBusLane [38][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][24].cb_test                                      ;
                vDownstreamStackBusLane [38][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][25].cb_test                                      ;
                vDownstreamStackBusLane [38][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][26].cb_test                                      ;
                vDownstreamStackBusLane [38][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][27].cb_test                                      ;
                vDownstreamStackBusLane [38][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][28].cb_test                                      ;
                vDownstreamStackBusLane [38][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][29].cb_test                                      ;
                vDownstreamStackBusLane [38][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][30].cb_test                                      ;
                vDownstreamStackBusLane [38][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[38][31].cb_test                                      ;
                vDownstreamStackBusLane [38][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [38][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[39][0].cb_test                                      ;
                vDownstreamStackBusLane [39][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][1].cb_test                                      ;
                vDownstreamStackBusLane [39][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][2].cb_test                                      ;
                vDownstreamStackBusLane [39][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][3].cb_test                                      ;
                vDownstreamStackBusLane [39][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][4].cb_test                                      ;
                vDownstreamStackBusLane [39][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][5].cb_test                                      ;
                vDownstreamStackBusLane [39][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][6].cb_test                                      ;
                vDownstreamStackBusLane [39][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][7].cb_test                                      ;
                vDownstreamStackBusLane [39][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][8].cb_test                                      ;
                vDownstreamStackBusLane [39][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][9].cb_test                                      ;
                vDownstreamStackBusLane [39][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][10].cb_test                                      ;
                vDownstreamStackBusLane [39][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][11].cb_test                                      ;
                vDownstreamStackBusLane [39][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][12].cb_test                                      ;
                vDownstreamStackBusLane [39][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][13].cb_test                                      ;
                vDownstreamStackBusLane [39][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][14].cb_test                                      ;
                vDownstreamStackBusLane [39][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][15].cb_test                                      ;
                vDownstreamStackBusLane [39][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][16].cb_test                                      ;
                vDownstreamStackBusLane [39][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][17].cb_test                                      ;
                vDownstreamStackBusLane [39][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][18].cb_test                                      ;
                vDownstreamStackBusLane [39][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][19].cb_test                                      ;
                vDownstreamStackBusLane [39][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][20].cb_test                                      ;
                vDownstreamStackBusLane [39][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][21].cb_test                                      ;
                vDownstreamStackBusLane [39][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][22].cb_test                                      ;
                vDownstreamStackBusLane [39][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][23].cb_test                                      ;
                vDownstreamStackBusLane [39][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][24].cb_test                                      ;
                vDownstreamStackBusLane [39][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][25].cb_test                                      ;
                vDownstreamStackBusLane [39][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][26].cb_test                                      ;
                vDownstreamStackBusLane [39][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][27].cb_test                                      ;
                vDownstreamStackBusLane [39][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][28].cb_test                                      ;
                vDownstreamStackBusLane [39][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][29].cb_test                                      ;
                vDownstreamStackBusLane [39][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][30].cb_test                                      ;
                vDownstreamStackBusLane [39][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[39][31].cb_test                                      ;
                vDownstreamStackBusLane [39][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [39][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[40][0].cb_test                                      ;
                vDownstreamStackBusLane [40][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][1].cb_test                                      ;
                vDownstreamStackBusLane [40][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][2].cb_test                                      ;
                vDownstreamStackBusLane [40][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][3].cb_test                                      ;
                vDownstreamStackBusLane [40][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][4].cb_test                                      ;
                vDownstreamStackBusLane [40][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][5].cb_test                                      ;
                vDownstreamStackBusLane [40][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][6].cb_test                                      ;
                vDownstreamStackBusLane [40][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][7].cb_test                                      ;
                vDownstreamStackBusLane [40][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][8].cb_test                                      ;
                vDownstreamStackBusLane [40][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][9].cb_test                                      ;
                vDownstreamStackBusLane [40][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][10].cb_test                                      ;
                vDownstreamStackBusLane [40][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][11].cb_test                                      ;
                vDownstreamStackBusLane [40][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][12].cb_test                                      ;
                vDownstreamStackBusLane [40][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][13].cb_test                                      ;
                vDownstreamStackBusLane [40][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][14].cb_test                                      ;
                vDownstreamStackBusLane [40][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][15].cb_test                                      ;
                vDownstreamStackBusLane [40][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][16].cb_test                                      ;
                vDownstreamStackBusLane [40][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][17].cb_test                                      ;
                vDownstreamStackBusLane [40][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][18].cb_test                                      ;
                vDownstreamStackBusLane [40][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][19].cb_test                                      ;
                vDownstreamStackBusLane [40][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][20].cb_test                                      ;
                vDownstreamStackBusLane [40][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][21].cb_test                                      ;
                vDownstreamStackBusLane [40][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][22].cb_test                                      ;
                vDownstreamStackBusLane [40][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][23].cb_test                                      ;
                vDownstreamStackBusLane [40][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][24].cb_test                                      ;
                vDownstreamStackBusLane [40][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][25].cb_test                                      ;
                vDownstreamStackBusLane [40][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][26].cb_test                                      ;
                vDownstreamStackBusLane [40][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][27].cb_test                                      ;
                vDownstreamStackBusLane [40][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][28].cb_test                                      ;
                vDownstreamStackBusLane [40][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][29].cb_test                                      ;
                vDownstreamStackBusLane [40][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][30].cb_test                                      ;
                vDownstreamStackBusLane [40][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[40][31].cb_test                                      ;
                vDownstreamStackBusLane [40][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [40][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[41][0].cb_test                                      ;
                vDownstreamStackBusLane [41][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][1].cb_test                                      ;
                vDownstreamStackBusLane [41][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][2].cb_test                                      ;
                vDownstreamStackBusLane [41][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][3].cb_test                                      ;
                vDownstreamStackBusLane [41][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][4].cb_test                                      ;
                vDownstreamStackBusLane [41][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][5].cb_test                                      ;
                vDownstreamStackBusLane [41][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][6].cb_test                                      ;
                vDownstreamStackBusLane [41][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][7].cb_test                                      ;
                vDownstreamStackBusLane [41][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][8].cb_test                                      ;
                vDownstreamStackBusLane [41][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][9].cb_test                                      ;
                vDownstreamStackBusLane [41][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][10].cb_test                                      ;
                vDownstreamStackBusLane [41][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][11].cb_test                                      ;
                vDownstreamStackBusLane [41][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][12].cb_test                                      ;
                vDownstreamStackBusLane [41][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][13].cb_test                                      ;
                vDownstreamStackBusLane [41][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][14].cb_test                                      ;
                vDownstreamStackBusLane [41][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][15].cb_test                                      ;
                vDownstreamStackBusLane [41][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][16].cb_test                                      ;
                vDownstreamStackBusLane [41][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][17].cb_test                                      ;
                vDownstreamStackBusLane [41][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][18].cb_test                                      ;
                vDownstreamStackBusLane [41][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][19].cb_test                                      ;
                vDownstreamStackBusLane [41][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][20].cb_test                                      ;
                vDownstreamStackBusLane [41][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][21].cb_test                                      ;
                vDownstreamStackBusLane [41][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][22].cb_test                                      ;
                vDownstreamStackBusLane [41][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][23].cb_test                                      ;
                vDownstreamStackBusLane [41][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][24].cb_test                                      ;
                vDownstreamStackBusLane [41][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][25].cb_test                                      ;
                vDownstreamStackBusLane [41][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][26].cb_test                                      ;
                vDownstreamStackBusLane [41][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][27].cb_test                                      ;
                vDownstreamStackBusLane [41][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][28].cb_test                                      ;
                vDownstreamStackBusLane [41][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][29].cb_test                                      ;
                vDownstreamStackBusLane [41][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][30].cb_test                                      ;
                vDownstreamStackBusLane [41][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[41][31].cb_test                                      ;
                vDownstreamStackBusLane [41][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [41][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[42][0].cb_test                                      ;
                vDownstreamStackBusLane [42][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][1].cb_test                                      ;
                vDownstreamStackBusLane [42][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][2].cb_test                                      ;
                vDownstreamStackBusLane [42][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][3].cb_test                                      ;
                vDownstreamStackBusLane [42][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][4].cb_test                                      ;
                vDownstreamStackBusLane [42][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][5].cb_test                                      ;
                vDownstreamStackBusLane [42][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][6].cb_test                                      ;
                vDownstreamStackBusLane [42][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][7].cb_test                                      ;
                vDownstreamStackBusLane [42][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][8].cb_test                                      ;
                vDownstreamStackBusLane [42][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][9].cb_test                                      ;
                vDownstreamStackBusLane [42][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][10].cb_test                                      ;
                vDownstreamStackBusLane [42][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][11].cb_test                                      ;
                vDownstreamStackBusLane [42][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][12].cb_test                                      ;
                vDownstreamStackBusLane [42][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][13].cb_test                                      ;
                vDownstreamStackBusLane [42][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][14].cb_test                                      ;
                vDownstreamStackBusLane [42][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][15].cb_test                                      ;
                vDownstreamStackBusLane [42][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][16].cb_test                                      ;
                vDownstreamStackBusLane [42][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][17].cb_test                                      ;
                vDownstreamStackBusLane [42][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][18].cb_test                                      ;
                vDownstreamStackBusLane [42][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][19].cb_test                                      ;
                vDownstreamStackBusLane [42][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][20].cb_test                                      ;
                vDownstreamStackBusLane [42][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][21].cb_test                                      ;
                vDownstreamStackBusLane [42][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][22].cb_test                                      ;
                vDownstreamStackBusLane [42][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][23].cb_test                                      ;
                vDownstreamStackBusLane [42][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][24].cb_test                                      ;
                vDownstreamStackBusLane [42][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][25].cb_test                                      ;
                vDownstreamStackBusLane [42][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][26].cb_test                                      ;
                vDownstreamStackBusLane [42][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][27].cb_test                                      ;
                vDownstreamStackBusLane [42][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][28].cb_test                                      ;
                vDownstreamStackBusLane [42][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][29].cb_test                                      ;
                vDownstreamStackBusLane [42][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][30].cb_test                                      ;
                vDownstreamStackBusLane [42][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[42][31].cb_test                                      ;
                vDownstreamStackBusLane [42][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [42][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[43][0].cb_test                                      ;
                vDownstreamStackBusLane [43][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][1].cb_test                                      ;
                vDownstreamStackBusLane [43][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][2].cb_test                                      ;
                vDownstreamStackBusLane [43][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][3].cb_test                                      ;
                vDownstreamStackBusLane [43][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][4].cb_test                                      ;
                vDownstreamStackBusLane [43][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][5].cb_test                                      ;
                vDownstreamStackBusLane [43][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][6].cb_test                                      ;
                vDownstreamStackBusLane [43][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][7].cb_test                                      ;
                vDownstreamStackBusLane [43][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][8].cb_test                                      ;
                vDownstreamStackBusLane [43][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][9].cb_test                                      ;
                vDownstreamStackBusLane [43][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][10].cb_test                                      ;
                vDownstreamStackBusLane [43][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][11].cb_test                                      ;
                vDownstreamStackBusLane [43][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][12].cb_test                                      ;
                vDownstreamStackBusLane [43][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][13].cb_test                                      ;
                vDownstreamStackBusLane [43][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][14].cb_test                                      ;
                vDownstreamStackBusLane [43][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][15].cb_test                                      ;
                vDownstreamStackBusLane [43][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][16].cb_test                                      ;
                vDownstreamStackBusLane [43][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][17].cb_test                                      ;
                vDownstreamStackBusLane [43][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][18].cb_test                                      ;
                vDownstreamStackBusLane [43][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][19].cb_test                                      ;
                vDownstreamStackBusLane [43][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][20].cb_test                                      ;
                vDownstreamStackBusLane [43][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][21].cb_test                                      ;
                vDownstreamStackBusLane [43][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][22].cb_test                                      ;
                vDownstreamStackBusLane [43][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][23].cb_test                                      ;
                vDownstreamStackBusLane [43][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][24].cb_test                                      ;
                vDownstreamStackBusLane [43][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][25].cb_test                                      ;
                vDownstreamStackBusLane [43][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][26].cb_test                                      ;
                vDownstreamStackBusLane [43][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][27].cb_test                                      ;
                vDownstreamStackBusLane [43][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][28].cb_test                                      ;
                vDownstreamStackBusLane [43][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][29].cb_test                                      ;
                vDownstreamStackBusLane [43][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][30].cb_test                                      ;
                vDownstreamStackBusLane [43][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[43][31].cb_test                                      ;
                vDownstreamStackBusLane [43][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [43][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[44][0].cb_test                                      ;
                vDownstreamStackBusLane [44][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][1].cb_test                                      ;
                vDownstreamStackBusLane [44][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][2].cb_test                                      ;
                vDownstreamStackBusLane [44][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][3].cb_test                                      ;
                vDownstreamStackBusLane [44][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][4].cb_test                                      ;
                vDownstreamStackBusLane [44][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][5].cb_test                                      ;
                vDownstreamStackBusLane [44][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][6].cb_test                                      ;
                vDownstreamStackBusLane [44][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][7].cb_test                                      ;
                vDownstreamStackBusLane [44][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][8].cb_test                                      ;
                vDownstreamStackBusLane [44][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][9].cb_test                                      ;
                vDownstreamStackBusLane [44][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][10].cb_test                                      ;
                vDownstreamStackBusLane [44][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][11].cb_test                                      ;
                vDownstreamStackBusLane [44][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][12].cb_test                                      ;
                vDownstreamStackBusLane [44][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][13].cb_test                                      ;
                vDownstreamStackBusLane [44][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][14].cb_test                                      ;
                vDownstreamStackBusLane [44][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][15].cb_test                                      ;
                vDownstreamStackBusLane [44][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][16].cb_test                                      ;
                vDownstreamStackBusLane [44][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][17].cb_test                                      ;
                vDownstreamStackBusLane [44][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][18].cb_test                                      ;
                vDownstreamStackBusLane [44][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][19].cb_test                                      ;
                vDownstreamStackBusLane [44][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][20].cb_test                                      ;
                vDownstreamStackBusLane [44][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][21].cb_test                                      ;
                vDownstreamStackBusLane [44][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][22].cb_test                                      ;
                vDownstreamStackBusLane [44][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][23].cb_test                                      ;
                vDownstreamStackBusLane [44][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][24].cb_test                                      ;
                vDownstreamStackBusLane [44][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][25].cb_test                                      ;
                vDownstreamStackBusLane [44][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][26].cb_test                                      ;
                vDownstreamStackBusLane [44][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][27].cb_test                                      ;
                vDownstreamStackBusLane [44][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][28].cb_test                                      ;
                vDownstreamStackBusLane [44][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][29].cb_test                                      ;
                vDownstreamStackBusLane [44][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][30].cb_test                                      ;
                vDownstreamStackBusLane [44][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[44][31].cb_test                                      ;
                vDownstreamStackBusLane [44][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [44][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[45][0].cb_test                                      ;
                vDownstreamStackBusLane [45][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][1].cb_test                                      ;
                vDownstreamStackBusLane [45][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][2].cb_test                                      ;
                vDownstreamStackBusLane [45][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][3].cb_test                                      ;
                vDownstreamStackBusLane [45][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][4].cb_test                                      ;
                vDownstreamStackBusLane [45][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][5].cb_test                                      ;
                vDownstreamStackBusLane [45][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][6].cb_test                                      ;
                vDownstreamStackBusLane [45][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][7].cb_test                                      ;
                vDownstreamStackBusLane [45][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][8].cb_test                                      ;
                vDownstreamStackBusLane [45][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][9].cb_test                                      ;
                vDownstreamStackBusLane [45][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][10].cb_test                                      ;
                vDownstreamStackBusLane [45][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][11].cb_test                                      ;
                vDownstreamStackBusLane [45][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][12].cb_test                                      ;
                vDownstreamStackBusLane [45][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][13].cb_test                                      ;
                vDownstreamStackBusLane [45][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][14].cb_test                                      ;
                vDownstreamStackBusLane [45][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][15].cb_test                                      ;
                vDownstreamStackBusLane [45][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][16].cb_test                                      ;
                vDownstreamStackBusLane [45][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][17].cb_test                                      ;
                vDownstreamStackBusLane [45][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][18].cb_test                                      ;
                vDownstreamStackBusLane [45][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][19].cb_test                                      ;
                vDownstreamStackBusLane [45][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][20].cb_test                                      ;
                vDownstreamStackBusLane [45][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][21].cb_test                                      ;
                vDownstreamStackBusLane [45][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][22].cb_test                                      ;
                vDownstreamStackBusLane [45][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][23].cb_test                                      ;
                vDownstreamStackBusLane [45][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][24].cb_test                                      ;
                vDownstreamStackBusLane [45][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][25].cb_test                                      ;
                vDownstreamStackBusLane [45][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][26].cb_test                                      ;
                vDownstreamStackBusLane [45][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][27].cb_test                                      ;
                vDownstreamStackBusLane [45][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][28].cb_test                                      ;
                vDownstreamStackBusLane [45][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][29].cb_test                                      ;
                vDownstreamStackBusLane [45][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][30].cb_test                                      ;
                vDownstreamStackBusLane [45][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[45][31].cb_test                                      ;
                vDownstreamStackBusLane [45][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [45][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[46][0].cb_test                                      ;
                vDownstreamStackBusLane [46][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][1].cb_test                                      ;
                vDownstreamStackBusLane [46][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][2].cb_test                                      ;
                vDownstreamStackBusLane [46][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][3].cb_test                                      ;
                vDownstreamStackBusLane [46][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][4].cb_test                                      ;
                vDownstreamStackBusLane [46][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][5].cb_test                                      ;
                vDownstreamStackBusLane [46][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][6].cb_test                                      ;
                vDownstreamStackBusLane [46][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][7].cb_test                                      ;
                vDownstreamStackBusLane [46][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][8].cb_test                                      ;
                vDownstreamStackBusLane [46][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][9].cb_test                                      ;
                vDownstreamStackBusLane [46][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][10].cb_test                                      ;
                vDownstreamStackBusLane [46][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][11].cb_test                                      ;
                vDownstreamStackBusLane [46][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][12].cb_test                                      ;
                vDownstreamStackBusLane [46][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][13].cb_test                                      ;
                vDownstreamStackBusLane [46][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][14].cb_test                                      ;
                vDownstreamStackBusLane [46][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][15].cb_test                                      ;
                vDownstreamStackBusLane [46][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][16].cb_test                                      ;
                vDownstreamStackBusLane [46][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][17].cb_test                                      ;
                vDownstreamStackBusLane [46][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][18].cb_test                                      ;
                vDownstreamStackBusLane [46][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][19].cb_test                                      ;
                vDownstreamStackBusLane [46][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][20].cb_test                                      ;
                vDownstreamStackBusLane [46][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][21].cb_test                                      ;
                vDownstreamStackBusLane [46][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][22].cb_test                                      ;
                vDownstreamStackBusLane [46][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][23].cb_test                                      ;
                vDownstreamStackBusLane [46][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][24].cb_test                                      ;
                vDownstreamStackBusLane [46][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][25].cb_test                                      ;
                vDownstreamStackBusLane [46][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][26].cb_test                                      ;
                vDownstreamStackBusLane [46][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][27].cb_test                                      ;
                vDownstreamStackBusLane [46][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][28].cb_test                                      ;
                vDownstreamStackBusLane [46][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][29].cb_test                                      ;
                vDownstreamStackBusLane [46][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][30].cb_test                                      ;
                vDownstreamStackBusLane [46][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[46][31].cb_test                                      ;
                vDownstreamStackBusLane [46][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [46][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[47][0].cb_test                                      ;
                vDownstreamStackBusLane [47][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][1].cb_test                                      ;
                vDownstreamStackBusLane [47][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][2].cb_test                                      ;
                vDownstreamStackBusLane [47][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][3].cb_test                                      ;
                vDownstreamStackBusLane [47][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][4].cb_test                                      ;
                vDownstreamStackBusLane [47][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][5].cb_test                                      ;
                vDownstreamStackBusLane [47][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][6].cb_test                                      ;
                vDownstreamStackBusLane [47][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][7].cb_test                                      ;
                vDownstreamStackBusLane [47][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][8].cb_test                                      ;
                vDownstreamStackBusLane [47][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][9].cb_test                                      ;
                vDownstreamStackBusLane [47][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][10].cb_test                                      ;
                vDownstreamStackBusLane [47][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][11].cb_test                                      ;
                vDownstreamStackBusLane [47][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][12].cb_test                                      ;
                vDownstreamStackBusLane [47][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][13].cb_test                                      ;
                vDownstreamStackBusLane [47][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][14].cb_test                                      ;
                vDownstreamStackBusLane [47][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][15].cb_test                                      ;
                vDownstreamStackBusLane [47][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][16].cb_test                                      ;
                vDownstreamStackBusLane [47][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][17].cb_test                                      ;
                vDownstreamStackBusLane [47][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][18].cb_test                                      ;
                vDownstreamStackBusLane [47][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][19].cb_test                                      ;
                vDownstreamStackBusLane [47][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][20].cb_test                                      ;
                vDownstreamStackBusLane [47][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][21].cb_test                                      ;
                vDownstreamStackBusLane [47][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][22].cb_test                                      ;
                vDownstreamStackBusLane [47][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][23].cb_test                                      ;
                vDownstreamStackBusLane [47][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][24].cb_test                                      ;
                vDownstreamStackBusLane [47][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][25].cb_test                                      ;
                vDownstreamStackBusLane [47][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][26].cb_test                                      ;
                vDownstreamStackBusLane [47][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][27].cb_test                                      ;
                vDownstreamStackBusLane [47][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][28].cb_test                                      ;
                vDownstreamStackBusLane [47][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][29].cb_test                                      ;
                vDownstreamStackBusLane [47][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][30].cb_test                                      ;
                vDownstreamStackBusLane [47][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[47][31].cb_test                                      ;
                vDownstreamStackBusLane [47][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [47][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[48][0].cb_test                                      ;
                vDownstreamStackBusLane [48][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][1].cb_test                                      ;
                vDownstreamStackBusLane [48][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][2].cb_test                                      ;
                vDownstreamStackBusLane [48][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][3].cb_test                                      ;
                vDownstreamStackBusLane [48][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][4].cb_test                                      ;
                vDownstreamStackBusLane [48][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][5].cb_test                                      ;
                vDownstreamStackBusLane [48][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][6].cb_test                                      ;
                vDownstreamStackBusLane [48][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][7].cb_test                                      ;
                vDownstreamStackBusLane [48][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][8].cb_test                                      ;
                vDownstreamStackBusLane [48][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][9].cb_test                                      ;
                vDownstreamStackBusLane [48][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][10].cb_test                                      ;
                vDownstreamStackBusLane [48][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][11].cb_test                                      ;
                vDownstreamStackBusLane [48][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][12].cb_test                                      ;
                vDownstreamStackBusLane [48][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][13].cb_test                                      ;
                vDownstreamStackBusLane [48][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][14].cb_test                                      ;
                vDownstreamStackBusLane [48][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][15].cb_test                                      ;
                vDownstreamStackBusLane [48][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][16].cb_test                                      ;
                vDownstreamStackBusLane [48][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][17].cb_test                                      ;
                vDownstreamStackBusLane [48][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][18].cb_test                                      ;
                vDownstreamStackBusLane [48][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][19].cb_test                                      ;
                vDownstreamStackBusLane [48][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][20].cb_test                                      ;
                vDownstreamStackBusLane [48][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][21].cb_test                                      ;
                vDownstreamStackBusLane [48][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][22].cb_test                                      ;
                vDownstreamStackBusLane [48][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][23].cb_test                                      ;
                vDownstreamStackBusLane [48][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][24].cb_test                                      ;
                vDownstreamStackBusLane [48][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][25].cb_test                                      ;
                vDownstreamStackBusLane [48][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][26].cb_test                                      ;
                vDownstreamStackBusLane [48][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][27].cb_test                                      ;
                vDownstreamStackBusLane [48][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][28].cb_test                                      ;
                vDownstreamStackBusLane [48][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][29].cb_test                                      ;
                vDownstreamStackBusLane [48][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][30].cb_test                                      ;
                vDownstreamStackBusLane [48][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[48][31].cb_test                                      ;
                vDownstreamStackBusLane [48][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [48][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[49][0].cb_test                                      ;
                vDownstreamStackBusLane [49][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][1].cb_test                                      ;
                vDownstreamStackBusLane [49][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][2].cb_test                                      ;
                vDownstreamStackBusLane [49][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][3].cb_test                                      ;
                vDownstreamStackBusLane [49][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][4].cb_test                                      ;
                vDownstreamStackBusLane [49][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][5].cb_test                                      ;
                vDownstreamStackBusLane [49][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][6].cb_test                                      ;
                vDownstreamStackBusLane [49][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][7].cb_test                                      ;
                vDownstreamStackBusLane [49][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][8].cb_test                                      ;
                vDownstreamStackBusLane [49][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][9].cb_test                                      ;
                vDownstreamStackBusLane [49][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][10].cb_test                                      ;
                vDownstreamStackBusLane [49][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][11].cb_test                                      ;
                vDownstreamStackBusLane [49][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][12].cb_test                                      ;
                vDownstreamStackBusLane [49][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][13].cb_test                                      ;
                vDownstreamStackBusLane [49][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][14].cb_test                                      ;
                vDownstreamStackBusLane [49][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][15].cb_test                                      ;
                vDownstreamStackBusLane [49][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][16].cb_test                                      ;
                vDownstreamStackBusLane [49][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][17].cb_test                                      ;
                vDownstreamStackBusLane [49][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][18].cb_test                                      ;
                vDownstreamStackBusLane [49][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][19].cb_test                                      ;
                vDownstreamStackBusLane [49][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][20].cb_test                                      ;
                vDownstreamStackBusLane [49][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][21].cb_test                                      ;
                vDownstreamStackBusLane [49][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][22].cb_test                                      ;
                vDownstreamStackBusLane [49][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][23].cb_test                                      ;
                vDownstreamStackBusLane [49][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][24].cb_test                                      ;
                vDownstreamStackBusLane [49][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][25].cb_test                                      ;
                vDownstreamStackBusLane [49][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][26].cb_test                                      ;
                vDownstreamStackBusLane [49][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][27].cb_test                                      ;
                vDownstreamStackBusLane [49][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][28].cb_test                                      ;
                vDownstreamStackBusLane [49][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][29].cb_test                                      ;
                vDownstreamStackBusLane [49][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][30].cb_test                                      ;
                vDownstreamStackBusLane [49][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[49][31].cb_test                                      ;
                vDownstreamStackBusLane [49][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [49][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[50][0].cb_test                                      ;
                vDownstreamStackBusLane [50][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][1].cb_test                                      ;
                vDownstreamStackBusLane [50][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][2].cb_test                                      ;
                vDownstreamStackBusLane [50][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][3].cb_test                                      ;
                vDownstreamStackBusLane [50][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][4].cb_test                                      ;
                vDownstreamStackBusLane [50][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][5].cb_test                                      ;
                vDownstreamStackBusLane [50][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][6].cb_test                                      ;
                vDownstreamStackBusLane [50][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][7].cb_test                                      ;
                vDownstreamStackBusLane [50][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][8].cb_test                                      ;
                vDownstreamStackBusLane [50][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][9].cb_test                                      ;
                vDownstreamStackBusLane [50][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][10].cb_test                                      ;
                vDownstreamStackBusLane [50][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][11].cb_test                                      ;
                vDownstreamStackBusLane [50][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][12].cb_test                                      ;
                vDownstreamStackBusLane [50][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][13].cb_test                                      ;
                vDownstreamStackBusLane [50][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][14].cb_test                                      ;
                vDownstreamStackBusLane [50][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][15].cb_test                                      ;
                vDownstreamStackBusLane [50][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][16].cb_test                                      ;
                vDownstreamStackBusLane [50][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][17].cb_test                                      ;
                vDownstreamStackBusLane [50][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][18].cb_test                                      ;
                vDownstreamStackBusLane [50][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][19].cb_test                                      ;
                vDownstreamStackBusLane [50][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][20].cb_test                                      ;
                vDownstreamStackBusLane [50][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][21].cb_test                                      ;
                vDownstreamStackBusLane [50][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][22].cb_test                                      ;
                vDownstreamStackBusLane [50][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][23].cb_test                                      ;
                vDownstreamStackBusLane [50][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][24].cb_test                                      ;
                vDownstreamStackBusLane [50][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][25].cb_test                                      ;
                vDownstreamStackBusLane [50][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][26].cb_test                                      ;
                vDownstreamStackBusLane [50][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][27].cb_test                                      ;
                vDownstreamStackBusLane [50][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][28].cb_test                                      ;
                vDownstreamStackBusLane [50][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][29].cb_test                                      ;
                vDownstreamStackBusLane [50][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][30].cb_test                                      ;
                vDownstreamStackBusLane [50][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[50][31].cb_test                                      ;
                vDownstreamStackBusLane [50][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [50][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[51][0].cb_test                                      ;
                vDownstreamStackBusLane [51][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][1].cb_test                                      ;
                vDownstreamStackBusLane [51][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][2].cb_test                                      ;
                vDownstreamStackBusLane [51][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][3].cb_test                                      ;
                vDownstreamStackBusLane [51][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][4].cb_test                                      ;
                vDownstreamStackBusLane [51][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][5].cb_test                                      ;
                vDownstreamStackBusLane [51][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][6].cb_test                                      ;
                vDownstreamStackBusLane [51][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][7].cb_test                                      ;
                vDownstreamStackBusLane [51][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][8].cb_test                                      ;
                vDownstreamStackBusLane [51][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][9].cb_test                                      ;
                vDownstreamStackBusLane [51][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][10].cb_test                                      ;
                vDownstreamStackBusLane [51][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][11].cb_test                                      ;
                vDownstreamStackBusLane [51][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][12].cb_test                                      ;
                vDownstreamStackBusLane [51][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][13].cb_test                                      ;
                vDownstreamStackBusLane [51][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][14].cb_test                                      ;
                vDownstreamStackBusLane [51][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][15].cb_test                                      ;
                vDownstreamStackBusLane [51][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][16].cb_test                                      ;
                vDownstreamStackBusLane [51][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][17].cb_test                                      ;
                vDownstreamStackBusLane [51][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][18].cb_test                                      ;
                vDownstreamStackBusLane [51][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][19].cb_test                                      ;
                vDownstreamStackBusLane [51][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][20].cb_test                                      ;
                vDownstreamStackBusLane [51][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][21].cb_test                                      ;
                vDownstreamStackBusLane [51][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][22].cb_test                                      ;
                vDownstreamStackBusLane [51][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][23].cb_test                                      ;
                vDownstreamStackBusLane [51][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][24].cb_test                                      ;
                vDownstreamStackBusLane [51][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][25].cb_test                                      ;
                vDownstreamStackBusLane [51][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][26].cb_test                                      ;
                vDownstreamStackBusLane [51][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][27].cb_test                                      ;
                vDownstreamStackBusLane [51][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][28].cb_test                                      ;
                vDownstreamStackBusLane [51][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][29].cb_test                                      ;
                vDownstreamStackBusLane [51][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][30].cb_test                                      ;
                vDownstreamStackBusLane [51][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[51][31].cb_test                                      ;
                vDownstreamStackBusLane [51][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [51][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[52][0].cb_test                                      ;
                vDownstreamStackBusLane [52][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][1].cb_test                                      ;
                vDownstreamStackBusLane [52][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][2].cb_test                                      ;
                vDownstreamStackBusLane [52][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][3].cb_test                                      ;
                vDownstreamStackBusLane [52][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][4].cb_test                                      ;
                vDownstreamStackBusLane [52][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][5].cb_test                                      ;
                vDownstreamStackBusLane [52][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][6].cb_test                                      ;
                vDownstreamStackBusLane [52][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][7].cb_test                                      ;
                vDownstreamStackBusLane [52][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][8].cb_test                                      ;
                vDownstreamStackBusLane [52][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][9].cb_test                                      ;
                vDownstreamStackBusLane [52][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][10].cb_test                                      ;
                vDownstreamStackBusLane [52][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][11].cb_test                                      ;
                vDownstreamStackBusLane [52][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][12].cb_test                                      ;
                vDownstreamStackBusLane [52][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][13].cb_test                                      ;
                vDownstreamStackBusLane [52][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][14].cb_test                                      ;
                vDownstreamStackBusLane [52][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][15].cb_test                                      ;
                vDownstreamStackBusLane [52][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][16].cb_test                                      ;
                vDownstreamStackBusLane [52][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][17].cb_test                                      ;
                vDownstreamStackBusLane [52][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][18].cb_test                                      ;
                vDownstreamStackBusLane [52][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][19].cb_test                                      ;
                vDownstreamStackBusLane [52][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][20].cb_test                                      ;
                vDownstreamStackBusLane [52][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][21].cb_test                                      ;
                vDownstreamStackBusLane [52][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][22].cb_test                                      ;
                vDownstreamStackBusLane [52][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][23].cb_test                                      ;
                vDownstreamStackBusLane [52][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][24].cb_test                                      ;
                vDownstreamStackBusLane [52][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][25].cb_test                                      ;
                vDownstreamStackBusLane [52][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][26].cb_test                                      ;
                vDownstreamStackBusLane [52][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][27].cb_test                                      ;
                vDownstreamStackBusLane [52][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][28].cb_test                                      ;
                vDownstreamStackBusLane [52][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][29].cb_test                                      ;
                vDownstreamStackBusLane [52][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][30].cb_test                                      ;
                vDownstreamStackBusLane [52][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[52][31].cb_test                                      ;
                vDownstreamStackBusLane [52][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [52][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[53][0].cb_test                                      ;
                vDownstreamStackBusLane [53][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][1].cb_test                                      ;
                vDownstreamStackBusLane [53][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][2].cb_test                                      ;
                vDownstreamStackBusLane [53][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][3].cb_test                                      ;
                vDownstreamStackBusLane [53][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][4].cb_test                                      ;
                vDownstreamStackBusLane [53][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][5].cb_test                                      ;
                vDownstreamStackBusLane [53][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][6].cb_test                                      ;
                vDownstreamStackBusLane [53][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][7].cb_test                                      ;
                vDownstreamStackBusLane [53][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][8].cb_test                                      ;
                vDownstreamStackBusLane [53][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][9].cb_test                                      ;
                vDownstreamStackBusLane [53][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][10].cb_test                                      ;
                vDownstreamStackBusLane [53][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][11].cb_test                                      ;
                vDownstreamStackBusLane [53][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][12].cb_test                                      ;
                vDownstreamStackBusLane [53][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][13].cb_test                                      ;
                vDownstreamStackBusLane [53][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][14].cb_test                                      ;
                vDownstreamStackBusLane [53][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][15].cb_test                                      ;
                vDownstreamStackBusLane [53][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][16].cb_test                                      ;
                vDownstreamStackBusLane [53][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][17].cb_test                                      ;
                vDownstreamStackBusLane [53][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][18].cb_test                                      ;
                vDownstreamStackBusLane [53][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][19].cb_test                                      ;
                vDownstreamStackBusLane [53][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][20].cb_test                                      ;
                vDownstreamStackBusLane [53][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][21].cb_test                                      ;
                vDownstreamStackBusLane [53][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][22].cb_test                                      ;
                vDownstreamStackBusLane [53][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][23].cb_test                                      ;
                vDownstreamStackBusLane [53][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][24].cb_test                                      ;
                vDownstreamStackBusLane [53][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][25].cb_test                                      ;
                vDownstreamStackBusLane [53][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][26].cb_test                                      ;
                vDownstreamStackBusLane [53][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][27].cb_test                                      ;
                vDownstreamStackBusLane [53][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][28].cb_test                                      ;
                vDownstreamStackBusLane [53][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][29].cb_test                                      ;
                vDownstreamStackBusLane [53][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][30].cb_test                                      ;
                vDownstreamStackBusLane [53][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[53][31].cb_test                                      ;
                vDownstreamStackBusLane [53][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [53][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[54][0].cb_test                                      ;
                vDownstreamStackBusLane [54][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][1].cb_test                                      ;
                vDownstreamStackBusLane [54][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][2].cb_test                                      ;
                vDownstreamStackBusLane [54][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][3].cb_test                                      ;
                vDownstreamStackBusLane [54][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][4].cb_test                                      ;
                vDownstreamStackBusLane [54][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][5].cb_test                                      ;
                vDownstreamStackBusLane [54][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][6].cb_test                                      ;
                vDownstreamStackBusLane [54][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][7].cb_test                                      ;
                vDownstreamStackBusLane [54][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][8].cb_test                                      ;
                vDownstreamStackBusLane [54][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][9].cb_test                                      ;
                vDownstreamStackBusLane [54][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][10].cb_test                                      ;
                vDownstreamStackBusLane [54][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][11].cb_test                                      ;
                vDownstreamStackBusLane [54][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][12].cb_test                                      ;
                vDownstreamStackBusLane [54][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][13].cb_test                                      ;
                vDownstreamStackBusLane [54][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][14].cb_test                                      ;
                vDownstreamStackBusLane [54][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][15].cb_test                                      ;
                vDownstreamStackBusLane [54][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][16].cb_test                                      ;
                vDownstreamStackBusLane [54][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][17].cb_test                                      ;
                vDownstreamStackBusLane [54][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][18].cb_test                                      ;
                vDownstreamStackBusLane [54][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][19].cb_test                                      ;
                vDownstreamStackBusLane [54][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][20].cb_test                                      ;
                vDownstreamStackBusLane [54][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][21].cb_test                                      ;
                vDownstreamStackBusLane [54][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][22].cb_test                                      ;
                vDownstreamStackBusLane [54][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][23].cb_test                                      ;
                vDownstreamStackBusLane [54][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][24].cb_test                                      ;
                vDownstreamStackBusLane [54][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][25].cb_test                                      ;
                vDownstreamStackBusLane [54][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][26].cb_test                                      ;
                vDownstreamStackBusLane [54][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][27].cb_test                                      ;
                vDownstreamStackBusLane [54][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][28].cb_test                                      ;
                vDownstreamStackBusLane [54][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][29].cb_test                                      ;
                vDownstreamStackBusLane [54][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][30].cb_test                                      ;
                vDownstreamStackBusLane [54][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[54][31].cb_test                                      ;
                vDownstreamStackBusLane [54][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [54][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[55][0].cb_test                                      ;
                vDownstreamStackBusLane [55][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][1].cb_test                                      ;
                vDownstreamStackBusLane [55][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][2].cb_test                                      ;
                vDownstreamStackBusLane [55][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][3].cb_test                                      ;
                vDownstreamStackBusLane [55][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][4].cb_test                                      ;
                vDownstreamStackBusLane [55][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][5].cb_test                                      ;
                vDownstreamStackBusLane [55][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][6].cb_test                                      ;
                vDownstreamStackBusLane [55][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][7].cb_test                                      ;
                vDownstreamStackBusLane [55][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][8].cb_test                                      ;
                vDownstreamStackBusLane [55][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][9].cb_test                                      ;
                vDownstreamStackBusLane [55][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][10].cb_test                                      ;
                vDownstreamStackBusLane [55][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][11].cb_test                                      ;
                vDownstreamStackBusLane [55][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][12].cb_test                                      ;
                vDownstreamStackBusLane [55][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][13].cb_test                                      ;
                vDownstreamStackBusLane [55][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][14].cb_test                                      ;
                vDownstreamStackBusLane [55][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][15].cb_test                                      ;
                vDownstreamStackBusLane [55][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][16].cb_test                                      ;
                vDownstreamStackBusLane [55][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][17].cb_test                                      ;
                vDownstreamStackBusLane [55][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][18].cb_test                                      ;
                vDownstreamStackBusLane [55][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][19].cb_test                                      ;
                vDownstreamStackBusLane [55][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][20].cb_test                                      ;
                vDownstreamStackBusLane [55][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][21].cb_test                                      ;
                vDownstreamStackBusLane [55][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][22].cb_test                                      ;
                vDownstreamStackBusLane [55][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][23].cb_test                                      ;
                vDownstreamStackBusLane [55][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][24].cb_test                                      ;
                vDownstreamStackBusLane [55][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][25].cb_test                                      ;
                vDownstreamStackBusLane [55][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][26].cb_test                                      ;
                vDownstreamStackBusLane [55][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][27].cb_test                                      ;
                vDownstreamStackBusLane [55][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][28].cb_test                                      ;
                vDownstreamStackBusLane [55][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][29].cb_test                                      ;
                vDownstreamStackBusLane [55][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][30].cb_test                                      ;
                vDownstreamStackBusLane [55][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[55][31].cb_test                                      ;
                vDownstreamStackBusLane [55][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [55][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[56][0].cb_test                                      ;
                vDownstreamStackBusLane [56][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][1].cb_test                                      ;
                vDownstreamStackBusLane [56][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][2].cb_test                                      ;
                vDownstreamStackBusLane [56][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][3].cb_test                                      ;
                vDownstreamStackBusLane [56][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][4].cb_test                                      ;
                vDownstreamStackBusLane [56][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][5].cb_test                                      ;
                vDownstreamStackBusLane [56][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][6].cb_test                                      ;
                vDownstreamStackBusLane [56][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][7].cb_test                                      ;
                vDownstreamStackBusLane [56][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][8].cb_test                                      ;
                vDownstreamStackBusLane [56][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][9].cb_test                                      ;
                vDownstreamStackBusLane [56][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][10].cb_test                                      ;
                vDownstreamStackBusLane [56][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][11].cb_test                                      ;
                vDownstreamStackBusLane [56][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][12].cb_test                                      ;
                vDownstreamStackBusLane [56][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][13].cb_test                                      ;
                vDownstreamStackBusLane [56][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][14].cb_test                                      ;
                vDownstreamStackBusLane [56][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][15].cb_test                                      ;
                vDownstreamStackBusLane [56][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][16].cb_test                                      ;
                vDownstreamStackBusLane [56][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][17].cb_test                                      ;
                vDownstreamStackBusLane [56][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][18].cb_test                                      ;
                vDownstreamStackBusLane [56][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][19].cb_test                                      ;
                vDownstreamStackBusLane [56][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][20].cb_test                                      ;
                vDownstreamStackBusLane [56][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][21].cb_test                                      ;
                vDownstreamStackBusLane [56][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][22].cb_test                                      ;
                vDownstreamStackBusLane [56][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][23].cb_test                                      ;
                vDownstreamStackBusLane [56][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][24].cb_test                                      ;
                vDownstreamStackBusLane [56][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][25].cb_test                                      ;
                vDownstreamStackBusLane [56][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][26].cb_test                                      ;
                vDownstreamStackBusLane [56][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][27].cb_test                                      ;
                vDownstreamStackBusLane [56][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][28].cb_test                                      ;
                vDownstreamStackBusLane [56][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][29].cb_test                                      ;
                vDownstreamStackBusLane [56][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][30].cb_test                                      ;
                vDownstreamStackBusLane [56][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[56][31].cb_test                                      ;
                vDownstreamStackBusLane [56][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [56][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[57][0].cb_test                                      ;
                vDownstreamStackBusLane [57][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][1].cb_test                                      ;
                vDownstreamStackBusLane [57][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][2].cb_test                                      ;
                vDownstreamStackBusLane [57][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][3].cb_test                                      ;
                vDownstreamStackBusLane [57][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][4].cb_test                                      ;
                vDownstreamStackBusLane [57][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][5].cb_test                                      ;
                vDownstreamStackBusLane [57][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][6].cb_test                                      ;
                vDownstreamStackBusLane [57][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][7].cb_test                                      ;
                vDownstreamStackBusLane [57][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][8].cb_test                                      ;
                vDownstreamStackBusLane [57][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][9].cb_test                                      ;
                vDownstreamStackBusLane [57][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][10].cb_test                                      ;
                vDownstreamStackBusLane [57][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][11].cb_test                                      ;
                vDownstreamStackBusLane [57][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][12].cb_test                                      ;
                vDownstreamStackBusLane [57][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][13].cb_test                                      ;
                vDownstreamStackBusLane [57][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][14].cb_test                                      ;
                vDownstreamStackBusLane [57][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][15].cb_test                                      ;
                vDownstreamStackBusLane [57][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][16].cb_test                                      ;
                vDownstreamStackBusLane [57][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][17].cb_test                                      ;
                vDownstreamStackBusLane [57][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][18].cb_test                                      ;
                vDownstreamStackBusLane [57][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][19].cb_test                                      ;
                vDownstreamStackBusLane [57][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][20].cb_test                                      ;
                vDownstreamStackBusLane [57][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][21].cb_test                                      ;
                vDownstreamStackBusLane [57][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][22].cb_test                                      ;
                vDownstreamStackBusLane [57][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][23].cb_test                                      ;
                vDownstreamStackBusLane [57][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][24].cb_test                                      ;
                vDownstreamStackBusLane [57][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][25].cb_test                                      ;
                vDownstreamStackBusLane [57][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][26].cb_test                                      ;
                vDownstreamStackBusLane [57][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][27].cb_test                                      ;
                vDownstreamStackBusLane [57][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][28].cb_test                                      ;
                vDownstreamStackBusLane [57][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][29].cb_test                                      ;
                vDownstreamStackBusLane [57][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][30].cb_test                                      ;
                vDownstreamStackBusLane [57][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[57][31].cb_test                                      ;
                vDownstreamStackBusLane [57][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [57][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[58][0].cb_test                                      ;
                vDownstreamStackBusLane [58][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][1].cb_test                                      ;
                vDownstreamStackBusLane [58][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][2].cb_test                                      ;
                vDownstreamStackBusLane [58][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][3].cb_test                                      ;
                vDownstreamStackBusLane [58][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][4].cb_test                                      ;
                vDownstreamStackBusLane [58][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][5].cb_test                                      ;
                vDownstreamStackBusLane [58][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][6].cb_test                                      ;
                vDownstreamStackBusLane [58][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][7].cb_test                                      ;
                vDownstreamStackBusLane [58][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][8].cb_test                                      ;
                vDownstreamStackBusLane [58][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][9].cb_test                                      ;
                vDownstreamStackBusLane [58][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][10].cb_test                                      ;
                vDownstreamStackBusLane [58][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][11].cb_test                                      ;
                vDownstreamStackBusLane [58][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][12].cb_test                                      ;
                vDownstreamStackBusLane [58][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][13].cb_test                                      ;
                vDownstreamStackBusLane [58][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][14].cb_test                                      ;
                vDownstreamStackBusLane [58][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][15].cb_test                                      ;
                vDownstreamStackBusLane [58][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][16].cb_test                                      ;
                vDownstreamStackBusLane [58][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][17].cb_test                                      ;
                vDownstreamStackBusLane [58][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][18].cb_test                                      ;
                vDownstreamStackBusLane [58][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][19].cb_test                                      ;
                vDownstreamStackBusLane [58][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][20].cb_test                                      ;
                vDownstreamStackBusLane [58][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][21].cb_test                                      ;
                vDownstreamStackBusLane [58][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][22].cb_test                                      ;
                vDownstreamStackBusLane [58][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][23].cb_test                                      ;
                vDownstreamStackBusLane [58][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][24].cb_test                                      ;
                vDownstreamStackBusLane [58][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][25].cb_test                                      ;
                vDownstreamStackBusLane [58][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][26].cb_test                                      ;
                vDownstreamStackBusLane [58][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][27].cb_test                                      ;
                vDownstreamStackBusLane [58][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][28].cb_test                                      ;
                vDownstreamStackBusLane [58][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][29].cb_test                                      ;
                vDownstreamStackBusLane [58][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][30].cb_test                                      ;
                vDownstreamStackBusLane [58][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[58][31].cb_test                                      ;
                vDownstreamStackBusLane [58][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [58][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[59][0].cb_test                                      ;
                vDownstreamStackBusLane [59][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][1].cb_test                                      ;
                vDownstreamStackBusLane [59][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][2].cb_test                                      ;
                vDownstreamStackBusLane [59][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][3].cb_test                                      ;
                vDownstreamStackBusLane [59][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][4].cb_test                                      ;
                vDownstreamStackBusLane [59][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][5].cb_test                                      ;
                vDownstreamStackBusLane [59][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][6].cb_test                                      ;
                vDownstreamStackBusLane [59][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][7].cb_test                                      ;
                vDownstreamStackBusLane [59][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][8].cb_test                                      ;
                vDownstreamStackBusLane [59][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][9].cb_test                                      ;
                vDownstreamStackBusLane [59][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][10].cb_test                                      ;
                vDownstreamStackBusLane [59][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][11].cb_test                                      ;
                vDownstreamStackBusLane [59][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][12].cb_test                                      ;
                vDownstreamStackBusLane [59][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][13].cb_test                                      ;
                vDownstreamStackBusLane [59][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][14].cb_test                                      ;
                vDownstreamStackBusLane [59][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][15].cb_test                                      ;
                vDownstreamStackBusLane [59][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][16].cb_test                                      ;
                vDownstreamStackBusLane [59][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][17].cb_test                                      ;
                vDownstreamStackBusLane [59][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][18].cb_test                                      ;
                vDownstreamStackBusLane [59][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][19].cb_test                                      ;
                vDownstreamStackBusLane [59][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][20].cb_test                                      ;
                vDownstreamStackBusLane [59][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][21].cb_test                                      ;
                vDownstreamStackBusLane [59][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][22].cb_test                                      ;
                vDownstreamStackBusLane [59][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][23].cb_test                                      ;
                vDownstreamStackBusLane [59][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][24].cb_test                                      ;
                vDownstreamStackBusLane [59][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][25].cb_test                                      ;
                vDownstreamStackBusLane [59][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][26].cb_test                                      ;
                vDownstreamStackBusLane [59][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][27].cb_test                                      ;
                vDownstreamStackBusLane [59][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][28].cb_test                                      ;
                vDownstreamStackBusLane [59][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][29].cb_test                                      ;
                vDownstreamStackBusLane [59][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][30].cb_test                                      ;
                vDownstreamStackBusLane [59][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[59][31].cb_test                                      ;
                vDownstreamStackBusLane [59][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [59][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[60][0].cb_test                                      ;
                vDownstreamStackBusLane [60][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][1].cb_test                                      ;
                vDownstreamStackBusLane [60][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][2].cb_test                                      ;
                vDownstreamStackBusLane [60][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][3].cb_test                                      ;
                vDownstreamStackBusLane [60][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][4].cb_test                                      ;
                vDownstreamStackBusLane [60][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][5].cb_test                                      ;
                vDownstreamStackBusLane [60][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][6].cb_test                                      ;
                vDownstreamStackBusLane [60][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][7].cb_test                                      ;
                vDownstreamStackBusLane [60][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][8].cb_test                                      ;
                vDownstreamStackBusLane [60][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][9].cb_test                                      ;
                vDownstreamStackBusLane [60][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][10].cb_test                                      ;
                vDownstreamStackBusLane [60][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][11].cb_test                                      ;
                vDownstreamStackBusLane [60][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][12].cb_test                                      ;
                vDownstreamStackBusLane [60][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][13].cb_test                                      ;
                vDownstreamStackBusLane [60][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][14].cb_test                                      ;
                vDownstreamStackBusLane [60][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][15].cb_test                                      ;
                vDownstreamStackBusLane [60][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][16].cb_test                                      ;
                vDownstreamStackBusLane [60][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][17].cb_test                                      ;
                vDownstreamStackBusLane [60][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][18].cb_test                                      ;
                vDownstreamStackBusLane [60][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][19].cb_test                                      ;
                vDownstreamStackBusLane [60][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][20].cb_test                                      ;
                vDownstreamStackBusLane [60][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][21].cb_test                                      ;
                vDownstreamStackBusLane [60][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][22].cb_test                                      ;
                vDownstreamStackBusLane [60][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][23].cb_test                                      ;
                vDownstreamStackBusLane [60][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][24].cb_test                                      ;
                vDownstreamStackBusLane [60][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][25].cb_test                                      ;
                vDownstreamStackBusLane [60][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][26].cb_test                                      ;
                vDownstreamStackBusLane [60][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][27].cb_test                                      ;
                vDownstreamStackBusLane [60][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][28].cb_test                                      ;
                vDownstreamStackBusLane [60][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][29].cb_test                                      ;
                vDownstreamStackBusLane [60][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][30].cb_test                                      ;
                vDownstreamStackBusLane [60][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[60][31].cb_test                                      ;
                vDownstreamStackBusLane [60][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [60][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[61][0].cb_test                                      ;
                vDownstreamStackBusLane [61][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][1].cb_test                                      ;
                vDownstreamStackBusLane [61][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][2].cb_test                                      ;
                vDownstreamStackBusLane [61][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][3].cb_test                                      ;
                vDownstreamStackBusLane [61][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][4].cb_test                                      ;
                vDownstreamStackBusLane [61][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][5].cb_test                                      ;
                vDownstreamStackBusLane [61][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][6].cb_test                                      ;
                vDownstreamStackBusLane [61][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][7].cb_test                                      ;
                vDownstreamStackBusLane [61][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][8].cb_test                                      ;
                vDownstreamStackBusLane [61][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][9].cb_test                                      ;
                vDownstreamStackBusLane [61][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][10].cb_test                                      ;
                vDownstreamStackBusLane [61][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][11].cb_test                                      ;
                vDownstreamStackBusLane [61][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][12].cb_test                                      ;
                vDownstreamStackBusLane [61][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][13].cb_test                                      ;
                vDownstreamStackBusLane [61][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][14].cb_test                                      ;
                vDownstreamStackBusLane [61][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][15].cb_test                                      ;
                vDownstreamStackBusLane [61][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][16].cb_test                                      ;
                vDownstreamStackBusLane [61][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][17].cb_test                                      ;
                vDownstreamStackBusLane [61][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][18].cb_test                                      ;
                vDownstreamStackBusLane [61][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][19].cb_test                                      ;
                vDownstreamStackBusLane [61][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][20].cb_test                                      ;
                vDownstreamStackBusLane [61][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][21].cb_test                                      ;
                vDownstreamStackBusLane [61][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][22].cb_test                                      ;
                vDownstreamStackBusLane [61][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][23].cb_test                                      ;
                vDownstreamStackBusLane [61][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][24].cb_test                                      ;
                vDownstreamStackBusLane [61][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][25].cb_test                                      ;
                vDownstreamStackBusLane [61][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][26].cb_test                                      ;
                vDownstreamStackBusLane [61][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][27].cb_test                                      ;
                vDownstreamStackBusLane [61][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][28].cb_test                                      ;
                vDownstreamStackBusLane [61][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][29].cb_test                                      ;
                vDownstreamStackBusLane [61][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][30].cb_test                                      ;
                vDownstreamStackBusLane [61][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[61][31].cb_test                                      ;
                vDownstreamStackBusLane [61][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [61][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[62][0].cb_test                                      ;
                vDownstreamStackBusLane [62][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][1].cb_test                                      ;
                vDownstreamStackBusLane [62][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][2].cb_test                                      ;
                vDownstreamStackBusLane [62][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][3].cb_test                                      ;
                vDownstreamStackBusLane [62][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][4].cb_test                                      ;
                vDownstreamStackBusLane [62][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][5].cb_test                                      ;
                vDownstreamStackBusLane [62][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][6].cb_test                                      ;
                vDownstreamStackBusLane [62][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][7].cb_test                                      ;
                vDownstreamStackBusLane [62][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][8].cb_test                                      ;
                vDownstreamStackBusLane [62][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][9].cb_test                                      ;
                vDownstreamStackBusLane [62][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][10].cb_test                                      ;
                vDownstreamStackBusLane [62][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][11].cb_test                                      ;
                vDownstreamStackBusLane [62][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][12].cb_test                                      ;
                vDownstreamStackBusLane [62][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][13].cb_test                                      ;
                vDownstreamStackBusLane [62][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][14].cb_test                                      ;
                vDownstreamStackBusLane [62][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][15].cb_test                                      ;
                vDownstreamStackBusLane [62][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][16].cb_test                                      ;
                vDownstreamStackBusLane [62][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][17].cb_test                                      ;
                vDownstreamStackBusLane [62][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][18].cb_test                                      ;
                vDownstreamStackBusLane [62][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][19].cb_test                                      ;
                vDownstreamStackBusLane [62][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][20].cb_test                                      ;
                vDownstreamStackBusLane [62][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][21].cb_test                                      ;
                vDownstreamStackBusLane [62][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][22].cb_test                                      ;
                vDownstreamStackBusLane [62][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][23].cb_test                                      ;
                vDownstreamStackBusLane [62][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][24].cb_test                                      ;
                vDownstreamStackBusLane [62][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][25].cb_test                                      ;
                vDownstreamStackBusLane [62][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][26].cb_test                                      ;
                vDownstreamStackBusLane [62][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][27].cb_test                                      ;
                vDownstreamStackBusLane [62][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][28].cb_test                                      ;
                vDownstreamStackBusLane [62][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][29].cb_test                                      ;
                vDownstreamStackBusLane [62][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][30].cb_test                                      ;
                vDownstreamStackBusLane [62][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[62][31].cb_test                                      ;
                vDownstreamStackBusLane [62][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [62][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vDownstreamStackBusLane[63][0].cb_test                                      ;
                vDownstreamStackBusLane [63][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][1].cb_test                                      ;
                vDownstreamStackBusLane [63][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][2].cb_test                                      ;
                vDownstreamStackBusLane [63][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][3].cb_test                                      ;
                vDownstreamStackBusLane [63][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][4].cb_test                                      ;
                vDownstreamStackBusLane [63][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][5].cb_test                                      ;
                vDownstreamStackBusLane [63][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][6].cb_test                                      ;
                vDownstreamStackBusLane [63][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][7].cb_test                                      ;
                vDownstreamStackBusLane [63][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][8].cb_test                                      ;
                vDownstreamStackBusLane [63][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][9].cb_test                                      ;
                vDownstreamStackBusLane [63][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][10].cb_test                                      ;
                vDownstreamStackBusLane [63][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][11].cb_test                                      ;
                vDownstreamStackBusLane [63][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][12].cb_test                                      ;
                vDownstreamStackBusLane [63][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][13].cb_test                                      ;
                vDownstreamStackBusLane [63][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][14].cb_test                                      ;
                vDownstreamStackBusLane [63][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][15].cb_test                                      ;
                vDownstreamStackBusLane [63][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][16].cb_test                                      ;
                vDownstreamStackBusLane [63][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][17].cb_test                                      ;
                vDownstreamStackBusLane [63][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][18].cb_test                                      ;
                vDownstreamStackBusLane [63][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][19].cb_test                                      ;
                vDownstreamStackBusLane [63][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][20].cb_test                                      ;
                vDownstreamStackBusLane [63][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][21].cb_test                                      ;
                vDownstreamStackBusLane [63][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][22].cb_test                                      ;
                vDownstreamStackBusLane [63][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][23].cb_test                                      ;
                vDownstreamStackBusLane [63][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][24].cb_test                                      ;
                vDownstreamStackBusLane [63][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][25].cb_test                                      ;
                vDownstreamStackBusLane [63][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][26].cb_test                                      ;
                vDownstreamStackBusLane [63][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][27].cb_test                                      ;
                vDownstreamStackBusLane [63][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][28].cb_test                                      ;
                vDownstreamStackBusLane [63][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][29].cb_test                                      ;
                vDownstreamStackBusLane [63][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][30].cb_test                                      ;
                vDownstreamStackBusLane [63][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vDownstreamStackBusLane[63][31].cb_test                                      ;
                vDownstreamStackBusLane [63][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vDownstreamStackBusLane [63][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
