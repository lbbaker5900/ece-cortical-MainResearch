

            // ##################################################
            // DMA Stream start addresses

            // Stream 0 start address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [0] = 32'h0010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [1] = 32'h1010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [2] = 32'h2010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [3] = 32'h3010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [4] = 32'h4010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [5] = 32'h5010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [6] = 32'h6010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [7] = 32'h7010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [8] = 32'h8010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [9] = 32'h9010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [10] = 32'ha010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [11] = 32'hb010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [12] = 32'hc010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [13] = 32'hd010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [14] = 32'he010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [15] = 32'hf010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [16] = 32'h10010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [17] = 32'h11010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [18] = 32'h12010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [19] = 32'h13010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [20] = 32'h14010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [21] = 32'h15010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [22] = 32'h16010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [23] = 32'h17010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [24] = 32'h18010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [25] = 32'h19010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [26] = 32'h1a010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [27] = 32'h1b010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [28] = 32'h1c010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [29] = 32'h1d010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [30] = 32'h1e010;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r134 [31] = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [0] = 32'h0800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [1] = 32'h1800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [2] = 32'h2800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [3] = 32'h3800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [4] = 32'h4800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [5] = 32'h5800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [6] = 32'h6800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [7] = 32'h7800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [8] = 32'h8800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [9] = 32'h9800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [10] = 32'ha800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [11] = 32'hb800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [12] = 32'hc800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [13] = 32'hd800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [14] = 32'he800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [15] = 32'hf800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [16] = 32'h10800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [17] = 32'h11800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [18] = 32'h12800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [19] = 32'h13800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [20] = 32'h14800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [21] = 32'h15800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [22] = 32'h16800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [23] = 32'h17800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [24] = 32'h18800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [25] = 32'h19800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [26] = 32'h1a800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [27] = 32'h1b800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [28] = 32'h1c800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [29] = 32'h1d800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [30] = 32'h1e800;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r135 [31] = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [0] = 32'h0010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [1] = 32'h1010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [2] = 32'h2010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [3] = 32'h3010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [4] = 32'h4010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [5] = 32'h5010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [6] = 32'h6010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [7] = 32'h7010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [8] = 32'h8010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [9] = 32'h9010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [10] = 32'ha010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [11] = 32'hb010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [12] = 32'hc010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [13] = 32'hd010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [14] = 32'he010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [15] = 32'hf010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [16] = 32'h10010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [17] = 32'h11010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [18] = 32'h12010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [19] = 32'h13010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [20] = 32'h14010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [21] = 32'h15010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [22] = 32'h16010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [23] = 32'h17010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [24] = 32'h18010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [25] = 32'h19010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [26] = 32'h1a010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [27] = 32'h1b010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [28] = 32'h1c010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [29] = 32'h1d010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [30] = 32'h1e010;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r134 [31] = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [0] = 32'h0800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [1] = 32'h1800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [2] = 32'h2800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [3] = 32'h3800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [4] = 32'h4800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [5] = 32'h5800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [6] = 32'h6800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [7] = 32'h7800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [8] = 32'h8800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [9] = 32'h9800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [10] = 32'ha800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [11] = 32'hb800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [12] = 32'hc800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [13] = 32'hd800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [14] = 32'he800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [15] = 32'hf800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [16] = 32'h10800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [17] = 32'h11800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [18] = 32'h12800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [19] = 32'h13800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [20] = 32'h14800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [21] = 32'h15800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [22] = 32'h16800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [23] = 32'h17800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [24] = 32'h18800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [25] = 32'h19800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [26] = 32'h1a800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [27] = 32'h1b800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [28] = 32'h1c800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [29] = 32'h1d800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [30] = 32'h1e800;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r135 [31] = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [0] = 32'h0010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [1] = 32'h1010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [2] = 32'h2010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [3] = 32'h3010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [4] = 32'h4010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [5] = 32'h5010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [6] = 32'h6010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [7] = 32'h7010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [8] = 32'h8010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [9] = 32'h9010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [10] = 32'ha010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [11] = 32'hb010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [12] = 32'hc010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [13] = 32'hd010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [14] = 32'he010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [15] = 32'hf010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [16] = 32'h10010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [17] = 32'h11010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [18] = 32'h12010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [19] = 32'h13010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [20] = 32'h14010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [21] = 32'h15010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [22] = 32'h16010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [23] = 32'h17010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [24] = 32'h18010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [25] = 32'h19010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [26] = 32'h1a010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [27] = 32'h1b010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [28] = 32'h1c010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [29] = 32'h1d010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [30] = 32'h1e010;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r134 [31] = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [0] = 32'h0800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [1] = 32'h1800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [2] = 32'h2800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [3] = 32'h3800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [4] = 32'h4800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [5] = 32'h5800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [6] = 32'h6800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [7] = 32'h7800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [8] = 32'h8800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [9] = 32'h9800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [10] = 32'ha800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [11] = 32'hb800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [12] = 32'hc800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [13] = 32'hd800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [14] = 32'he800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [15] = 32'hf800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [16] = 32'h10800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [17] = 32'h11800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [18] = 32'h12800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [19] = 32'h13800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [20] = 32'h14800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [21] = 32'h15800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [22] = 32'h16800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [23] = 32'h17800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [24] = 32'h18800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [25] = 32'h19800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [26] = 32'h1a800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [27] = 32'h1b800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [28] = 32'h1c800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [29] = 32'h1d800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [30] = 32'h1e800;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r135 [31] = 32'h1f800;
            // Stream 0 start address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [0] = 32'h0010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [1] = 32'h1010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [2] = 32'h2010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [3] = 32'h3010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [4] = 32'h4010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [5] = 32'h5010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [6] = 32'h6010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [7] = 32'h7010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [8] = 32'h8010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [9] = 32'h9010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [10] = 32'ha010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [11] = 32'hb010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [12] = 32'hc010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [13] = 32'hd010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [14] = 32'he010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [15] = 32'hf010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [16] = 32'h10010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [17] = 32'h11010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [18] = 32'h12010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [19] = 32'h13010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [20] = 32'h14010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [21] = 32'h15010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [22] = 32'h16010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [23] = 32'h17010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [24] = 32'h18010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [25] = 32'h19010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [26] = 32'h1a010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [27] = 32'h1b010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [28] = 32'h1c010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [29] = 32'h1d010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [30] = 32'h1e010;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r134 [31] = 32'h1f010;
            // Stream 1 start address
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [0] = 32'h0800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [1] = 32'h1800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [2] = 32'h2800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [3] = 32'h3800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [4] = 32'h4800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [5] = 32'h5800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [6] = 32'h6800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [7] = 32'h7800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [8] = 32'h8800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [9] = 32'h9800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [10] = 32'ha800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [11] = 32'hb800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [12] = 32'hc800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [13] = 32'hd800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [14] = 32'he800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [15] = 32'hf800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [16] = 32'h10800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [17] = 32'h11800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [18] = 32'h12800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [19] = 32'h13800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [20] = 32'h14800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [21] = 32'h15800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [22] = 32'h16800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [23] = 32'h17800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [24] = 32'h18800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [25] = 32'h19800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [26] = 32'h1a800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [27] = 32'h1b800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [28] = 32'h1c800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [29] = 32'h1d800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [30] = 32'h1e800;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r135 [31] = 32'h1f800;

            // ##################################################
            // DMA Type and length of stream

            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r132[31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[0].pe.simd__scntl__lane_r133[31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r132[31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__lane_r133[31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r132[31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__lane_r133[31][15:0]  = numOfTypes;
            // Set data type and size of stream0 (in types)
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r132[31][15:0]  = numOfTypes;
            // Set data type and size of stream1 (in types)
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[0][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[0][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[1][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[1][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[2][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[2][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[3][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[3][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[4][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[4][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[5][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[5][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[6][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[6][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[7][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[7][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[8][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[8][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[9][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[9][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[10][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[10][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[11][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[11][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[12][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[12][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[13][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[13][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[14][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[14][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[15][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[15][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[16][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[16][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[17][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[17][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[18][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[18][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[19][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[19][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[20][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[20][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[21][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[21][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[22][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[22][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[23][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[23][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[24][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[24][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[25][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[25][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[26][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[26][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[27][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[27][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[28][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[28][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[29][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[29][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[30][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[30][15:0]  = numOfTypes;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[31][19:16] = 4'd4;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__lane_r133[31][15:0]  = numOfTypes;

            // ##################################################
            // Enable and set transfer type

            repeat(10) @(negedge clk); 

            // Enable
            force pe_array_inst.pe_inst[0].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__rs0[0]           = 1'b1;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__rs0[0]           = 1'b1;

            // Operation
            force pe_array_inst.pe_inst[0].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[1].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[2].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;
            force pe_array_inst.pe_inst[3].pe.simd__scntl__rs0[31:1] = `STREAMING_OP_CNTL_OPERATION_NOP_FROM_TWO_EXT_TO_MEM ;

            repeat(50) @(negedge clk);