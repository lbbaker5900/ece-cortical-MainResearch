
  assign   pe_inst[0].sys__pe__allSynchronized    =  sys__pe0__allSynchronized                ;
  assign   pe0__sys__thisSynchronized             =  pe_inst[0].pe__sys__thisSynchronized     ;
  assign   pe0__sys__ready                        =  pe_inst[0].pe__sys__ready                ;
  assign   pe0__sys__complete                     =  pe_inst[0].pe__sys__complete             ;
  assign   pe_inst[0].std__pe__oob_cntl           =  std__pe0__oob_cntl                       ;
  assign   pe_inst[0].std__pe__oob_valid          =  std__pe0__oob_valid                      ;
  assign   pe0__std__oob_ready                    =  pe_inst[0].pe__std__oob_ready            ;
  assign   pe_inst[0].std__pe__oob_type           =  std__pe0__oob_type                       ;
  assign   pe_inst[0].std__pe__oob_data           =  std__pe0__oob_data                       ;
  assign   pe_inst[1].sys__pe__allSynchronized    =  sys__pe1__allSynchronized                ;
  assign   pe1__sys__thisSynchronized             =  pe_inst[1].pe__sys__thisSynchronized     ;
  assign   pe1__sys__ready                        =  pe_inst[1].pe__sys__ready                ;
  assign   pe1__sys__complete                     =  pe_inst[1].pe__sys__complete             ;
  assign   pe_inst[1].std__pe__oob_cntl           =  std__pe1__oob_cntl                       ;
  assign   pe_inst[1].std__pe__oob_valid          =  std__pe1__oob_valid                      ;
  assign   pe1__std__oob_ready                    =  pe_inst[1].pe__std__oob_ready            ;
  assign   pe_inst[1].std__pe__oob_type           =  std__pe1__oob_type                       ;
  assign   pe_inst[1].std__pe__oob_data           =  std__pe1__oob_data                       ;
  assign   pe_inst[2].sys__pe__allSynchronized    =  sys__pe2__allSynchronized                ;
  assign   pe2__sys__thisSynchronized             =  pe_inst[2].pe__sys__thisSynchronized     ;
  assign   pe2__sys__ready                        =  pe_inst[2].pe__sys__ready                ;
  assign   pe2__sys__complete                     =  pe_inst[2].pe__sys__complete             ;
  assign   pe_inst[2].std__pe__oob_cntl           =  std__pe2__oob_cntl                       ;
  assign   pe_inst[2].std__pe__oob_valid          =  std__pe2__oob_valid                      ;
  assign   pe2__std__oob_ready                    =  pe_inst[2].pe__std__oob_ready            ;
  assign   pe_inst[2].std__pe__oob_type           =  std__pe2__oob_type                       ;
  assign   pe_inst[2].std__pe__oob_data           =  std__pe2__oob_data                       ;
  assign   pe_inst[3].sys__pe__allSynchronized    =  sys__pe3__allSynchronized                ;
  assign   pe3__sys__thisSynchronized             =  pe_inst[3].pe__sys__thisSynchronized     ;
  assign   pe3__sys__ready                        =  pe_inst[3].pe__sys__ready                ;
  assign   pe3__sys__complete                     =  pe_inst[3].pe__sys__complete             ;
  assign   pe_inst[3].std__pe__oob_cntl           =  std__pe3__oob_cntl                       ;
  assign   pe_inst[3].std__pe__oob_valid          =  std__pe3__oob_valid                      ;
  assign   pe3__std__oob_ready                    =  pe_inst[3].pe__std__oob_ready            ;
  assign   pe_inst[3].std__pe__oob_type           =  std__pe3__oob_type                       ;
  assign   pe_inst[3].std__pe__oob_data           =  std__pe3__oob_data                       ;
  assign   pe_inst[4].sys__pe__allSynchronized    =  sys__pe4__allSynchronized                ;
  assign   pe4__sys__thisSynchronized             =  pe_inst[4].pe__sys__thisSynchronized     ;
  assign   pe4__sys__ready                        =  pe_inst[4].pe__sys__ready                ;
  assign   pe4__sys__complete                     =  pe_inst[4].pe__sys__complete             ;
  assign   pe_inst[4].std__pe__oob_cntl           =  std__pe4__oob_cntl                       ;
  assign   pe_inst[4].std__pe__oob_valid          =  std__pe4__oob_valid                      ;
  assign   pe4__std__oob_ready                    =  pe_inst[4].pe__std__oob_ready            ;
  assign   pe_inst[4].std__pe__oob_type           =  std__pe4__oob_type                       ;
  assign   pe_inst[4].std__pe__oob_data           =  std__pe4__oob_data                       ;
  assign   pe_inst[5].sys__pe__allSynchronized    =  sys__pe5__allSynchronized                ;
  assign   pe5__sys__thisSynchronized             =  pe_inst[5].pe__sys__thisSynchronized     ;
  assign   pe5__sys__ready                        =  pe_inst[5].pe__sys__ready                ;
  assign   pe5__sys__complete                     =  pe_inst[5].pe__sys__complete             ;
  assign   pe_inst[5].std__pe__oob_cntl           =  std__pe5__oob_cntl                       ;
  assign   pe_inst[5].std__pe__oob_valid          =  std__pe5__oob_valid                      ;
  assign   pe5__std__oob_ready                    =  pe_inst[5].pe__std__oob_ready            ;
  assign   pe_inst[5].std__pe__oob_type           =  std__pe5__oob_type                       ;
  assign   pe_inst[5].std__pe__oob_data           =  std__pe5__oob_data                       ;
  assign   pe_inst[6].sys__pe__allSynchronized    =  sys__pe6__allSynchronized                ;
  assign   pe6__sys__thisSynchronized             =  pe_inst[6].pe__sys__thisSynchronized     ;
  assign   pe6__sys__ready                        =  pe_inst[6].pe__sys__ready                ;
  assign   pe6__sys__complete                     =  pe_inst[6].pe__sys__complete             ;
  assign   pe_inst[6].std__pe__oob_cntl           =  std__pe6__oob_cntl                       ;
  assign   pe_inst[6].std__pe__oob_valid          =  std__pe6__oob_valid                      ;
  assign   pe6__std__oob_ready                    =  pe_inst[6].pe__std__oob_ready            ;
  assign   pe_inst[6].std__pe__oob_type           =  std__pe6__oob_type                       ;
  assign   pe_inst[6].std__pe__oob_data           =  std__pe6__oob_data                       ;
  assign   pe_inst[7].sys__pe__allSynchronized    =  sys__pe7__allSynchronized                ;
  assign   pe7__sys__thisSynchronized             =  pe_inst[7].pe__sys__thisSynchronized     ;
  assign   pe7__sys__ready                        =  pe_inst[7].pe__sys__ready                ;
  assign   pe7__sys__complete                     =  pe_inst[7].pe__sys__complete             ;
  assign   pe_inst[7].std__pe__oob_cntl           =  std__pe7__oob_cntl                       ;
  assign   pe_inst[7].std__pe__oob_valid          =  std__pe7__oob_valid                      ;
  assign   pe7__std__oob_ready                    =  pe_inst[7].pe__std__oob_ready            ;
  assign   pe_inst[7].std__pe__oob_type           =  std__pe7__oob_type                       ;
  assign   pe_inst[7].std__pe__oob_data           =  std__pe7__oob_data                       ;
  assign   pe_inst[8].sys__pe__allSynchronized    =  sys__pe8__allSynchronized                ;
  assign   pe8__sys__thisSynchronized             =  pe_inst[8].pe__sys__thisSynchronized     ;
  assign   pe8__sys__ready                        =  pe_inst[8].pe__sys__ready                ;
  assign   pe8__sys__complete                     =  pe_inst[8].pe__sys__complete             ;
  assign   pe_inst[8].std__pe__oob_cntl           =  std__pe8__oob_cntl                       ;
  assign   pe_inst[8].std__pe__oob_valid          =  std__pe8__oob_valid                      ;
  assign   pe8__std__oob_ready                    =  pe_inst[8].pe__std__oob_ready            ;
  assign   pe_inst[8].std__pe__oob_type           =  std__pe8__oob_type                       ;
  assign   pe_inst[8].std__pe__oob_data           =  std__pe8__oob_data                       ;
  assign   pe_inst[9].sys__pe__allSynchronized    =  sys__pe9__allSynchronized                ;
  assign   pe9__sys__thisSynchronized             =  pe_inst[9].pe__sys__thisSynchronized     ;
  assign   pe9__sys__ready                        =  pe_inst[9].pe__sys__ready                ;
  assign   pe9__sys__complete                     =  pe_inst[9].pe__sys__complete             ;
  assign   pe_inst[9].std__pe__oob_cntl           =  std__pe9__oob_cntl                       ;
  assign   pe_inst[9].std__pe__oob_valid          =  std__pe9__oob_valid                      ;
  assign   pe9__std__oob_ready                    =  pe_inst[9].pe__std__oob_ready            ;
  assign   pe_inst[9].std__pe__oob_type           =  std__pe9__oob_type                       ;
  assign   pe_inst[9].std__pe__oob_data           =  std__pe9__oob_data                       ;
  assign   pe_inst[10].sys__pe__allSynchronized    =  sys__pe10__allSynchronized                ;
  assign   pe10__sys__thisSynchronized             =  pe_inst[10].pe__sys__thisSynchronized     ;
  assign   pe10__sys__ready                        =  pe_inst[10].pe__sys__ready                ;
  assign   pe10__sys__complete                     =  pe_inst[10].pe__sys__complete             ;
  assign   pe_inst[10].std__pe__oob_cntl           =  std__pe10__oob_cntl                       ;
  assign   pe_inst[10].std__pe__oob_valid          =  std__pe10__oob_valid                      ;
  assign   pe10__std__oob_ready                    =  pe_inst[10].pe__std__oob_ready            ;
  assign   pe_inst[10].std__pe__oob_type           =  std__pe10__oob_type                       ;
  assign   pe_inst[10].std__pe__oob_data           =  std__pe10__oob_data                       ;
  assign   pe_inst[11].sys__pe__allSynchronized    =  sys__pe11__allSynchronized                ;
  assign   pe11__sys__thisSynchronized             =  pe_inst[11].pe__sys__thisSynchronized     ;
  assign   pe11__sys__ready                        =  pe_inst[11].pe__sys__ready                ;
  assign   pe11__sys__complete                     =  pe_inst[11].pe__sys__complete             ;
  assign   pe_inst[11].std__pe__oob_cntl           =  std__pe11__oob_cntl                       ;
  assign   pe_inst[11].std__pe__oob_valid          =  std__pe11__oob_valid                      ;
  assign   pe11__std__oob_ready                    =  pe_inst[11].pe__std__oob_ready            ;
  assign   pe_inst[11].std__pe__oob_type           =  std__pe11__oob_type                       ;
  assign   pe_inst[11].std__pe__oob_data           =  std__pe11__oob_data                       ;
  assign   pe_inst[12].sys__pe__allSynchronized    =  sys__pe12__allSynchronized                ;
  assign   pe12__sys__thisSynchronized             =  pe_inst[12].pe__sys__thisSynchronized     ;
  assign   pe12__sys__ready                        =  pe_inst[12].pe__sys__ready                ;
  assign   pe12__sys__complete                     =  pe_inst[12].pe__sys__complete             ;
  assign   pe_inst[12].std__pe__oob_cntl           =  std__pe12__oob_cntl                       ;
  assign   pe_inst[12].std__pe__oob_valid          =  std__pe12__oob_valid                      ;
  assign   pe12__std__oob_ready                    =  pe_inst[12].pe__std__oob_ready            ;
  assign   pe_inst[12].std__pe__oob_type           =  std__pe12__oob_type                       ;
  assign   pe_inst[12].std__pe__oob_data           =  std__pe12__oob_data                       ;
  assign   pe_inst[13].sys__pe__allSynchronized    =  sys__pe13__allSynchronized                ;
  assign   pe13__sys__thisSynchronized             =  pe_inst[13].pe__sys__thisSynchronized     ;
  assign   pe13__sys__ready                        =  pe_inst[13].pe__sys__ready                ;
  assign   pe13__sys__complete                     =  pe_inst[13].pe__sys__complete             ;
  assign   pe_inst[13].std__pe__oob_cntl           =  std__pe13__oob_cntl                       ;
  assign   pe_inst[13].std__pe__oob_valid          =  std__pe13__oob_valid                      ;
  assign   pe13__std__oob_ready                    =  pe_inst[13].pe__std__oob_ready            ;
  assign   pe_inst[13].std__pe__oob_type           =  std__pe13__oob_type                       ;
  assign   pe_inst[13].std__pe__oob_data           =  std__pe13__oob_data                       ;
  assign   pe_inst[14].sys__pe__allSynchronized    =  sys__pe14__allSynchronized                ;
  assign   pe14__sys__thisSynchronized             =  pe_inst[14].pe__sys__thisSynchronized     ;
  assign   pe14__sys__ready                        =  pe_inst[14].pe__sys__ready                ;
  assign   pe14__sys__complete                     =  pe_inst[14].pe__sys__complete             ;
  assign   pe_inst[14].std__pe__oob_cntl           =  std__pe14__oob_cntl                       ;
  assign   pe_inst[14].std__pe__oob_valid          =  std__pe14__oob_valid                      ;
  assign   pe14__std__oob_ready                    =  pe_inst[14].pe__std__oob_ready            ;
  assign   pe_inst[14].std__pe__oob_type           =  std__pe14__oob_type                       ;
  assign   pe_inst[14].std__pe__oob_data           =  std__pe14__oob_data                       ;
  assign   pe_inst[15].sys__pe__allSynchronized    =  sys__pe15__allSynchronized                ;
  assign   pe15__sys__thisSynchronized             =  pe_inst[15].pe__sys__thisSynchronized     ;
  assign   pe15__sys__ready                        =  pe_inst[15].pe__sys__ready                ;
  assign   pe15__sys__complete                     =  pe_inst[15].pe__sys__complete             ;
  assign   pe_inst[15].std__pe__oob_cntl           =  std__pe15__oob_cntl                       ;
  assign   pe_inst[15].std__pe__oob_valid          =  std__pe15__oob_valid                      ;
  assign   pe15__std__oob_ready                    =  pe_inst[15].pe__std__oob_ready            ;
  assign   pe_inst[15].std__pe__oob_type           =  std__pe15__oob_type                       ;
  assign   pe_inst[15].std__pe__oob_data           =  std__pe15__oob_data                       ;
  assign   pe_inst[16].sys__pe__allSynchronized    =  sys__pe16__allSynchronized                ;
  assign   pe16__sys__thisSynchronized             =  pe_inst[16].pe__sys__thisSynchronized     ;
  assign   pe16__sys__ready                        =  pe_inst[16].pe__sys__ready                ;
  assign   pe16__sys__complete                     =  pe_inst[16].pe__sys__complete             ;
  assign   pe_inst[16].std__pe__oob_cntl           =  std__pe16__oob_cntl                       ;
  assign   pe_inst[16].std__pe__oob_valid          =  std__pe16__oob_valid                      ;
  assign   pe16__std__oob_ready                    =  pe_inst[16].pe__std__oob_ready            ;
  assign   pe_inst[16].std__pe__oob_type           =  std__pe16__oob_type                       ;
  assign   pe_inst[16].std__pe__oob_data           =  std__pe16__oob_data                       ;
  assign   pe_inst[17].sys__pe__allSynchronized    =  sys__pe17__allSynchronized                ;
  assign   pe17__sys__thisSynchronized             =  pe_inst[17].pe__sys__thisSynchronized     ;
  assign   pe17__sys__ready                        =  pe_inst[17].pe__sys__ready                ;
  assign   pe17__sys__complete                     =  pe_inst[17].pe__sys__complete             ;
  assign   pe_inst[17].std__pe__oob_cntl           =  std__pe17__oob_cntl                       ;
  assign   pe_inst[17].std__pe__oob_valid          =  std__pe17__oob_valid                      ;
  assign   pe17__std__oob_ready                    =  pe_inst[17].pe__std__oob_ready            ;
  assign   pe_inst[17].std__pe__oob_type           =  std__pe17__oob_type                       ;
  assign   pe_inst[17].std__pe__oob_data           =  std__pe17__oob_data                       ;
  assign   pe_inst[18].sys__pe__allSynchronized    =  sys__pe18__allSynchronized                ;
  assign   pe18__sys__thisSynchronized             =  pe_inst[18].pe__sys__thisSynchronized     ;
  assign   pe18__sys__ready                        =  pe_inst[18].pe__sys__ready                ;
  assign   pe18__sys__complete                     =  pe_inst[18].pe__sys__complete             ;
  assign   pe_inst[18].std__pe__oob_cntl           =  std__pe18__oob_cntl                       ;
  assign   pe_inst[18].std__pe__oob_valid          =  std__pe18__oob_valid                      ;
  assign   pe18__std__oob_ready                    =  pe_inst[18].pe__std__oob_ready            ;
  assign   pe_inst[18].std__pe__oob_type           =  std__pe18__oob_type                       ;
  assign   pe_inst[18].std__pe__oob_data           =  std__pe18__oob_data                       ;
  assign   pe_inst[19].sys__pe__allSynchronized    =  sys__pe19__allSynchronized                ;
  assign   pe19__sys__thisSynchronized             =  pe_inst[19].pe__sys__thisSynchronized     ;
  assign   pe19__sys__ready                        =  pe_inst[19].pe__sys__ready                ;
  assign   pe19__sys__complete                     =  pe_inst[19].pe__sys__complete             ;
  assign   pe_inst[19].std__pe__oob_cntl           =  std__pe19__oob_cntl                       ;
  assign   pe_inst[19].std__pe__oob_valid          =  std__pe19__oob_valid                      ;
  assign   pe19__std__oob_ready                    =  pe_inst[19].pe__std__oob_ready            ;
  assign   pe_inst[19].std__pe__oob_type           =  std__pe19__oob_type                       ;
  assign   pe_inst[19].std__pe__oob_data           =  std__pe19__oob_data                       ;
  assign   pe_inst[20].sys__pe__allSynchronized    =  sys__pe20__allSynchronized                ;
  assign   pe20__sys__thisSynchronized             =  pe_inst[20].pe__sys__thisSynchronized     ;
  assign   pe20__sys__ready                        =  pe_inst[20].pe__sys__ready                ;
  assign   pe20__sys__complete                     =  pe_inst[20].pe__sys__complete             ;
  assign   pe_inst[20].std__pe__oob_cntl           =  std__pe20__oob_cntl                       ;
  assign   pe_inst[20].std__pe__oob_valid          =  std__pe20__oob_valid                      ;
  assign   pe20__std__oob_ready                    =  pe_inst[20].pe__std__oob_ready            ;
  assign   pe_inst[20].std__pe__oob_type           =  std__pe20__oob_type                       ;
  assign   pe_inst[20].std__pe__oob_data           =  std__pe20__oob_data                       ;
  assign   pe_inst[21].sys__pe__allSynchronized    =  sys__pe21__allSynchronized                ;
  assign   pe21__sys__thisSynchronized             =  pe_inst[21].pe__sys__thisSynchronized     ;
  assign   pe21__sys__ready                        =  pe_inst[21].pe__sys__ready                ;
  assign   pe21__sys__complete                     =  pe_inst[21].pe__sys__complete             ;
  assign   pe_inst[21].std__pe__oob_cntl           =  std__pe21__oob_cntl                       ;
  assign   pe_inst[21].std__pe__oob_valid          =  std__pe21__oob_valid                      ;
  assign   pe21__std__oob_ready                    =  pe_inst[21].pe__std__oob_ready            ;
  assign   pe_inst[21].std__pe__oob_type           =  std__pe21__oob_type                       ;
  assign   pe_inst[21].std__pe__oob_data           =  std__pe21__oob_data                       ;
  assign   pe_inst[22].sys__pe__allSynchronized    =  sys__pe22__allSynchronized                ;
  assign   pe22__sys__thisSynchronized             =  pe_inst[22].pe__sys__thisSynchronized     ;
  assign   pe22__sys__ready                        =  pe_inst[22].pe__sys__ready                ;
  assign   pe22__sys__complete                     =  pe_inst[22].pe__sys__complete             ;
  assign   pe_inst[22].std__pe__oob_cntl           =  std__pe22__oob_cntl                       ;
  assign   pe_inst[22].std__pe__oob_valid          =  std__pe22__oob_valid                      ;
  assign   pe22__std__oob_ready                    =  pe_inst[22].pe__std__oob_ready            ;
  assign   pe_inst[22].std__pe__oob_type           =  std__pe22__oob_type                       ;
  assign   pe_inst[22].std__pe__oob_data           =  std__pe22__oob_data                       ;
  assign   pe_inst[23].sys__pe__allSynchronized    =  sys__pe23__allSynchronized                ;
  assign   pe23__sys__thisSynchronized             =  pe_inst[23].pe__sys__thisSynchronized     ;
  assign   pe23__sys__ready                        =  pe_inst[23].pe__sys__ready                ;
  assign   pe23__sys__complete                     =  pe_inst[23].pe__sys__complete             ;
  assign   pe_inst[23].std__pe__oob_cntl           =  std__pe23__oob_cntl                       ;
  assign   pe_inst[23].std__pe__oob_valid          =  std__pe23__oob_valid                      ;
  assign   pe23__std__oob_ready                    =  pe_inst[23].pe__std__oob_ready            ;
  assign   pe_inst[23].std__pe__oob_type           =  std__pe23__oob_type                       ;
  assign   pe_inst[23].std__pe__oob_data           =  std__pe23__oob_data                       ;
  assign   pe_inst[24].sys__pe__allSynchronized    =  sys__pe24__allSynchronized                ;
  assign   pe24__sys__thisSynchronized             =  pe_inst[24].pe__sys__thisSynchronized     ;
  assign   pe24__sys__ready                        =  pe_inst[24].pe__sys__ready                ;
  assign   pe24__sys__complete                     =  pe_inst[24].pe__sys__complete             ;
  assign   pe_inst[24].std__pe__oob_cntl           =  std__pe24__oob_cntl                       ;
  assign   pe_inst[24].std__pe__oob_valid          =  std__pe24__oob_valid                      ;
  assign   pe24__std__oob_ready                    =  pe_inst[24].pe__std__oob_ready            ;
  assign   pe_inst[24].std__pe__oob_type           =  std__pe24__oob_type                       ;
  assign   pe_inst[24].std__pe__oob_data           =  std__pe24__oob_data                       ;
  assign   pe_inst[25].sys__pe__allSynchronized    =  sys__pe25__allSynchronized                ;
  assign   pe25__sys__thisSynchronized             =  pe_inst[25].pe__sys__thisSynchronized     ;
  assign   pe25__sys__ready                        =  pe_inst[25].pe__sys__ready                ;
  assign   pe25__sys__complete                     =  pe_inst[25].pe__sys__complete             ;
  assign   pe_inst[25].std__pe__oob_cntl           =  std__pe25__oob_cntl                       ;
  assign   pe_inst[25].std__pe__oob_valid          =  std__pe25__oob_valid                      ;
  assign   pe25__std__oob_ready                    =  pe_inst[25].pe__std__oob_ready            ;
  assign   pe_inst[25].std__pe__oob_type           =  std__pe25__oob_type                       ;
  assign   pe_inst[25].std__pe__oob_data           =  std__pe25__oob_data                       ;
  assign   pe_inst[26].sys__pe__allSynchronized    =  sys__pe26__allSynchronized                ;
  assign   pe26__sys__thisSynchronized             =  pe_inst[26].pe__sys__thisSynchronized     ;
  assign   pe26__sys__ready                        =  pe_inst[26].pe__sys__ready                ;
  assign   pe26__sys__complete                     =  pe_inst[26].pe__sys__complete             ;
  assign   pe_inst[26].std__pe__oob_cntl           =  std__pe26__oob_cntl                       ;
  assign   pe_inst[26].std__pe__oob_valid          =  std__pe26__oob_valid                      ;
  assign   pe26__std__oob_ready                    =  pe_inst[26].pe__std__oob_ready            ;
  assign   pe_inst[26].std__pe__oob_type           =  std__pe26__oob_type                       ;
  assign   pe_inst[26].std__pe__oob_data           =  std__pe26__oob_data                       ;
  assign   pe_inst[27].sys__pe__allSynchronized    =  sys__pe27__allSynchronized                ;
  assign   pe27__sys__thisSynchronized             =  pe_inst[27].pe__sys__thisSynchronized     ;
  assign   pe27__sys__ready                        =  pe_inst[27].pe__sys__ready                ;
  assign   pe27__sys__complete                     =  pe_inst[27].pe__sys__complete             ;
  assign   pe_inst[27].std__pe__oob_cntl           =  std__pe27__oob_cntl                       ;
  assign   pe_inst[27].std__pe__oob_valid          =  std__pe27__oob_valid                      ;
  assign   pe27__std__oob_ready                    =  pe_inst[27].pe__std__oob_ready            ;
  assign   pe_inst[27].std__pe__oob_type           =  std__pe27__oob_type                       ;
  assign   pe_inst[27].std__pe__oob_data           =  std__pe27__oob_data                       ;
  assign   pe_inst[28].sys__pe__allSynchronized    =  sys__pe28__allSynchronized                ;
  assign   pe28__sys__thisSynchronized             =  pe_inst[28].pe__sys__thisSynchronized     ;
  assign   pe28__sys__ready                        =  pe_inst[28].pe__sys__ready                ;
  assign   pe28__sys__complete                     =  pe_inst[28].pe__sys__complete             ;
  assign   pe_inst[28].std__pe__oob_cntl           =  std__pe28__oob_cntl                       ;
  assign   pe_inst[28].std__pe__oob_valid          =  std__pe28__oob_valid                      ;
  assign   pe28__std__oob_ready                    =  pe_inst[28].pe__std__oob_ready            ;
  assign   pe_inst[28].std__pe__oob_type           =  std__pe28__oob_type                       ;
  assign   pe_inst[28].std__pe__oob_data           =  std__pe28__oob_data                       ;
  assign   pe_inst[29].sys__pe__allSynchronized    =  sys__pe29__allSynchronized                ;
  assign   pe29__sys__thisSynchronized             =  pe_inst[29].pe__sys__thisSynchronized     ;
  assign   pe29__sys__ready                        =  pe_inst[29].pe__sys__ready                ;
  assign   pe29__sys__complete                     =  pe_inst[29].pe__sys__complete             ;
  assign   pe_inst[29].std__pe__oob_cntl           =  std__pe29__oob_cntl                       ;
  assign   pe_inst[29].std__pe__oob_valid          =  std__pe29__oob_valid                      ;
  assign   pe29__std__oob_ready                    =  pe_inst[29].pe__std__oob_ready            ;
  assign   pe_inst[29].std__pe__oob_type           =  std__pe29__oob_type                       ;
  assign   pe_inst[29].std__pe__oob_data           =  std__pe29__oob_data                       ;
  assign   pe_inst[30].sys__pe__allSynchronized    =  sys__pe30__allSynchronized                ;
  assign   pe30__sys__thisSynchronized             =  pe_inst[30].pe__sys__thisSynchronized     ;
  assign   pe30__sys__ready                        =  pe_inst[30].pe__sys__ready                ;
  assign   pe30__sys__complete                     =  pe_inst[30].pe__sys__complete             ;
  assign   pe_inst[30].std__pe__oob_cntl           =  std__pe30__oob_cntl                       ;
  assign   pe_inst[30].std__pe__oob_valid          =  std__pe30__oob_valid                      ;
  assign   pe30__std__oob_ready                    =  pe_inst[30].pe__std__oob_ready            ;
  assign   pe_inst[30].std__pe__oob_type           =  std__pe30__oob_type                       ;
  assign   pe_inst[30].std__pe__oob_data           =  std__pe30__oob_data                       ;
  assign   pe_inst[31].sys__pe__allSynchronized    =  sys__pe31__allSynchronized                ;
  assign   pe31__sys__thisSynchronized             =  pe_inst[31].pe__sys__thisSynchronized     ;
  assign   pe31__sys__ready                        =  pe_inst[31].pe__sys__ready                ;
  assign   pe31__sys__complete                     =  pe_inst[31].pe__sys__complete             ;
  assign   pe_inst[31].std__pe__oob_cntl           =  std__pe31__oob_cntl                       ;
  assign   pe_inst[31].std__pe__oob_valid          =  std__pe31__oob_valid                      ;
  assign   pe31__std__oob_ready                    =  pe_inst[31].pe__std__oob_ready            ;
  assign   pe_inst[31].std__pe__oob_type           =  std__pe31__oob_type                       ;
  assign   pe_inst[31].std__pe__oob_data           =  std__pe31__oob_data                       ;
  assign   pe_inst[32].sys__pe__allSynchronized    =  sys__pe32__allSynchronized                ;
  assign   pe32__sys__thisSynchronized             =  pe_inst[32].pe__sys__thisSynchronized     ;
  assign   pe32__sys__ready                        =  pe_inst[32].pe__sys__ready                ;
  assign   pe32__sys__complete                     =  pe_inst[32].pe__sys__complete             ;
  assign   pe_inst[32].std__pe__oob_cntl           =  std__pe32__oob_cntl                       ;
  assign   pe_inst[32].std__pe__oob_valid          =  std__pe32__oob_valid                      ;
  assign   pe32__std__oob_ready                    =  pe_inst[32].pe__std__oob_ready            ;
  assign   pe_inst[32].std__pe__oob_type           =  std__pe32__oob_type                       ;
  assign   pe_inst[32].std__pe__oob_data           =  std__pe32__oob_data                       ;
  assign   pe_inst[33].sys__pe__allSynchronized    =  sys__pe33__allSynchronized                ;
  assign   pe33__sys__thisSynchronized             =  pe_inst[33].pe__sys__thisSynchronized     ;
  assign   pe33__sys__ready                        =  pe_inst[33].pe__sys__ready                ;
  assign   pe33__sys__complete                     =  pe_inst[33].pe__sys__complete             ;
  assign   pe_inst[33].std__pe__oob_cntl           =  std__pe33__oob_cntl                       ;
  assign   pe_inst[33].std__pe__oob_valid          =  std__pe33__oob_valid                      ;
  assign   pe33__std__oob_ready                    =  pe_inst[33].pe__std__oob_ready            ;
  assign   pe_inst[33].std__pe__oob_type           =  std__pe33__oob_type                       ;
  assign   pe_inst[33].std__pe__oob_data           =  std__pe33__oob_data                       ;
  assign   pe_inst[34].sys__pe__allSynchronized    =  sys__pe34__allSynchronized                ;
  assign   pe34__sys__thisSynchronized             =  pe_inst[34].pe__sys__thisSynchronized     ;
  assign   pe34__sys__ready                        =  pe_inst[34].pe__sys__ready                ;
  assign   pe34__sys__complete                     =  pe_inst[34].pe__sys__complete             ;
  assign   pe_inst[34].std__pe__oob_cntl           =  std__pe34__oob_cntl                       ;
  assign   pe_inst[34].std__pe__oob_valid          =  std__pe34__oob_valid                      ;
  assign   pe34__std__oob_ready                    =  pe_inst[34].pe__std__oob_ready            ;
  assign   pe_inst[34].std__pe__oob_type           =  std__pe34__oob_type                       ;
  assign   pe_inst[34].std__pe__oob_data           =  std__pe34__oob_data                       ;
  assign   pe_inst[35].sys__pe__allSynchronized    =  sys__pe35__allSynchronized                ;
  assign   pe35__sys__thisSynchronized             =  pe_inst[35].pe__sys__thisSynchronized     ;
  assign   pe35__sys__ready                        =  pe_inst[35].pe__sys__ready                ;
  assign   pe35__sys__complete                     =  pe_inst[35].pe__sys__complete             ;
  assign   pe_inst[35].std__pe__oob_cntl           =  std__pe35__oob_cntl                       ;
  assign   pe_inst[35].std__pe__oob_valid          =  std__pe35__oob_valid                      ;
  assign   pe35__std__oob_ready                    =  pe_inst[35].pe__std__oob_ready            ;
  assign   pe_inst[35].std__pe__oob_type           =  std__pe35__oob_type                       ;
  assign   pe_inst[35].std__pe__oob_data           =  std__pe35__oob_data                       ;
  assign   pe_inst[36].sys__pe__allSynchronized    =  sys__pe36__allSynchronized                ;
  assign   pe36__sys__thisSynchronized             =  pe_inst[36].pe__sys__thisSynchronized     ;
  assign   pe36__sys__ready                        =  pe_inst[36].pe__sys__ready                ;
  assign   pe36__sys__complete                     =  pe_inst[36].pe__sys__complete             ;
  assign   pe_inst[36].std__pe__oob_cntl           =  std__pe36__oob_cntl                       ;
  assign   pe_inst[36].std__pe__oob_valid          =  std__pe36__oob_valid                      ;
  assign   pe36__std__oob_ready                    =  pe_inst[36].pe__std__oob_ready            ;
  assign   pe_inst[36].std__pe__oob_type           =  std__pe36__oob_type                       ;
  assign   pe_inst[36].std__pe__oob_data           =  std__pe36__oob_data                       ;
  assign   pe_inst[37].sys__pe__allSynchronized    =  sys__pe37__allSynchronized                ;
  assign   pe37__sys__thisSynchronized             =  pe_inst[37].pe__sys__thisSynchronized     ;
  assign   pe37__sys__ready                        =  pe_inst[37].pe__sys__ready                ;
  assign   pe37__sys__complete                     =  pe_inst[37].pe__sys__complete             ;
  assign   pe_inst[37].std__pe__oob_cntl           =  std__pe37__oob_cntl                       ;
  assign   pe_inst[37].std__pe__oob_valid          =  std__pe37__oob_valid                      ;
  assign   pe37__std__oob_ready                    =  pe_inst[37].pe__std__oob_ready            ;
  assign   pe_inst[37].std__pe__oob_type           =  std__pe37__oob_type                       ;
  assign   pe_inst[37].std__pe__oob_data           =  std__pe37__oob_data                       ;
  assign   pe_inst[38].sys__pe__allSynchronized    =  sys__pe38__allSynchronized                ;
  assign   pe38__sys__thisSynchronized             =  pe_inst[38].pe__sys__thisSynchronized     ;
  assign   pe38__sys__ready                        =  pe_inst[38].pe__sys__ready                ;
  assign   pe38__sys__complete                     =  pe_inst[38].pe__sys__complete             ;
  assign   pe_inst[38].std__pe__oob_cntl           =  std__pe38__oob_cntl                       ;
  assign   pe_inst[38].std__pe__oob_valid          =  std__pe38__oob_valid                      ;
  assign   pe38__std__oob_ready                    =  pe_inst[38].pe__std__oob_ready            ;
  assign   pe_inst[38].std__pe__oob_type           =  std__pe38__oob_type                       ;
  assign   pe_inst[38].std__pe__oob_data           =  std__pe38__oob_data                       ;
  assign   pe_inst[39].sys__pe__allSynchronized    =  sys__pe39__allSynchronized                ;
  assign   pe39__sys__thisSynchronized             =  pe_inst[39].pe__sys__thisSynchronized     ;
  assign   pe39__sys__ready                        =  pe_inst[39].pe__sys__ready                ;
  assign   pe39__sys__complete                     =  pe_inst[39].pe__sys__complete             ;
  assign   pe_inst[39].std__pe__oob_cntl           =  std__pe39__oob_cntl                       ;
  assign   pe_inst[39].std__pe__oob_valid          =  std__pe39__oob_valid                      ;
  assign   pe39__std__oob_ready                    =  pe_inst[39].pe__std__oob_ready            ;
  assign   pe_inst[39].std__pe__oob_type           =  std__pe39__oob_type                       ;
  assign   pe_inst[39].std__pe__oob_data           =  std__pe39__oob_data                       ;
  assign   pe_inst[40].sys__pe__allSynchronized    =  sys__pe40__allSynchronized                ;
  assign   pe40__sys__thisSynchronized             =  pe_inst[40].pe__sys__thisSynchronized     ;
  assign   pe40__sys__ready                        =  pe_inst[40].pe__sys__ready                ;
  assign   pe40__sys__complete                     =  pe_inst[40].pe__sys__complete             ;
  assign   pe_inst[40].std__pe__oob_cntl           =  std__pe40__oob_cntl                       ;
  assign   pe_inst[40].std__pe__oob_valid          =  std__pe40__oob_valid                      ;
  assign   pe40__std__oob_ready                    =  pe_inst[40].pe__std__oob_ready            ;
  assign   pe_inst[40].std__pe__oob_type           =  std__pe40__oob_type                       ;
  assign   pe_inst[40].std__pe__oob_data           =  std__pe40__oob_data                       ;
  assign   pe_inst[41].sys__pe__allSynchronized    =  sys__pe41__allSynchronized                ;
  assign   pe41__sys__thisSynchronized             =  pe_inst[41].pe__sys__thisSynchronized     ;
  assign   pe41__sys__ready                        =  pe_inst[41].pe__sys__ready                ;
  assign   pe41__sys__complete                     =  pe_inst[41].pe__sys__complete             ;
  assign   pe_inst[41].std__pe__oob_cntl           =  std__pe41__oob_cntl                       ;
  assign   pe_inst[41].std__pe__oob_valid          =  std__pe41__oob_valid                      ;
  assign   pe41__std__oob_ready                    =  pe_inst[41].pe__std__oob_ready            ;
  assign   pe_inst[41].std__pe__oob_type           =  std__pe41__oob_type                       ;
  assign   pe_inst[41].std__pe__oob_data           =  std__pe41__oob_data                       ;
  assign   pe_inst[42].sys__pe__allSynchronized    =  sys__pe42__allSynchronized                ;
  assign   pe42__sys__thisSynchronized             =  pe_inst[42].pe__sys__thisSynchronized     ;
  assign   pe42__sys__ready                        =  pe_inst[42].pe__sys__ready                ;
  assign   pe42__sys__complete                     =  pe_inst[42].pe__sys__complete             ;
  assign   pe_inst[42].std__pe__oob_cntl           =  std__pe42__oob_cntl                       ;
  assign   pe_inst[42].std__pe__oob_valid          =  std__pe42__oob_valid                      ;
  assign   pe42__std__oob_ready                    =  pe_inst[42].pe__std__oob_ready            ;
  assign   pe_inst[42].std__pe__oob_type           =  std__pe42__oob_type                       ;
  assign   pe_inst[42].std__pe__oob_data           =  std__pe42__oob_data                       ;
  assign   pe_inst[43].sys__pe__allSynchronized    =  sys__pe43__allSynchronized                ;
  assign   pe43__sys__thisSynchronized             =  pe_inst[43].pe__sys__thisSynchronized     ;
  assign   pe43__sys__ready                        =  pe_inst[43].pe__sys__ready                ;
  assign   pe43__sys__complete                     =  pe_inst[43].pe__sys__complete             ;
  assign   pe_inst[43].std__pe__oob_cntl           =  std__pe43__oob_cntl                       ;
  assign   pe_inst[43].std__pe__oob_valid          =  std__pe43__oob_valid                      ;
  assign   pe43__std__oob_ready                    =  pe_inst[43].pe__std__oob_ready            ;
  assign   pe_inst[43].std__pe__oob_type           =  std__pe43__oob_type                       ;
  assign   pe_inst[43].std__pe__oob_data           =  std__pe43__oob_data                       ;
  assign   pe_inst[44].sys__pe__allSynchronized    =  sys__pe44__allSynchronized                ;
  assign   pe44__sys__thisSynchronized             =  pe_inst[44].pe__sys__thisSynchronized     ;
  assign   pe44__sys__ready                        =  pe_inst[44].pe__sys__ready                ;
  assign   pe44__sys__complete                     =  pe_inst[44].pe__sys__complete             ;
  assign   pe_inst[44].std__pe__oob_cntl           =  std__pe44__oob_cntl                       ;
  assign   pe_inst[44].std__pe__oob_valid          =  std__pe44__oob_valid                      ;
  assign   pe44__std__oob_ready                    =  pe_inst[44].pe__std__oob_ready            ;
  assign   pe_inst[44].std__pe__oob_type           =  std__pe44__oob_type                       ;
  assign   pe_inst[44].std__pe__oob_data           =  std__pe44__oob_data                       ;
  assign   pe_inst[45].sys__pe__allSynchronized    =  sys__pe45__allSynchronized                ;
  assign   pe45__sys__thisSynchronized             =  pe_inst[45].pe__sys__thisSynchronized     ;
  assign   pe45__sys__ready                        =  pe_inst[45].pe__sys__ready                ;
  assign   pe45__sys__complete                     =  pe_inst[45].pe__sys__complete             ;
  assign   pe_inst[45].std__pe__oob_cntl           =  std__pe45__oob_cntl                       ;
  assign   pe_inst[45].std__pe__oob_valid          =  std__pe45__oob_valid                      ;
  assign   pe45__std__oob_ready                    =  pe_inst[45].pe__std__oob_ready            ;
  assign   pe_inst[45].std__pe__oob_type           =  std__pe45__oob_type                       ;
  assign   pe_inst[45].std__pe__oob_data           =  std__pe45__oob_data                       ;
  assign   pe_inst[46].sys__pe__allSynchronized    =  sys__pe46__allSynchronized                ;
  assign   pe46__sys__thisSynchronized             =  pe_inst[46].pe__sys__thisSynchronized     ;
  assign   pe46__sys__ready                        =  pe_inst[46].pe__sys__ready                ;
  assign   pe46__sys__complete                     =  pe_inst[46].pe__sys__complete             ;
  assign   pe_inst[46].std__pe__oob_cntl           =  std__pe46__oob_cntl                       ;
  assign   pe_inst[46].std__pe__oob_valid          =  std__pe46__oob_valid                      ;
  assign   pe46__std__oob_ready                    =  pe_inst[46].pe__std__oob_ready            ;
  assign   pe_inst[46].std__pe__oob_type           =  std__pe46__oob_type                       ;
  assign   pe_inst[46].std__pe__oob_data           =  std__pe46__oob_data                       ;
  assign   pe_inst[47].sys__pe__allSynchronized    =  sys__pe47__allSynchronized                ;
  assign   pe47__sys__thisSynchronized             =  pe_inst[47].pe__sys__thisSynchronized     ;
  assign   pe47__sys__ready                        =  pe_inst[47].pe__sys__ready                ;
  assign   pe47__sys__complete                     =  pe_inst[47].pe__sys__complete             ;
  assign   pe_inst[47].std__pe__oob_cntl           =  std__pe47__oob_cntl                       ;
  assign   pe_inst[47].std__pe__oob_valid          =  std__pe47__oob_valid                      ;
  assign   pe47__std__oob_ready                    =  pe_inst[47].pe__std__oob_ready            ;
  assign   pe_inst[47].std__pe__oob_type           =  std__pe47__oob_type                       ;
  assign   pe_inst[47].std__pe__oob_data           =  std__pe47__oob_data                       ;
  assign   pe_inst[48].sys__pe__allSynchronized    =  sys__pe48__allSynchronized                ;
  assign   pe48__sys__thisSynchronized             =  pe_inst[48].pe__sys__thisSynchronized     ;
  assign   pe48__sys__ready                        =  pe_inst[48].pe__sys__ready                ;
  assign   pe48__sys__complete                     =  pe_inst[48].pe__sys__complete             ;
  assign   pe_inst[48].std__pe__oob_cntl           =  std__pe48__oob_cntl                       ;
  assign   pe_inst[48].std__pe__oob_valid          =  std__pe48__oob_valid                      ;
  assign   pe48__std__oob_ready                    =  pe_inst[48].pe__std__oob_ready            ;
  assign   pe_inst[48].std__pe__oob_type           =  std__pe48__oob_type                       ;
  assign   pe_inst[48].std__pe__oob_data           =  std__pe48__oob_data                       ;
  assign   pe_inst[49].sys__pe__allSynchronized    =  sys__pe49__allSynchronized                ;
  assign   pe49__sys__thisSynchronized             =  pe_inst[49].pe__sys__thisSynchronized     ;
  assign   pe49__sys__ready                        =  pe_inst[49].pe__sys__ready                ;
  assign   pe49__sys__complete                     =  pe_inst[49].pe__sys__complete             ;
  assign   pe_inst[49].std__pe__oob_cntl           =  std__pe49__oob_cntl                       ;
  assign   pe_inst[49].std__pe__oob_valid          =  std__pe49__oob_valid                      ;
  assign   pe49__std__oob_ready                    =  pe_inst[49].pe__std__oob_ready            ;
  assign   pe_inst[49].std__pe__oob_type           =  std__pe49__oob_type                       ;
  assign   pe_inst[49].std__pe__oob_data           =  std__pe49__oob_data                       ;
  assign   pe_inst[50].sys__pe__allSynchronized    =  sys__pe50__allSynchronized                ;
  assign   pe50__sys__thisSynchronized             =  pe_inst[50].pe__sys__thisSynchronized     ;
  assign   pe50__sys__ready                        =  pe_inst[50].pe__sys__ready                ;
  assign   pe50__sys__complete                     =  pe_inst[50].pe__sys__complete             ;
  assign   pe_inst[50].std__pe__oob_cntl           =  std__pe50__oob_cntl                       ;
  assign   pe_inst[50].std__pe__oob_valid          =  std__pe50__oob_valid                      ;
  assign   pe50__std__oob_ready                    =  pe_inst[50].pe__std__oob_ready            ;
  assign   pe_inst[50].std__pe__oob_type           =  std__pe50__oob_type                       ;
  assign   pe_inst[50].std__pe__oob_data           =  std__pe50__oob_data                       ;
  assign   pe_inst[51].sys__pe__allSynchronized    =  sys__pe51__allSynchronized                ;
  assign   pe51__sys__thisSynchronized             =  pe_inst[51].pe__sys__thisSynchronized     ;
  assign   pe51__sys__ready                        =  pe_inst[51].pe__sys__ready                ;
  assign   pe51__sys__complete                     =  pe_inst[51].pe__sys__complete             ;
  assign   pe_inst[51].std__pe__oob_cntl           =  std__pe51__oob_cntl                       ;
  assign   pe_inst[51].std__pe__oob_valid          =  std__pe51__oob_valid                      ;
  assign   pe51__std__oob_ready                    =  pe_inst[51].pe__std__oob_ready            ;
  assign   pe_inst[51].std__pe__oob_type           =  std__pe51__oob_type                       ;
  assign   pe_inst[51].std__pe__oob_data           =  std__pe51__oob_data                       ;
  assign   pe_inst[52].sys__pe__allSynchronized    =  sys__pe52__allSynchronized                ;
  assign   pe52__sys__thisSynchronized             =  pe_inst[52].pe__sys__thisSynchronized     ;
  assign   pe52__sys__ready                        =  pe_inst[52].pe__sys__ready                ;
  assign   pe52__sys__complete                     =  pe_inst[52].pe__sys__complete             ;
  assign   pe_inst[52].std__pe__oob_cntl           =  std__pe52__oob_cntl                       ;
  assign   pe_inst[52].std__pe__oob_valid          =  std__pe52__oob_valid                      ;
  assign   pe52__std__oob_ready                    =  pe_inst[52].pe__std__oob_ready            ;
  assign   pe_inst[52].std__pe__oob_type           =  std__pe52__oob_type                       ;
  assign   pe_inst[52].std__pe__oob_data           =  std__pe52__oob_data                       ;
  assign   pe_inst[53].sys__pe__allSynchronized    =  sys__pe53__allSynchronized                ;
  assign   pe53__sys__thisSynchronized             =  pe_inst[53].pe__sys__thisSynchronized     ;
  assign   pe53__sys__ready                        =  pe_inst[53].pe__sys__ready                ;
  assign   pe53__sys__complete                     =  pe_inst[53].pe__sys__complete             ;
  assign   pe_inst[53].std__pe__oob_cntl           =  std__pe53__oob_cntl                       ;
  assign   pe_inst[53].std__pe__oob_valid          =  std__pe53__oob_valid                      ;
  assign   pe53__std__oob_ready                    =  pe_inst[53].pe__std__oob_ready            ;
  assign   pe_inst[53].std__pe__oob_type           =  std__pe53__oob_type                       ;
  assign   pe_inst[53].std__pe__oob_data           =  std__pe53__oob_data                       ;
  assign   pe_inst[54].sys__pe__allSynchronized    =  sys__pe54__allSynchronized                ;
  assign   pe54__sys__thisSynchronized             =  pe_inst[54].pe__sys__thisSynchronized     ;
  assign   pe54__sys__ready                        =  pe_inst[54].pe__sys__ready                ;
  assign   pe54__sys__complete                     =  pe_inst[54].pe__sys__complete             ;
  assign   pe_inst[54].std__pe__oob_cntl           =  std__pe54__oob_cntl                       ;
  assign   pe_inst[54].std__pe__oob_valid          =  std__pe54__oob_valid                      ;
  assign   pe54__std__oob_ready                    =  pe_inst[54].pe__std__oob_ready            ;
  assign   pe_inst[54].std__pe__oob_type           =  std__pe54__oob_type                       ;
  assign   pe_inst[54].std__pe__oob_data           =  std__pe54__oob_data                       ;
  assign   pe_inst[55].sys__pe__allSynchronized    =  sys__pe55__allSynchronized                ;
  assign   pe55__sys__thisSynchronized             =  pe_inst[55].pe__sys__thisSynchronized     ;
  assign   pe55__sys__ready                        =  pe_inst[55].pe__sys__ready                ;
  assign   pe55__sys__complete                     =  pe_inst[55].pe__sys__complete             ;
  assign   pe_inst[55].std__pe__oob_cntl           =  std__pe55__oob_cntl                       ;
  assign   pe_inst[55].std__pe__oob_valid          =  std__pe55__oob_valid                      ;
  assign   pe55__std__oob_ready                    =  pe_inst[55].pe__std__oob_ready            ;
  assign   pe_inst[55].std__pe__oob_type           =  std__pe55__oob_type                       ;
  assign   pe_inst[55].std__pe__oob_data           =  std__pe55__oob_data                       ;
  assign   pe_inst[56].sys__pe__allSynchronized    =  sys__pe56__allSynchronized                ;
  assign   pe56__sys__thisSynchronized             =  pe_inst[56].pe__sys__thisSynchronized     ;
  assign   pe56__sys__ready                        =  pe_inst[56].pe__sys__ready                ;
  assign   pe56__sys__complete                     =  pe_inst[56].pe__sys__complete             ;
  assign   pe_inst[56].std__pe__oob_cntl           =  std__pe56__oob_cntl                       ;
  assign   pe_inst[56].std__pe__oob_valid          =  std__pe56__oob_valid                      ;
  assign   pe56__std__oob_ready                    =  pe_inst[56].pe__std__oob_ready            ;
  assign   pe_inst[56].std__pe__oob_type           =  std__pe56__oob_type                       ;
  assign   pe_inst[56].std__pe__oob_data           =  std__pe56__oob_data                       ;
  assign   pe_inst[57].sys__pe__allSynchronized    =  sys__pe57__allSynchronized                ;
  assign   pe57__sys__thisSynchronized             =  pe_inst[57].pe__sys__thisSynchronized     ;
  assign   pe57__sys__ready                        =  pe_inst[57].pe__sys__ready                ;
  assign   pe57__sys__complete                     =  pe_inst[57].pe__sys__complete             ;
  assign   pe_inst[57].std__pe__oob_cntl           =  std__pe57__oob_cntl                       ;
  assign   pe_inst[57].std__pe__oob_valid          =  std__pe57__oob_valid                      ;
  assign   pe57__std__oob_ready                    =  pe_inst[57].pe__std__oob_ready            ;
  assign   pe_inst[57].std__pe__oob_type           =  std__pe57__oob_type                       ;
  assign   pe_inst[57].std__pe__oob_data           =  std__pe57__oob_data                       ;
  assign   pe_inst[58].sys__pe__allSynchronized    =  sys__pe58__allSynchronized                ;
  assign   pe58__sys__thisSynchronized             =  pe_inst[58].pe__sys__thisSynchronized     ;
  assign   pe58__sys__ready                        =  pe_inst[58].pe__sys__ready                ;
  assign   pe58__sys__complete                     =  pe_inst[58].pe__sys__complete             ;
  assign   pe_inst[58].std__pe__oob_cntl           =  std__pe58__oob_cntl                       ;
  assign   pe_inst[58].std__pe__oob_valid          =  std__pe58__oob_valid                      ;
  assign   pe58__std__oob_ready                    =  pe_inst[58].pe__std__oob_ready            ;
  assign   pe_inst[58].std__pe__oob_type           =  std__pe58__oob_type                       ;
  assign   pe_inst[58].std__pe__oob_data           =  std__pe58__oob_data                       ;
  assign   pe_inst[59].sys__pe__allSynchronized    =  sys__pe59__allSynchronized                ;
  assign   pe59__sys__thisSynchronized             =  pe_inst[59].pe__sys__thisSynchronized     ;
  assign   pe59__sys__ready                        =  pe_inst[59].pe__sys__ready                ;
  assign   pe59__sys__complete                     =  pe_inst[59].pe__sys__complete             ;
  assign   pe_inst[59].std__pe__oob_cntl           =  std__pe59__oob_cntl                       ;
  assign   pe_inst[59].std__pe__oob_valid          =  std__pe59__oob_valid                      ;
  assign   pe59__std__oob_ready                    =  pe_inst[59].pe__std__oob_ready            ;
  assign   pe_inst[59].std__pe__oob_type           =  std__pe59__oob_type                       ;
  assign   pe_inst[59].std__pe__oob_data           =  std__pe59__oob_data                       ;
  assign   pe_inst[60].sys__pe__allSynchronized    =  sys__pe60__allSynchronized                ;
  assign   pe60__sys__thisSynchronized             =  pe_inst[60].pe__sys__thisSynchronized     ;
  assign   pe60__sys__ready                        =  pe_inst[60].pe__sys__ready                ;
  assign   pe60__sys__complete                     =  pe_inst[60].pe__sys__complete             ;
  assign   pe_inst[60].std__pe__oob_cntl           =  std__pe60__oob_cntl                       ;
  assign   pe_inst[60].std__pe__oob_valid          =  std__pe60__oob_valid                      ;
  assign   pe60__std__oob_ready                    =  pe_inst[60].pe__std__oob_ready            ;
  assign   pe_inst[60].std__pe__oob_type           =  std__pe60__oob_type                       ;
  assign   pe_inst[60].std__pe__oob_data           =  std__pe60__oob_data                       ;
  assign   pe_inst[61].sys__pe__allSynchronized    =  sys__pe61__allSynchronized                ;
  assign   pe61__sys__thisSynchronized             =  pe_inst[61].pe__sys__thisSynchronized     ;
  assign   pe61__sys__ready                        =  pe_inst[61].pe__sys__ready                ;
  assign   pe61__sys__complete                     =  pe_inst[61].pe__sys__complete             ;
  assign   pe_inst[61].std__pe__oob_cntl           =  std__pe61__oob_cntl                       ;
  assign   pe_inst[61].std__pe__oob_valid          =  std__pe61__oob_valid                      ;
  assign   pe61__std__oob_ready                    =  pe_inst[61].pe__std__oob_ready            ;
  assign   pe_inst[61].std__pe__oob_type           =  std__pe61__oob_type                       ;
  assign   pe_inst[61].std__pe__oob_data           =  std__pe61__oob_data                       ;
  assign   pe_inst[62].sys__pe__allSynchronized    =  sys__pe62__allSynchronized                ;
  assign   pe62__sys__thisSynchronized             =  pe_inst[62].pe__sys__thisSynchronized     ;
  assign   pe62__sys__ready                        =  pe_inst[62].pe__sys__ready                ;
  assign   pe62__sys__complete                     =  pe_inst[62].pe__sys__complete             ;
  assign   pe_inst[62].std__pe__oob_cntl           =  std__pe62__oob_cntl                       ;
  assign   pe_inst[62].std__pe__oob_valid          =  std__pe62__oob_valid                      ;
  assign   pe62__std__oob_ready                    =  pe_inst[62].pe__std__oob_ready            ;
  assign   pe_inst[62].std__pe__oob_type           =  std__pe62__oob_type                       ;
  assign   pe_inst[62].std__pe__oob_data           =  std__pe62__oob_data                       ;
  assign   pe_inst[63].sys__pe__allSynchronized    =  sys__pe63__allSynchronized                ;
  assign   pe63__sys__thisSynchronized             =  pe_inst[63].pe__sys__thisSynchronized     ;
  assign   pe63__sys__ready                        =  pe_inst[63].pe__sys__ready                ;
  assign   pe63__sys__complete                     =  pe_inst[63].pe__sys__complete             ;
  assign   pe_inst[63].std__pe__oob_cntl           =  std__pe63__oob_cntl                       ;
  assign   pe_inst[63].std__pe__oob_valid          =  std__pe63__oob_valid                      ;
  assign   pe63__std__oob_ready                    =  pe_inst[63].pe__std__oob_ready            ;
  assign   pe_inst[63].std__pe__oob_type           =  std__pe63__oob_type                       ;
  assign   pe_inst[63].std__pe__oob_data           =  std__pe63__oob_data                       ;
