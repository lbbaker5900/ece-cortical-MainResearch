
            .std__mgr0__lane0_strm0_ready           ( std__mgr0__lane0_strm0_ready       ),
            .mgr0__std__lane0_strm0_cntl            ( mgr0__std__lane0_strm0_cntl        ),
            .mgr0__std__lane0_strm0_data            ( mgr0__std__lane0_strm0_data        ),
            .mgr0__std__lane0_strm0_data_valid      ( mgr0__std__lane0_strm0_data_valid  ),

            .std__mgr0__lane0_strm1_ready           ( std__mgr0__lane0_strm1_ready       ),
            .mgr0__std__lane0_strm1_cntl            ( mgr0__std__lane0_strm1_cntl        ),
            .mgr0__std__lane0_strm1_data            ( mgr0__std__lane0_strm1_data        ),
            .mgr0__std__lane0_strm1_data_valid      ( mgr0__std__lane0_strm1_data_valid  ),

            .std__mgr0__lane1_strm0_ready           ( std__mgr0__lane1_strm0_ready       ),
            .mgr0__std__lane1_strm0_cntl            ( mgr0__std__lane1_strm0_cntl        ),
            .mgr0__std__lane1_strm0_data            ( mgr0__std__lane1_strm0_data        ),
            .mgr0__std__lane1_strm0_data_valid      ( mgr0__std__lane1_strm0_data_valid  ),

            .std__mgr0__lane1_strm1_ready           ( std__mgr0__lane1_strm1_ready       ),
            .mgr0__std__lane1_strm1_cntl            ( mgr0__std__lane1_strm1_cntl        ),
            .mgr0__std__lane1_strm1_data            ( mgr0__std__lane1_strm1_data        ),
            .mgr0__std__lane1_strm1_data_valid      ( mgr0__std__lane1_strm1_data_valid  ),

            .std__mgr0__lane2_strm0_ready           ( std__mgr0__lane2_strm0_ready       ),
            .mgr0__std__lane2_strm0_cntl            ( mgr0__std__lane2_strm0_cntl        ),
            .mgr0__std__lane2_strm0_data            ( mgr0__std__lane2_strm0_data        ),
            .mgr0__std__lane2_strm0_data_valid      ( mgr0__std__lane2_strm0_data_valid  ),

            .std__mgr0__lane2_strm1_ready           ( std__mgr0__lane2_strm1_ready       ),
            .mgr0__std__lane2_strm1_cntl            ( mgr0__std__lane2_strm1_cntl        ),
            .mgr0__std__lane2_strm1_data            ( mgr0__std__lane2_strm1_data        ),
            .mgr0__std__lane2_strm1_data_valid      ( mgr0__std__lane2_strm1_data_valid  ),

            .std__mgr0__lane3_strm0_ready           ( std__mgr0__lane3_strm0_ready       ),
            .mgr0__std__lane3_strm0_cntl            ( mgr0__std__lane3_strm0_cntl        ),
            .mgr0__std__lane3_strm0_data            ( mgr0__std__lane3_strm0_data        ),
            .mgr0__std__lane3_strm0_data_valid      ( mgr0__std__lane3_strm0_data_valid  ),

            .std__mgr0__lane3_strm1_ready           ( std__mgr0__lane3_strm1_ready       ),
            .mgr0__std__lane3_strm1_cntl            ( mgr0__std__lane3_strm1_cntl        ),
            .mgr0__std__lane3_strm1_data            ( mgr0__std__lane3_strm1_data        ),
            .mgr0__std__lane3_strm1_data_valid      ( mgr0__std__lane3_strm1_data_valid  ),

            .std__mgr0__lane4_strm0_ready           ( std__mgr0__lane4_strm0_ready       ),
            .mgr0__std__lane4_strm0_cntl            ( mgr0__std__lane4_strm0_cntl        ),
            .mgr0__std__lane4_strm0_data            ( mgr0__std__lane4_strm0_data        ),
            .mgr0__std__lane4_strm0_data_valid      ( mgr0__std__lane4_strm0_data_valid  ),

            .std__mgr0__lane4_strm1_ready           ( std__mgr0__lane4_strm1_ready       ),
            .mgr0__std__lane4_strm1_cntl            ( mgr0__std__lane4_strm1_cntl        ),
            .mgr0__std__lane4_strm1_data            ( mgr0__std__lane4_strm1_data        ),
            .mgr0__std__lane4_strm1_data_valid      ( mgr0__std__lane4_strm1_data_valid  ),

            .std__mgr0__lane5_strm0_ready           ( std__mgr0__lane5_strm0_ready       ),
            .mgr0__std__lane5_strm0_cntl            ( mgr0__std__lane5_strm0_cntl        ),
            .mgr0__std__lane5_strm0_data            ( mgr0__std__lane5_strm0_data        ),
            .mgr0__std__lane5_strm0_data_valid      ( mgr0__std__lane5_strm0_data_valid  ),

            .std__mgr0__lane5_strm1_ready           ( std__mgr0__lane5_strm1_ready       ),
            .mgr0__std__lane5_strm1_cntl            ( mgr0__std__lane5_strm1_cntl        ),
            .mgr0__std__lane5_strm1_data            ( mgr0__std__lane5_strm1_data        ),
            .mgr0__std__lane5_strm1_data_valid      ( mgr0__std__lane5_strm1_data_valid  ),

            .std__mgr0__lane6_strm0_ready           ( std__mgr0__lane6_strm0_ready       ),
            .mgr0__std__lane6_strm0_cntl            ( mgr0__std__lane6_strm0_cntl        ),
            .mgr0__std__lane6_strm0_data            ( mgr0__std__lane6_strm0_data        ),
            .mgr0__std__lane6_strm0_data_valid      ( mgr0__std__lane6_strm0_data_valid  ),

            .std__mgr0__lane6_strm1_ready           ( std__mgr0__lane6_strm1_ready       ),
            .mgr0__std__lane6_strm1_cntl            ( mgr0__std__lane6_strm1_cntl        ),
            .mgr0__std__lane6_strm1_data            ( mgr0__std__lane6_strm1_data        ),
            .mgr0__std__lane6_strm1_data_valid      ( mgr0__std__lane6_strm1_data_valid  ),

            .std__mgr0__lane7_strm0_ready           ( std__mgr0__lane7_strm0_ready       ),
            .mgr0__std__lane7_strm0_cntl            ( mgr0__std__lane7_strm0_cntl        ),
            .mgr0__std__lane7_strm0_data            ( mgr0__std__lane7_strm0_data        ),
            .mgr0__std__lane7_strm0_data_valid      ( mgr0__std__lane7_strm0_data_valid  ),

            .std__mgr0__lane7_strm1_ready           ( std__mgr0__lane7_strm1_ready       ),
            .mgr0__std__lane7_strm1_cntl            ( mgr0__std__lane7_strm1_cntl        ),
            .mgr0__std__lane7_strm1_data            ( mgr0__std__lane7_strm1_data        ),
            .mgr0__std__lane7_strm1_data_valid      ( mgr0__std__lane7_strm1_data_valid  ),

            .std__mgr0__lane8_strm0_ready           ( std__mgr0__lane8_strm0_ready       ),
            .mgr0__std__lane8_strm0_cntl            ( mgr0__std__lane8_strm0_cntl        ),
            .mgr0__std__lane8_strm0_data            ( mgr0__std__lane8_strm0_data        ),
            .mgr0__std__lane8_strm0_data_valid      ( mgr0__std__lane8_strm0_data_valid  ),

            .std__mgr0__lane8_strm1_ready           ( std__mgr0__lane8_strm1_ready       ),
            .mgr0__std__lane8_strm1_cntl            ( mgr0__std__lane8_strm1_cntl        ),
            .mgr0__std__lane8_strm1_data            ( mgr0__std__lane8_strm1_data        ),
            .mgr0__std__lane8_strm1_data_valid      ( mgr0__std__lane8_strm1_data_valid  ),

            .std__mgr0__lane9_strm0_ready           ( std__mgr0__lane9_strm0_ready       ),
            .mgr0__std__lane9_strm0_cntl            ( mgr0__std__lane9_strm0_cntl        ),
            .mgr0__std__lane9_strm0_data            ( mgr0__std__lane9_strm0_data        ),
            .mgr0__std__lane9_strm0_data_valid      ( mgr0__std__lane9_strm0_data_valid  ),

            .std__mgr0__lane9_strm1_ready           ( std__mgr0__lane9_strm1_ready       ),
            .mgr0__std__lane9_strm1_cntl            ( mgr0__std__lane9_strm1_cntl        ),
            .mgr0__std__lane9_strm1_data            ( mgr0__std__lane9_strm1_data        ),
            .mgr0__std__lane9_strm1_data_valid      ( mgr0__std__lane9_strm1_data_valid  ),

            .std__mgr0__lane10_strm0_ready           ( std__mgr0__lane10_strm0_ready       ),
            .mgr0__std__lane10_strm0_cntl            ( mgr0__std__lane10_strm0_cntl        ),
            .mgr0__std__lane10_strm0_data            ( mgr0__std__lane10_strm0_data        ),
            .mgr0__std__lane10_strm0_data_valid      ( mgr0__std__lane10_strm0_data_valid  ),

            .std__mgr0__lane10_strm1_ready           ( std__mgr0__lane10_strm1_ready       ),
            .mgr0__std__lane10_strm1_cntl            ( mgr0__std__lane10_strm1_cntl        ),
            .mgr0__std__lane10_strm1_data            ( mgr0__std__lane10_strm1_data        ),
            .mgr0__std__lane10_strm1_data_valid      ( mgr0__std__lane10_strm1_data_valid  ),

            .std__mgr0__lane11_strm0_ready           ( std__mgr0__lane11_strm0_ready       ),
            .mgr0__std__lane11_strm0_cntl            ( mgr0__std__lane11_strm0_cntl        ),
            .mgr0__std__lane11_strm0_data            ( mgr0__std__lane11_strm0_data        ),
            .mgr0__std__lane11_strm0_data_valid      ( mgr0__std__lane11_strm0_data_valid  ),

            .std__mgr0__lane11_strm1_ready           ( std__mgr0__lane11_strm1_ready       ),
            .mgr0__std__lane11_strm1_cntl            ( mgr0__std__lane11_strm1_cntl        ),
            .mgr0__std__lane11_strm1_data            ( mgr0__std__lane11_strm1_data        ),
            .mgr0__std__lane11_strm1_data_valid      ( mgr0__std__lane11_strm1_data_valid  ),

            .std__mgr0__lane12_strm0_ready           ( std__mgr0__lane12_strm0_ready       ),
            .mgr0__std__lane12_strm0_cntl            ( mgr0__std__lane12_strm0_cntl        ),
            .mgr0__std__lane12_strm0_data            ( mgr0__std__lane12_strm0_data        ),
            .mgr0__std__lane12_strm0_data_valid      ( mgr0__std__lane12_strm0_data_valid  ),

            .std__mgr0__lane12_strm1_ready           ( std__mgr0__lane12_strm1_ready       ),
            .mgr0__std__lane12_strm1_cntl            ( mgr0__std__lane12_strm1_cntl        ),
            .mgr0__std__lane12_strm1_data            ( mgr0__std__lane12_strm1_data        ),
            .mgr0__std__lane12_strm1_data_valid      ( mgr0__std__lane12_strm1_data_valid  ),

            .std__mgr0__lane13_strm0_ready           ( std__mgr0__lane13_strm0_ready       ),
            .mgr0__std__lane13_strm0_cntl            ( mgr0__std__lane13_strm0_cntl        ),
            .mgr0__std__lane13_strm0_data            ( mgr0__std__lane13_strm0_data        ),
            .mgr0__std__lane13_strm0_data_valid      ( mgr0__std__lane13_strm0_data_valid  ),

            .std__mgr0__lane13_strm1_ready           ( std__mgr0__lane13_strm1_ready       ),
            .mgr0__std__lane13_strm1_cntl            ( mgr0__std__lane13_strm1_cntl        ),
            .mgr0__std__lane13_strm1_data            ( mgr0__std__lane13_strm1_data        ),
            .mgr0__std__lane13_strm1_data_valid      ( mgr0__std__lane13_strm1_data_valid  ),

            .std__mgr0__lane14_strm0_ready           ( std__mgr0__lane14_strm0_ready       ),
            .mgr0__std__lane14_strm0_cntl            ( mgr0__std__lane14_strm0_cntl        ),
            .mgr0__std__lane14_strm0_data            ( mgr0__std__lane14_strm0_data        ),
            .mgr0__std__lane14_strm0_data_valid      ( mgr0__std__lane14_strm0_data_valid  ),

            .std__mgr0__lane14_strm1_ready           ( std__mgr0__lane14_strm1_ready       ),
            .mgr0__std__lane14_strm1_cntl            ( mgr0__std__lane14_strm1_cntl        ),
            .mgr0__std__lane14_strm1_data            ( mgr0__std__lane14_strm1_data        ),
            .mgr0__std__lane14_strm1_data_valid      ( mgr0__std__lane14_strm1_data_valid  ),

            .std__mgr0__lane15_strm0_ready           ( std__mgr0__lane15_strm0_ready       ),
            .mgr0__std__lane15_strm0_cntl            ( mgr0__std__lane15_strm0_cntl        ),
            .mgr0__std__lane15_strm0_data            ( mgr0__std__lane15_strm0_data        ),
            .mgr0__std__lane15_strm0_data_valid      ( mgr0__std__lane15_strm0_data_valid  ),

            .std__mgr0__lane15_strm1_ready           ( std__mgr0__lane15_strm1_ready       ),
            .mgr0__std__lane15_strm1_cntl            ( mgr0__std__lane15_strm1_cntl        ),
            .mgr0__std__lane15_strm1_data            ( mgr0__std__lane15_strm1_data        ),
            .mgr0__std__lane15_strm1_data_valid      ( mgr0__std__lane15_strm1_data_valid  ),

            .std__mgr0__lane16_strm0_ready           ( std__mgr0__lane16_strm0_ready       ),
            .mgr0__std__lane16_strm0_cntl            ( mgr0__std__lane16_strm0_cntl        ),
            .mgr0__std__lane16_strm0_data            ( mgr0__std__lane16_strm0_data        ),
            .mgr0__std__lane16_strm0_data_valid      ( mgr0__std__lane16_strm0_data_valid  ),

            .std__mgr0__lane16_strm1_ready           ( std__mgr0__lane16_strm1_ready       ),
            .mgr0__std__lane16_strm1_cntl            ( mgr0__std__lane16_strm1_cntl        ),
            .mgr0__std__lane16_strm1_data            ( mgr0__std__lane16_strm1_data        ),
            .mgr0__std__lane16_strm1_data_valid      ( mgr0__std__lane16_strm1_data_valid  ),

            .std__mgr0__lane17_strm0_ready           ( std__mgr0__lane17_strm0_ready       ),
            .mgr0__std__lane17_strm0_cntl            ( mgr0__std__lane17_strm0_cntl        ),
            .mgr0__std__lane17_strm0_data            ( mgr0__std__lane17_strm0_data        ),
            .mgr0__std__lane17_strm0_data_valid      ( mgr0__std__lane17_strm0_data_valid  ),

            .std__mgr0__lane17_strm1_ready           ( std__mgr0__lane17_strm1_ready       ),
            .mgr0__std__lane17_strm1_cntl            ( mgr0__std__lane17_strm1_cntl        ),
            .mgr0__std__lane17_strm1_data            ( mgr0__std__lane17_strm1_data        ),
            .mgr0__std__lane17_strm1_data_valid      ( mgr0__std__lane17_strm1_data_valid  ),

            .std__mgr0__lane18_strm0_ready           ( std__mgr0__lane18_strm0_ready       ),
            .mgr0__std__lane18_strm0_cntl            ( mgr0__std__lane18_strm0_cntl        ),
            .mgr0__std__lane18_strm0_data            ( mgr0__std__lane18_strm0_data        ),
            .mgr0__std__lane18_strm0_data_valid      ( mgr0__std__lane18_strm0_data_valid  ),

            .std__mgr0__lane18_strm1_ready           ( std__mgr0__lane18_strm1_ready       ),
            .mgr0__std__lane18_strm1_cntl            ( mgr0__std__lane18_strm1_cntl        ),
            .mgr0__std__lane18_strm1_data            ( mgr0__std__lane18_strm1_data        ),
            .mgr0__std__lane18_strm1_data_valid      ( mgr0__std__lane18_strm1_data_valid  ),

            .std__mgr0__lane19_strm0_ready           ( std__mgr0__lane19_strm0_ready       ),
            .mgr0__std__lane19_strm0_cntl            ( mgr0__std__lane19_strm0_cntl        ),
            .mgr0__std__lane19_strm0_data            ( mgr0__std__lane19_strm0_data        ),
            .mgr0__std__lane19_strm0_data_valid      ( mgr0__std__lane19_strm0_data_valid  ),

            .std__mgr0__lane19_strm1_ready           ( std__mgr0__lane19_strm1_ready       ),
            .mgr0__std__lane19_strm1_cntl            ( mgr0__std__lane19_strm1_cntl        ),
            .mgr0__std__lane19_strm1_data            ( mgr0__std__lane19_strm1_data        ),
            .mgr0__std__lane19_strm1_data_valid      ( mgr0__std__lane19_strm1_data_valid  ),

            .std__mgr0__lane20_strm0_ready           ( std__mgr0__lane20_strm0_ready       ),
            .mgr0__std__lane20_strm0_cntl            ( mgr0__std__lane20_strm0_cntl        ),
            .mgr0__std__lane20_strm0_data            ( mgr0__std__lane20_strm0_data        ),
            .mgr0__std__lane20_strm0_data_valid      ( mgr0__std__lane20_strm0_data_valid  ),

            .std__mgr0__lane20_strm1_ready           ( std__mgr0__lane20_strm1_ready       ),
            .mgr0__std__lane20_strm1_cntl            ( mgr0__std__lane20_strm1_cntl        ),
            .mgr0__std__lane20_strm1_data            ( mgr0__std__lane20_strm1_data        ),
            .mgr0__std__lane20_strm1_data_valid      ( mgr0__std__lane20_strm1_data_valid  ),

            .std__mgr0__lane21_strm0_ready           ( std__mgr0__lane21_strm0_ready       ),
            .mgr0__std__lane21_strm0_cntl            ( mgr0__std__lane21_strm0_cntl        ),
            .mgr0__std__lane21_strm0_data            ( mgr0__std__lane21_strm0_data        ),
            .mgr0__std__lane21_strm0_data_valid      ( mgr0__std__lane21_strm0_data_valid  ),

            .std__mgr0__lane21_strm1_ready           ( std__mgr0__lane21_strm1_ready       ),
            .mgr0__std__lane21_strm1_cntl            ( mgr0__std__lane21_strm1_cntl        ),
            .mgr0__std__lane21_strm1_data            ( mgr0__std__lane21_strm1_data        ),
            .mgr0__std__lane21_strm1_data_valid      ( mgr0__std__lane21_strm1_data_valid  ),

            .std__mgr0__lane22_strm0_ready           ( std__mgr0__lane22_strm0_ready       ),
            .mgr0__std__lane22_strm0_cntl            ( mgr0__std__lane22_strm0_cntl        ),
            .mgr0__std__lane22_strm0_data            ( mgr0__std__lane22_strm0_data        ),
            .mgr0__std__lane22_strm0_data_valid      ( mgr0__std__lane22_strm0_data_valid  ),

            .std__mgr0__lane22_strm1_ready           ( std__mgr0__lane22_strm1_ready       ),
            .mgr0__std__lane22_strm1_cntl            ( mgr0__std__lane22_strm1_cntl        ),
            .mgr0__std__lane22_strm1_data            ( mgr0__std__lane22_strm1_data        ),
            .mgr0__std__lane22_strm1_data_valid      ( mgr0__std__lane22_strm1_data_valid  ),

            .std__mgr0__lane23_strm0_ready           ( std__mgr0__lane23_strm0_ready       ),
            .mgr0__std__lane23_strm0_cntl            ( mgr0__std__lane23_strm0_cntl        ),
            .mgr0__std__lane23_strm0_data            ( mgr0__std__lane23_strm0_data        ),
            .mgr0__std__lane23_strm0_data_valid      ( mgr0__std__lane23_strm0_data_valid  ),

            .std__mgr0__lane23_strm1_ready           ( std__mgr0__lane23_strm1_ready       ),
            .mgr0__std__lane23_strm1_cntl            ( mgr0__std__lane23_strm1_cntl        ),
            .mgr0__std__lane23_strm1_data            ( mgr0__std__lane23_strm1_data        ),
            .mgr0__std__lane23_strm1_data_valid      ( mgr0__std__lane23_strm1_data_valid  ),

            .std__mgr0__lane24_strm0_ready           ( std__mgr0__lane24_strm0_ready       ),
            .mgr0__std__lane24_strm0_cntl            ( mgr0__std__lane24_strm0_cntl        ),
            .mgr0__std__lane24_strm0_data            ( mgr0__std__lane24_strm0_data        ),
            .mgr0__std__lane24_strm0_data_valid      ( mgr0__std__lane24_strm0_data_valid  ),

            .std__mgr0__lane24_strm1_ready           ( std__mgr0__lane24_strm1_ready       ),
            .mgr0__std__lane24_strm1_cntl            ( mgr0__std__lane24_strm1_cntl        ),
            .mgr0__std__lane24_strm1_data            ( mgr0__std__lane24_strm1_data        ),
            .mgr0__std__lane24_strm1_data_valid      ( mgr0__std__lane24_strm1_data_valid  ),

            .std__mgr0__lane25_strm0_ready           ( std__mgr0__lane25_strm0_ready       ),
            .mgr0__std__lane25_strm0_cntl            ( mgr0__std__lane25_strm0_cntl        ),
            .mgr0__std__lane25_strm0_data            ( mgr0__std__lane25_strm0_data        ),
            .mgr0__std__lane25_strm0_data_valid      ( mgr0__std__lane25_strm0_data_valid  ),

            .std__mgr0__lane25_strm1_ready           ( std__mgr0__lane25_strm1_ready       ),
            .mgr0__std__lane25_strm1_cntl            ( mgr0__std__lane25_strm1_cntl        ),
            .mgr0__std__lane25_strm1_data            ( mgr0__std__lane25_strm1_data        ),
            .mgr0__std__lane25_strm1_data_valid      ( mgr0__std__lane25_strm1_data_valid  ),

            .std__mgr0__lane26_strm0_ready           ( std__mgr0__lane26_strm0_ready       ),
            .mgr0__std__lane26_strm0_cntl            ( mgr0__std__lane26_strm0_cntl        ),
            .mgr0__std__lane26_strm0_data            ( mgr0__std__lane26_strm0_data        ),
            .mgr0__std__lane26_strm0_data_valid      ( mgr0__std__lane26_strm0_data_valid  ),

            .std__mgr0__lane26_strm1_ready           ( std__mgr0__lane26_strm1_ready       ),
            .mgr0__std__lane26_strm1_cntl            ( mgr0__std__lane26_strm1_cntl        ),
            .mgr0__std__lane26_strm1_data            ( mgr0__std__lane26_strm1_data        ),
            .mgr0__std__lane26_strm1_data_valid      ( mgr0__std__lane26_strm1_data_valid  ),

            .std__mgr0__lane27_strm0_ready           ( std__mgr0__lane27_strm0_ready       ),
            .mgr0__std__lane27_strm0_cntl            ( mgr0__std__lane27_strm0_cntl        ),
            .mgr0__std__lane27_strm0_data            ( mgr0__std__lane27_strm0_data        ),
            .mgr0__std__lane27_strm0_data_valid      ( mgr0__std__lane27_strm0_data_valid  ),

            .std__mgr0__lane27_strm1_ready           ( std__mgr0__lane27_strm1_ready       ),
            .mgr0__std__lane27_strm1_cntl            ( mgr0__std__lane27_strm1_cntl        ),
            .mgr0__std__lane27_strm1_data            ( mgr0__std__lane27_strm1_data        ),
            .mgr0__std__lane27_strm1_data_valid      ( mgr0__std__lane27_strm1_data_valid  ),

            .std__mgr0__lane28_strm0_ready           ( std__mgr0__lane28_strm0_ready       ),
            .mgr0__std__lane28_strm0_cntl            ( mgr0__std__lane28_strm0_cntl        ),
            .mgr0__std__lane28_strm0_data            ( mgr0__std__lane28_strm0_data        ),
            .mgr0__std__lane28_strm0_data_valid      ( mgr0__std__lane28_strm0_data_valid  ),

            .std__mgr0__lane28_strm1_ready           ( std__mgr0__lane28_strm1_ready       ),
            .mgr0__std__lane28_strm1_cntl            ( mgr0__std__lane28_strm1_cntl        ),
            .mgr0__std__lane28_strm1_data            ( mgr0__std__lane28_strm1_data        ),
            .mgr0__std__lane28_strm1_data_valid      ( mgr0__std__lane28_strm1_data_valid  ),

            .std__mgr0__lane29_strm0_ready           ( std__mgr0__lane29_strm0_ready       ),
            .mgr0__std__lane29_strm0_cntl            ( mgr0__std__lane29_strm0_cntl        ),
            .mgr0__std__lane29_strm0_data            ( mgr0__std__lane29_strm0_data        ),
            .mgr0__std__lane29_strm0_data_valid      ( mgr0__std__lane29_strm0_data_valid  ),

            .std__mgr0__lane29_strm1_ready           ( std__mgr0__lane29_strm1_ready       ),
            .mgr0__std__lane29_strm1_cntl            ( mgr0__std__lane29_strm1_cntl        ),
            .mgr0__std__lane29_strm1_data            ( mgr0__std__lane29_strm1_data        ),
            .mgr0__std__lane29_strm1_data_valid      ( mgr0__std__lane29_strm1_data_valid  ),

            .std__mgr0__lane30_strm0_ready           ( std__mgr0__lane30_strm0_ready       ),
            .mgr0__std__lane30_strm0_cntl            ( mgr0__std__lane30_strm0_cntl        ),
            .mgr0__std__lane30_strm0_data            ( mgr0__std__lane30_strm0_data        ),
            .mgr0__std__lane30_strm0_data_valid      ( mgr0__std__lane30_strm0_data_valid  ),

            .std__mgr0__lane30_strm1_ready           ( std__mgr0__lane30_strm1_ready       ),
            .mgr0__std__lane30_strm1_cntl            ( mgr0__std__lane30_strm1_cntl        ),
            .mgr0__std__lane30_strm1_data            ( mgr0__std__lane30_strm1_data        ),
            .mgr0__std__lane30_strm1_data_valid      ( mgr0__std__lane30_strm1_data_valid  ),

            .std__mgr0__lane31_strm0_ready           ( std__mgr0__lane31_strm0_ready       ),
            .mgr0__std__lane31_strm0_cntl            ( mgr0__std__lane31_strm0_cntl        ),
            .mgr0__std__lane31_strm0_data            ( mgr0__std__lane31_strm0_data        ),
            .mgr0__std__lane31_strm0_data_valid      ( mgr0__std__lane31_strm0_data_valid  ),

            .std__mgr0__lane31_strm1_ready           ( std__mgr0__lane31_strm1_ready       ),
            .mgr0__std__lane31_strm1_cntl            ( mgr0__std__lane31_strm1_cntl        ),
            .mgr0__std__lane31_strm1_data            ( mgr0__std__lane31_strm1_data        ),
            .mgr0__std__lane31_strm1_data_valid      ( mgr0__std__lane31_strm1_data_valid  ),

            .std__mgr1__lane0_strm0_ready           ( std__mgr1__lane0_strm0_ready       ),
            .mgr1__std__lane0_strm0_cntl            ( mgr1__std__lane0_strm0_cntl        ),
            .mgr1__std__lane0_strm0_data            ( mgr1__std__lane0_strm0_data        ),
            .mgr1__std__lane0_strm0_data_valid      ( mgr1__std__lane0_strm0_data_valid  ),

            .std__mgr1__lane0_strm1_ready           ( std__mgr1__lane0_strm1_ready       ),
            .mgr1__std__lane0_strm1_cntl            ( mgr1__std__lane0_strm1_cntl        ),
            .mgr1__std__lane0_strm1_data            ( mgr1__std__lane0_strm1_data        ),
            .mgr1__std__lane0_strm1_data_valid      ( mgr1__std__lane0_strm1_data_valid  ),

            .std__mgr1__lane1_strm0_ready           ( std__mgr1__lane1_strm0_ready       ),
            .mgr1__std__lane1_strm0_cntl            ( mgr1__std__lane1_strm0_cntl        ),
            .mgr1__std__lane1_strm0_data            ( mgr1__std__lane1_strm0_data        ),
            .mgr1__std__lane1_strm0_data_valid      ( mgr1__std__lane1_strm0_data_valid  ),

            .std__mgr1__lane1_strm1_ready           ( std__mgr1__lane1_strm1_ready       ),
            .mgr1__std__lane1_strm1_cntl            ( mgr1__std__lane1_strm1_cntl        ),
            .mgr1__std__lane1_strm1_data            ( mgr1__std__lane1_strm1_data        ),
            .mgr1__std__lane1_strm1_data_valid      ( mgr1__std__lane1_strm1_data_valid  ),

            .std__mgr1__lane2_strm0_ready           ( std__mgr1__lane2_strm0_ready       ),
            .mgr1__std__lane2_strm0_cntl            ( mgr1__std__lane2_strm0_cntl        ),
            .mgr1__std__lane2_strm0_data            ( mgr1__std__lane2_strm0_data        ),
            .mgr1__std__lane2_strm0_data_valid      ( mgr1__std__lane2_strm0_data_valid  ),

            .std__mgr1__lane2_strm1_ready           ( std__mgr1__lane2_strm1_ready       ),
            .mgr1__std__lane2_strm1_cntl            ( mgr1__std__lane2_strm1_cntl        ),
            .mgr1__std__lane2_strm1_data            ( mgr1__std__lane2_strm1_data        ),
            .mgr1__std__lane2_strm1_data_valid      ( mgr1__std__lane2_strm1_data_valid  ),

            .std__mgr1__lane3_strm0_ready           ( std__mgr1__lane3_strm0_ready       ),
            .mgr1__std__lane3_strm0_cntl            ( mgr1__std__lane3_strm0_cntl        ),
            .mgr1__std__lane3_strm0_data            ( mgr1__std__lane3_strm0_data        ),
            .mgr1__std__lane3_strm0_data_valid      ( mgr1__std__lane3_strm0_data_valid  ),

            .std__mgr1__lane3_strm1_ready           ( std__mgr1__lane3_strm1_ready       ),
            .mgr1__std__lane3_strm1_cntl            ( mgr1__std__lane3_strm1_cntl        ),
            .mgr1__std__lane3_strm1_data            ( mgr1__std__lane3_strm1_data        ),
            .mgr1__std__lane3_strm1_data_valid      ( mgr1__std__lane3_strm1_data_valid  ),

            .std__mgr1__lane4_strm0_ready           ( std__mgr1__lane4_strm0_ready       ),
            .mgr1__std__lane4_strm0_cntl            ( mgr1__std__lane4_strm0_cntl        ),
            .mgr1__std__lane4_strm0_data            ( mgr1__std__lane4_strm0_data        ),
            .mgr1__std__lane4_strm0_data_valid      ( mgr1__std__lane4_strm0_data_valid  ),

            .std__mgr1__lane4_strm1_ready           ( std__mgr1__lane4_strm1_ready       ),
            .mgr1__std__lane4_strm1_cntl            ( mgr1__std__lane4_strm1_cntl        ),
            .mgr1__std__lane4_strm1_data            ( mgr1__std__lane4_strm1_data        ),
            .mgr1__std__lane4_strm1_data_valid      ( mgr1__std__lane4_strm1_data_valid  ),

            .std__mgr1__lane5_strm0_ready           ( std__mgr1__lane5_strm0_ready       ),
            .mgr1__std__lane5_strm0_cntl            ( mgr1__std__lane5_strm0_cntl        ),
            .mgr1__std__lane5_strm0_data            ( mgr1__std__lane5_strm0_data        ),
            .mgr1__std__lane5_strm0_data_valid      ( mgr1__std__lane5_strm0_data_valid  ),

            .std__mgr1__lane5_strm1_ready           ( std__mgr1__lane5_strm1_ready       ),
            .mgr1__std__lane5_strm1_cntl            ( mgr1__std__lane5_strm1_cntl        ),
            .mgr1__std__lane5_strm1_data            ( mgr1__std__lane5_strm1_data        ),
            .mgr1__std__lane5_strm1_data_valid      ( mgr1__std__lane5_strm1_data_valid  ),

            .std__mgr1__lane6_strm0_ready           ( std__mgr1__lane6_strm0_ready       ),
            .mgr1__std__lane6_strm0_cntl            ( mgr1__std__lane6_strm0_cntl        ),
            .mgr1__std__lane6_strm0_data            ( mgr1__std__lane6_strm0_data        ),
            .mgr1__std__lane6_strm0_data_valid      ( mgr1__std__lane6_strm0_data_valid  ),

            .std__mgr1__lane6_strm1_ready           ( std__mgr1__lane6_strm1_ready       ),
            .mgr1__std__lane6_strm1_cntl            ( mgr1__std__lane6_strm1_cntl        ),
            .mgr1__std__lane6_strm1_data            ( mgr1__std__lane6_strm1_data        ),
            .mgr1__std__lane6_strm1_data_valid      ( mgr1__std__lane6_strm1_data_valid  ),

            .std__mgr1__lane7_strm0_ready           ( std__mgr1__lane7_strm0_ready       ),
            .mgr1__std__lane7_strm0_cntl            ( mgr1__std__lane7_strm0_cntl        ),
            .mgr1__std__lane7_strm0_data            ( mgr1__std__lane7_strm0_data        ),
            .mgr1__std__lane7_strm0_data_valid      ( mgr1__std__lane7_strm0_data_valid  ),

            .std__mgr1__lane7_strm1_ready           ( std__mgr1__lane7_strm1_ready       ),
            .mgr1__std__lane7_strm1_cntl            ( mgr1__std__lane7_strm1_cntl        ),
            .mgr1__std__lane7_strm1_data            ( mgr1__std__lane7_strm1_data        ),
            .mgr1__std__lane7_strm1_data_valid      ( mgr1__std__lane7_strm1_data_valid  ),

            .std__mgr1__lane8_strm0_ready           ( std__mgr1__lane8_strm0_ready       ),
            .mgr1__std__lane8_strm0_cntl            ( mgr1__std__lane8_strm0_cntl        ),
            .mgr1__std__lane8_strm0_data            ( mgr1__std__lane8_strm0_data        ),
            .mgr1__std__lane8_strm0_data_valid      ( mgr1__std__lane8_strm0_data_valid  ),

            .std__mgr1__lane8_strm1_ready           ( std__mgr1__lane8_strm1_ready       ),
            .mgr1__std__lane8_strm1_cntl            ( mgr1__std__lane8_strm1_cntl        ),
            .mgr1__std__lane8_strm1_data            ( mgr1__std__lane8_strm1_data        ),
            .mgr1__std__lane8_strm1_data_valid      ( mgr1__std__lane8_strm1_data_valid  ),

            .std__mgr1__lane9_strm0_ready           ( std__mgr1__lane9_strm0_ready       ),
            .mgr1__std__lane9_strm0_cntl            ( mgr1__std__lane9_strm0_cntl        ),
            .mgr1__std__lane9_strm0_data            ( mgr1__std__lane9_strm0_data        ),
            .mgr1__std__lane9_strm0_data_valid      ( mgr1__std__lane9_strm0_data_valid  ),

            .std__mgr1__lane9_strm1_ready           ( std__mgr1__lane9_strm1_ready       ),
            .mgr1__std__lane9_strm1_cntl            ( mgr1__std__lane9_strm1_cntl        ),
            .mgr1__std__lane9_strm1_data            ( mgr1__std__lane9_strm1_data        ),
            .mgr1__std__lane9_strm1_data_valid      ( mgr1__std__lane9_strm1_data_valid  ),

            .std__mgr1__lane10_strm0_ready           ( std__mgr1__lane10_strm0_ready       ),
            .mgr1__std__lane10_strm0_cntl            ( mgr1__std__lane10_strm0_cntl        ),
            .mgr1__std__lane10_strm0_data            ( mgr1__std__lane10_strm0_data        ),
            .mgr1__std__lane10_strm0_data_valid      ( mgr1__std__lane10_strm0_data_valid  ),

            .std__mgr1__lane10_strm1_ready           ( std__mgr1__lane10_strm1_ready       ),
            .mgr1__std__lane10_strm1_cntl            ( mgr1__std__lane10_strm1_cntl        ),
            .mgr1__std__lane10_strm1_data            ( mgr1__std__lane10_strm1_data        ),
            .mgr1__std__lane10_strm1_data_valid      ( mgr1__std__lane10_strm1_data_valid  ),

            .std__mgr1__lane11_strm0_ready           ( std__mgr1__lane11_strm0_ready       ),
            .mgr1__std__lane11_strm0_cntl            ( mgr1__std__lane11_strm0_cntl        ),
            .mgr1__std__lane11_strm0_data            ( mgr1__std__lane11_strm0_data        ),
            .mgr1__std__lane11_strm0_data_valid      ( mgr1__std__lane11_strm0_data_valid  ),

            .std__mgr1__lane11_strm1_ready           ( std__mgr1__lane11_strm1_ready       ),
            .mgr1__std__lane11_strm1_cntl            ( mgr1__std__lane11_strm1_cntl        ),
            .mgr1__std__lane11_strm1_data            ( mgr1__std__lane11_strm1_data        ),
            .mgr1__std__lane11_strm1_data_valid      ( mgr1__std__lane11_strm1_data_valid  ),

            .std__mgr1__lane12_strm0_ready           ( std__mgr1__lane12_strm0_ready       ),
            .mgr1__std__lane12_strm0_cntl            ( mgr1__std__lane12_strm0_cntl        ),
            .mgr1__std__lane12_strm0_data            ( mgr1__std__lane12_strm0_data        ),
            .mgr1__std__lane12_strm0_data_valid      ( mgr1__std__lane12_strm0_data_valid  ),

            .std__mgr1__lane12_strm1_ready           ( std__mgr1__lane12_strm1_ready       ),
            .mgr1__std__lane12_strm1_cntl            ( mgr1__std__lane12_strm1_cntl        ),
            .mgr1__std__lane12_strm1_data            ( mgr1__std__lane12_strm1_data        ),
            .mgr1__std__lane12_strm1_data_valid      ( mgr1__std__lane12_strm1_data_valid  ),

            .std__mgr1__lane13_strm0_ready           ( std__mgr1__lane13_strm0_ready       ),
            .mgr1__std__lane13_strm0_cntl            ( mgr1__std__lane13_strm0_cntl        ),
            .mgr1__std__lane13_strm0_data            ( mgr1__std__lane13_strm0_data        ),
            .mgr1__std__lane13_strm0_data_valid      ( mgr1__std__lane13_strm0_data_valid  ),

            .std__mgr1__lane13_strm1_ready           ( std__mgr1__lane13_strm1_ready       ),
            .mgr1__std__lane13_strm1_cntl            ( mgr1__std__lane13_strm1_cntl        ),
            .mgr1__std__lane13_strm1_data            ( mgr1__std__lane13_strm1_data        ),
            .mgr1__std__lane13_strm1_data_valid      ( mgr1__std__lane13_strm1_data_valid  ),

            .std__mgr1__lane14_strm0_ready           ( std__mgr1__lane14_strm0_ready       ),
            .mgr1__std__lane14_strm0_cntl            ( mgr1__std__lane14_strm0_cntl        ),
            .mgr1__std__lane14_strm0_data            ( mgr1__std__lane14_strm0_data        ),
            .mgr1__std__lane14_strm0_data_valid      ( mgr1__std__lane14_strm0_data_valid  ),

            .std__mgr1__lane14_strm1_ready           ( std__mgr1__lane14_strm1_ready       ),
            .mgr1__std__lane14_strm1_cntl            ( mgr1__std__lane14_strm1_cntl        ),
            .mgr1__std__lane14_strm1_data            ( mgr1__std__lane14_strm1_data        ),
            .mgr1__std__lane14_strm1_data_valid      ( mgr1__std__lane14_strm1_data_valid  ),

            .std__mgr1__lane15_strm0_ready           ( std__mgr1__lane15_strm0_ready       ),
            .mgr1__std__lane15_strm0_cntl            ( mgr1__std__lane15_strm0_cntl        ),
            .mgr1__std__lane15_strm0_data            ( mgr1__std__lane15_strm0_data        ),
            .mgr1__std__lane15_strm0_data_valid      ( mgr1__std__lane15_strm0_data_valid  ),

            .std__mgr1__lane15_strm1_ready           ( std__mgr1__lane15_strm1_ready       ),
            .mgr1__std__lane15_strm1_cntl            ( mgr1__std__lane15_strm1_cntl        ),
            .mgr1__std__lane15_strm1_data            ( mgr1__std__lane15_strm1_data        ),
            .mgr1__std__lane15_strm1_data_valid      ( mgr1__std__lane15_strm1_data_valid  ),

            .std__mgr1__lane16_strm0_ready           ( std__mgr1__lane16_strm0_ready       ),
            .mgr1__std__lane16_strm0_cntl            ( mgr1__std__lane16_strm0_cntl        ),
            .mgr1__std__lane16_strm0_data            ( mgr1__std__lane16_strm0_data        ),
            .mgr1__std__lane16_strm0_data_valid      ( mgr1__std__lane16_strm0_data_valid  ),

            .std__mgr1__lane16_strm1_ready           ( std__mgr1__lane16_strm1_ready       ),
            .mgr1__std__lane16_strm1_cntl            ( mgr1__std__lane16_strm1_cntl        ),
            .mgr1__std__lane16_strm1_data            ( mgr1__std__lane16_strm1_data        ),
            .mgr1__std__lane16_strm1_data_valid      ( mgr1__std__lane16_strm1_data_valid  ),

            .std__mgr1__lane17_strm0_ready           ( std__mgr1__lane17_strm0_ready       ),
            .mgr1__std__lane17_strm0_cntl            ( mgr1__std__lane17_strm0_cntl        ),
            .mgr1__std__lane17_strm0_data            ( mgr1__std__lane17_strm0_data        ),
            .mgr1__std__lane17_strm0_data_valid      ( mgr1__std__lane17_strm0_data_valid  ),

            .std__mgr1__lane17_strm1_ready           ( std__mgr1__lane17_strm1_ready       ),
            .mgr1__std__lane17_strm1_cntl            ( mgr1__std__lane17_strm1_cntl        ),
            .mgr1__std__lane17_strm1_data            ( mgr1__std__lane17_strm1_data        ),
            .mgr1__std__lane17_strm1_data_valid      ( mgr1__std__lane17_strm1_data_valid  ),

            .std__mgr1__lane18_strm0_ready           ( std__mgr1__lane18_strm0_ready       ),
            .mgr1__std__lane18_strm0_cntl            ( mgr1__std__lane18_strm0_cntl        ),
            .mgr1__std__lane18_strm0_data            ( mgr1__std__lane18_strm0_data        ),
            .mgr1__std__lane18_strm0_data_valid      ( mgr1__std__lane18_strm0_data_valid  ),

            .std__mgr1__lane18_strm1_ready           ( std__mgr1__lane18_strm1_ready       ),
            .mgr1__std__lane18_strm1_cntl            ( mgr1__std__lane18_strm1_cntl        ),
            .mgr1__std__lane18_strm1_data            ( mgr1__std__lane18_strm1_data        ),
            .mgr1__std__lane18_strm1_data_valid      ( mgr1__std__lane18_strm1_data_valid  ),

            .std__mgr1__lane19_strm0_ready           ( std__mgr1__lane19_strm0_ready       ),
            .mgr1__std__lane19_strm0_cntl            ( mgr1__std__lane19_strm0_cntl        ),
            .mgr1__std__lane19_strm0_data            ( mgr1__std__lane19_strm0_data        ),
            .mgr1__std__lane19_strm0_data_valid      ( mgr1__std__lane19_strm0_data_valid  ),

            .std__mgr1__lane19_strm1_ready           ( std__mgr1__lane19_strm1_ready       ),
            .mgr1__std__lane19_strm1_cntl            ( mgr1__std__lane19_strm1_cntl        ),
            .mgr1__std__lane19_strm1_data            ( mgr1__std__lane19_strm1_data        ),
            .mgr1__std__lane19_strm1_data_valid      ( mgr1__std__lane19_strm1_data_valid  ),

            .std__mgr1__lane20_strm0_ready           ( std__mgr1__lane20_strm0_ready       ),
            .mgr1__std__lane20_strm0_cntl            ( mgr1__std__lane20_strm0_cntl        ),
            .mgr1__std__lane20_strm0_data            ( mgr1__std__lane20_strm0_data        ),
            .mgr1__std__lane20_strm0_data_valid      ( mgr1__std__lane20_strm0_data_valid  ),

            .std__mgr1__lane20_strm1_ready           ( std__mgr1__lane20_strm1_ready       ),
            .mgr1__std__lane20_strm1_cntl            ( mgr1__std__lane20_strm1_cntl        ),
            .mgr1__std__lane20_strm1_data            ( mgr1__std__lane20_strm1_data        ),
            .mgr1__std__lane20_strm1_data_valid      ( mgr1__std__lane20_strm1_data_valid  ),

            .std__mgr1__lane21_strm0_ready           ( std__mgr1__lane21_strm0_ready       ),
            .mgr1__std__lane21_strm0_cntl            ( mgr1__std__lane21_strm0_cntl        ),
            .mgr1__std__lane21_strm0_data            ( mgr1__std__lane21_strm0_data        ),
            .mgr1__std__lane21_strm0_data_valid      ( mgr1__std__lane21_strm0_data_valid  ),

            .std__mgr1__lane21_strm1_ready           ( std__mgr1__lane21_strm1_ready       ),
            .mgr1__std__lane21_strm1_cntl            ( mgr1__std__lane21_strm1_cntl        ),
            .mgr1__std__lane21_strm1_data            ( mgr1__std__lane21_strm1_data        ),
            .mgr1__std__lane21_strm1_data_valid      ( mgr1__std__lane21_strm1_data_valid  ),

            .std__mgr1__lane22_strm0_ready           ( std__mgr1__lane22_strm0_ready       ),
            .mgr1__std__lane22_strm0_cntl            ( mgr1__std__lane22_strm0_cntl        ),
            .mgr1__std__lane22_strm0_data            ( mgr1__std__lane22_strm0_data        ),
            .mgr1__std__lane22_strm0_data_valid      ( mgr1__std__lane22_strm0_data_valid  ),

            .std__mgr1__lane22_strm1_ready           ( std__mgr1__lane22_strm1_ready       ),
            .mgr1__std__lane22_strm1_cntl            ( mgr1__std__lane22_strm1_cntl        ),
            .mgr1__std__lane22_strm1_data            ( mgr1__std__lane22_strm1_data        ),
            .mgr1__std__lane22_strm1_data_valid      ( mgr1__std__lane22_strm1_data_valid  ),

            .std__mgr1__lane23_strm0_ready           ( std__mgr1__lane23_strm0_ready       ),
            .mgr1__std__lane23_strm0_cntl            ( mgr1__std__lane23_strm0_cntl        ),
            .mgr1__std__lane23_strm0_data            ( mgr1__std__lane23_strm0_data        ),
            .mgr1__std__lane23_strm0_data_valid      ( mgr1__std__lane23_strm0_data_valid  ),

            .std__mgr1__lane23_strm1_ready           ( std__mgr1__lane23_strm1_ready       ),
            .mgr1__std__lane23_strm1_cntl            ( mgr1__std__lane23_strm1_cntl        ),
            .mgr1__std__lane23_strm1_data            ( mgr1__std__lane23_strm1_data        ),
            .mgr1__std__lane23_strm1_data_valid      ( mgr1__std__lane23_strm1_data_valid  ),

            .std__mgr1__lane24_strm0_ready           ( std__mgr1__lane24_strm0_ready       ),
            .mgr1__std__lane24_strm0_cntl            ( mgr1__std__lane24_strm0_cntl        ),
            .mgr1__std__lane24_strm0_data            ( mgr1__std__lane24_strm0_data        ),
            .mgr1__std__lane24_strm0_data_valid      ( mgr1__std__lane24_strm0_data_valid  ),

            .std__mgr1__lane24_strm1_ready           ( std__mgr1__lane24_strm1_ready       ),
            .mgr1__std__lane24_strm1_cntl            ( mgr1__std__lane24_strm1_cntl        ),
            .mgr1__std__lane24_strm1_data            ( mgr1__std__lane24_strm1_data        ),
            .mgr1__std__lane24_strm1_data_valid      ( mgr1__std__lane24_strm1_data_valid  ),

            .std__mgr1__lane25_strm0_ready           ( std__mgr1__lane25_strm0_ready       ),
            .mgr1__std__lane25_strm0_cntl            ( mgr1__std__lane25_strm0_cntl        ),
            .mgr1__std__lane25_strm0_data            ( mgr1__std__lane25_strm0_data        ),
            .mgr1__std__lane25_strm0_data_valid      ( mgr1__std__lane25_strm0_data_valid  ),

            .std__mgr1__lane25_strm1_ready           ( std__mgr1__lane25_strm1_ready       ),
            .mgr1__std__lane25_strm1_cntl            ( mgr1__std__lane25_strm1_cntl        ),
            .mgr1__std__lane25_strm1_data            ( mgr1__std__lane25_strm1_data        ),
            .mgr1__std__lane25_strm1_data_valid      ( mgr1__std__lane25_strm1_data_valid  ),

            .std__mgr1__lane26_strm0_ready           ( std__mgr1__lane26_strm0_ready       ),
            .mgr1__std__lane26_strm0_cntl            ( mgr1__std__lane26_strm0_cntl        ),
            .mgr1__std__lane26_strm0_data            ( mgr1__std__lane26_strm0_data        ),
            .mgr1__std__lane26_strm0_data_valid      ( mgr1__std__lane26_strm0_data_valid  ),

            .std__mgr1__lane26_strm1_ready           ( std__mgr1__lane26_strm1_ready       ),
            .mgr1__std__lane26_strm1_cntl            ( mgr1__std__lane26_strm1_cntl        ),
            .mgr1__std__lane26_strm1_data            ( mgr1__std__lane26_strm1_data        ),
            .mgr1__std__lane26_strm1_data_valid      ( mgr1__std__lane26_strm1_data_valid  ),

            .std__mgr1__lane27_strm0_ready           ( std__mgr1__lane27_strm0_ready       ),
            .mgr1__std__lane27_strm0_cntl            ( mgr1__std__lane27_strm0_cntl        ),
            .mgr1__std__lane27_strm0_data            ( mgr1__std__lane27_strm0_data        ),
            .mgr1__std__lane27_strm0_data_valid      ( mgr1__std__lane27_strm0_data_valid  ),

            .std__mgr1__lane27_strm1_ready           ( std__mgr1__lane27_strm1_ready       ),
            .mgr1__std__lane27_strm1_cntl            ( mgr1__std__lane27_strm1_cntl        ),
            .mgr1__std__lane27_strm1_data            ( mgr1__std__lane27_strm1_data        ),
            .mgr1__std__lane27_strm1_data_valid      ( mgr1__std__lane27_strm1_data_valid  ),

            .std__mgr1__lane28_strm0_ready           ( std__mgr1__lane28_strm0_ready       ),
            .mgr1__std__lane28_strm0_cntl            ( mgr1__std__lane28_strm0_cntl        ),
            .mgr1__std__lane28_strm0_data            ( mgr1__std__lane28_strm0_data        ),
            .mgr1__std__lane28_strm0_data_valid      ( mgr1__std__lane28_strm0_data_valid  ),

            .std__mgr1__lane28_strm1_ready           ( std__mgr1__lane28_strm1_ready       ),
            .mgr1__std__lane28_strm1_cntl            ( mgr1__std__lane28_strm1_cntl        ),
            .mgr1__std__lane28_strm1_data            ( mgr1__std__lane28_strm1_data        ),
            .mgr1__std__lane28_strm1_data_valid      ( mgr1__std__lane28_strm1_data_valid  ),

            .std__mgr1__lane29_strm0_ready           ( std__mgr1__lane29_strm0_ready       ),
            .mgr1__std__lane29_strm0_cntl            ( mgr1__std__lane29_strm0_cntl        ),
            .mgr1__std__lane29_strm0_data            ( mgr1__std__lane29_strm0_data        ),
            .mgr1__std__lane29_strm0_data_valid      ( mgr1__std__lane29_strm0_data_valid  ),

            .std__mgr1__lane29_strm1_ready           ( std__mgr1__lane29_strm1_ready       ),
            .mgr1__std__lane29_strm1_cntl            ( mgr1__std__lane29_strm1_cntl        ),
            .mgr1__std__lane29_strm1_data            ( mgr1__std__lane29_strm1_data        ),
            .mgr1__std__lane29_strm1_data_valid      ( mgr1__std__lane29_strm1_data_valid  ),

            .std__mgr1__lane30_strm0_ready           ( std__mgr1__lane30_strm0_ready       ),
            .mgr1__std__lane30_strm0_cntl            ( mgr1__std__lane30_strm0_cntl        ),
            .mgr1__std__lane30_strm0_data            ( mgr1__std__lane30_strm0_data        ),
            .mgr1__std__lane30_strm0_data_valid      ( mgr1__std__lane30_strm0_data_valid  ),

            .std__mgr1__lane30_strm1_ready           ( std__mgr1__lane30_strm1_ready       ),
            .mgr1__std__lane30_strm1_cntl            ( mgr1__std__lane30_strm1_cntl        ),
            .mgr1__std__lane30_strm1_data            ( mgr1__std__lane30_strm1_data        ),
            .mgr1__std__lane30_strm1_data_valid      ( mgr1__std__lane30_strm1_data_valid  ),

            .std__mgr1__lane31_strm0_ready           ( std__mgr1__lane31_strm0_ready       ),
            .mgr1__std__lane31_strm0_cntl            ( mgr1__std__lane31_strm0_cntl        ),
            .mgr1__std__lane31_strm0_data            ( mgr1__std__lane31_strm0_data        ),
            .mgr1__std__lane31_strm0_data_valid      ( mgr1__std__lane31_strm0_data_valid  ),

            .std__mgr1__lane31_strm1_ready           ( std__mgr1__lane31_strm1_ready       ),
            .mgr1__std__lane31_strm1_cntl            ( mgr1__std__lane31_strm1_cntl        ),
            .mgr1__std__lane31_strm1_data            ( mgr1__std__lane31_strm1_data        ),
            .mgr1__std__lane31_strm1_data_valid      ( mgr1__std__lane31_strm1_data_valid  ),

            .std__mgr2__lane0_strm0_ready           ( std__mgr2__lane0_strm0_ready       ),
            .mgr2__std__lane0_strm0_cntl            ( mgr2__std__lane0_strm0_cntl        ),
            .mgr2__std__lane0_strm0_data            ( mgr2__std__lane0_strm0_data        ),
            .mgr2__std__lane0_strm0_data_valid      ( mgr2__std__lane0_strm0_data_valid  ),

            .std__mgr2__lane0_strm1_ready           ( std__mgr2__lane0_strm1_ready       ),
            .mgr2__std__lane0_strm1_cntl            ( mgr2__std__lane0_strm1_cntl        ),
            .mgr2__std__lane0_strm1_data            ( mgr2__std__lane0_strm1_data        ),
            .mgr2__std__lane0_strm1_data_valid      ( mgr2__std__lane0_strm1_data_valid  ),

            .std__mgr2__lane1_strm0_ready           ( std__mgr2__lane1_strm0_ready       ),
            .mgr2__std__lane1_strm0_cntl            ( mgr2__std__lane1_strm0_cntl        ),
            .mgr2__std__lane1_strm0_data            ( mgr2__std__lane1_strm0_data        ),
            .mgr2__std__lane1_strm0_data_valid      ( mgr2__std__lane1_strm0_data_valid  ),

            .std__mgr2__lane1_strm1_ready           ( std__mgr2__lane1_strm1_ready       ),
            .mgr2__std__lane1_strm1_cntl            ( mgr2__std__lane1_strm1_cntl        ),
            .mgr2__std__lane1_strm1_data            ( mgr2__std__lane1_strm1_data        ),
            .mgr2__std__lane1_strm1_data_valid      ( mgr2__std__lane1_strm1_data_valid  ),

            .std__mgr2__lane2_strm0_ready           ( std__mgr2__lane2_strm0_ready       ),
            .mgr2__std__lane2_strm0_cntl            ( mgr2__std__lane2_strm0_cntl        ),
            .mgr2__std__lane2_strm0_data            ( mgr2__std__lane2_strm0_data        ),
            .mgr2__std__lane2_strm0_data_valid      ( mgr2__std__lane2_strm0_data_valid  ),

            .std__mgr2__lane2_strm1_ready           ( std__mgr2__lane2_strm1_ready       ),
            .mgr2__std__lane2_strm1_cntl            ( mgr2__std__lane2_strm1_cntl        ),
            .mgr2__std__lane2_strm1_data            ( mgr2__std__lane2_strm1_data        ),
            .mgr2__std__lane2_strm1_data_valid      ( mgr2__std__lane2_strm1_data_valid  ),

            .std__mgr2__lane3_strm0_ready           ( std__mgr2__lane3_strm0_ready       ),
            .mgr2__std__lane3_strm0_cntl            ( mgr2__std__lane3_strm0_cntl        ),
            .mgr2__std__lane3_strm0_data            ( mgr2__std__lane3_strm0_data        ),
            .mgr2__std__lane3_strm0_data_valid      ( mgr2__std__lane3_strm0_data_valid  ),

            .std__mgr2__lane3_strm1_ready           ( std__mgr2__lane3_strm1_ready       ),
            .mgr2__std__lane3_strm1_cntl            ( mgr2__std__lane3_strm1_cntl        ),
            .mgr2__std__lane3_strm1_data            ( mgr2__std__lane3_strm1_data        ),
            .mgr2__std__lane3_strm1_data_valid      ( mgr2__std__lane3_strm1_data_valid  ),

            .std__mgr2__lane4_strm0_ready           ( std__mgr2__lane4_strm0_ready       ),
            .mgr2__std__lane4_strm0_cntl            ( mgr2__std__lane4_strm0_cntl        ),
            .mgr2__std__lane4_strm0_data            ( mgr2__std__lane4_strm0_data        ),
            .mgr2__std__lane4_strm0_data_valid      ( mgr2__std__lane4_strm0_data_valid  ),

            .std__mgr2__lane4_strm1_ready           ( std__mgr2__lane4_strm1_ready       ),
            .mgr2__std__lane4_strm1_cntl            ( mgr2__std__lane4_strm1_cntl        ),
            .mgr2__std__lane4_strm1_data            ( mgr2__std__lane4_strm1_data        ),
            .mgr2__std__lane4_strm1_data_valid      ( mgr2__std__lane4_strm1_data_valid  ),

            .std__mgr2__lane5_strm0_ready           ( std__mgr2__lane5_strm0_ready       ),
            .mgr2__std__lane5_strm0_cntl            ( mgr2__std__lane5_strm0_cntl        ),
            .mgr2__std__lane5_strm0_data            ( mgr2__std__lane5_strm0_data        ),
            .mgr2__std__lane5_strm0_data_valid      ( mgr2__std__lane5_strm0_data_valid  ),

            .std__mgr2__lane5_strm1_ready           ( std__mgr2__lane5_strm1_ready       ),
            .mgr2__std__lane5_strm1_cntl            ( mgr2__std__lane5_strm1_cntl        ),
            .mgr2__std__lane5_strm1_data            ( mgr2__std__lane5_strm1_data        ),
            .mgr2__std__lane5_strm1_data_valid      ( mgr2__std__lane5_strm1_data_valid  ),

            .std__mgr2__lane6_strm0_ready           ( std__mgr2__lane6_strm0_ready       ),
            .mgr2__std__lane6_strm0_cntl            ( mgr2__std__lane6_strm0_cntl        ),
            .mgr2__std__lane6_strm0_data            ( mgr2__std__lane6_strm0_data        ),
            .mgr2__std__lane6_strm0_data_valid      ( mgr2__std__lane6_strm0_data_valid  ),

            .std__mgr2__lane6_strm1_ready           ( std__mgr2__lane6_strm1_ready       ),
            .mgr2__std__lane6_strm1_cntl            ( mgr2__std__lane6_strm1_cntl        ),
            .mgr2__std__lane6_strm1_data            ( mgr2__std__lane6_strm1_data        ),
            .mgr2__std__lane6_strm1_data_valid      ( mgr2__std__lane6_strm1_data_valid  ),

            .std__mgr2__lane7_strm0_ready           ( std__mgr2__lane7_strm0_ready       ),
            .mgr2__std__lane7_strm0_cntl            ( mgr2__std__lane7_strm0_cntl        ),
            .mgr2__std__lane7_strm0_data            ( mgr2__std__lane7_strm0_data        ),
            .mgr2__std__lane7_strm0_data_valid      ( mgr2__std__lane7_strm0_data_valid  ),

            .std__mgr2__lane7_strm1_ready           ( std__mgr2__lane7_strm1_ready       ),
            .mgr2__std__lane7_strm1_cntl            ( mgr2__std__lane7_strm1_cntl        ),
            .mgr2__std__lane7_strm1_data            ( mgr2__std__lane7_strm1_data        ),
            .mgr2__std__lane7_strm1_data_valid      ( mgr2__std__lane7_strm1_data_valid  ),

            .std__mgr2__lane8_strm0_ready           ( std__mgr2__lane8_strm0_ready       ),
            .mgr2__std__lane8_strm0_cntl            ( mgr2__std__lane8_strm0_cntl        ),
            .mgr2__std__lane8_strm0_data            ( mgr2__std__lane8_strm0_data        ),
            .mgr2__std__lane8_strm0_data_valid      ( mgr2__std__lane8_strm0_data_valid  ),

            .std__mgr2__lane8_strm1_ready           ( std__mgr2__lane8_strm1_ready       ),
            .mgr2__std__lane8_strm1_cntl            ( mgr2__std__lane8_strm1_cntl        ),
            .mgr2__std__lane8_strm1_data            ( mgr2__std__lane8_strm1_data        ),
            .mgr2__std__lane8_strm1_data_valid      ( mgr2__std__lane8_strm1_data_valid  ),

            .std__mgr2__lane9_strm0_ready           ( std__mgr2__lane9_strm0_ready       ),
            .mgr2__std__lane9_strm0_cntl            ( mgr2__std__lane9_strm0_cntl        ),
            .mgr2__std__lane9_strm0_data            ( mgr2__std__lane9_strm0_data        ),
            .mgr2__std__lane9_strm0_data_valid      ( mgr2__std__lane9_strm0_data_valid  ),

            .std__mgr2__lane9_strm1_ready           ( std__mgr2__lane9_strm1_ready       ),
            .mgr2__std__lane9_strm1_cntl            ( mgr2__std__lane9_strm1_cntl        ),
            .mgr2__std__lane9_strm1_data            ( mgr2__std__lane9_strm1_data        ),
            .mgr2__std__lane9_strm1_data_valid      ( mgr2__std__lane9_strm1_data_valid  ),

            .std__mgr2__lane10_strm0_ready           ( std__mgr2__lane10_strm0_ready       ),
            .mgr2__std__lane10_strm0_cntl            ( mgr2__std__lane10_strm0_cntl        ),
            .mgr2__std__lane10_strm0_data            ( mgr2__std__lane10_strm0_data        ),
            .mgr2__std__lane10_strm0_data_valid      ( mgr2__std__lane10_strm0_data_valid  ),

            .std__mgr2__lane10_strm1_ready           ( std__mgr2__lane10_strm1_ready       ),
            .mgr2__std__lane10_strm1_cntl            ( mgr2__std__lane10_strm1_cntl        ),
            .mgr2__std__lane10_strm1_data            ( mgr2__std__lane10_strm1_data        ),
            .mgr2__std__lane10_strm1_data_valid      ( mgr2__std__lane10_strm1_data_valid  ),

            .std__mgr2__lane11_strm0_ready           ( std__mgr2__lane11_strm0_ready       ),
            .mgr2__std__lane11_strm0_cntl            ( mgr2__std__lane11_strm0_cntl        ),
            .mgr2__std__lane11_strm0_data            ( mgr2__std__lane11_strm0_data        ),
            .mgr2__std__lane11_strm0_data_valid      ( mgr2__std__lane11_strm0_data_valid  ),

            .std__mgr2__lane11_strm1_ready           ( std__mgr2__lane11_strm1_ready       ),
            .mgr2__std__lane11_strm1_cntl            ( mgr2__std__lane11_strm1_cntl        ),
            .mgr2__std__lane11_strm1_data            ( mgr2__std__lane11_strm1_data        ),
            .mgr2__std__lane11_strm1_data_valid      ( mgr2__std__lane11_strm1_data_valid  ),

            .std__mgr2__lane12_strm0_ready           ( std__mgr2__lane12_strm0_ready       ),
            .mgr2__std__lane12_strm0_cntl            ( mgr2__std__lane12_strm0_cntl        ),
            .mgr2__std__lane12_strm0_data            ( mgr2__std__lane12_strm0_data        ),
            .mgr2__std__lane12_strm0_data_valid      ( mgr2__std__lane12_strm0_data_valid  ),

            .std__mgr2__lane12_strm1_ready           ( std__mgr2__lane12_strm1_ready       ),
            .mgr2__std__lane12_strm1_cntl            ( mgr2__std__lane12_strm1_cntl        ),
            .mgr2__std__lane12_strm1_data            ( mgr2__std__lane12_strm1_data        ),
            .mgr2__std__lane12_strm1_data_valid      ( mgr2__std__lane12_strm1_data_valid  ),

            .std__mgr2__lane13_strm0_ready           ( std__mgr2__lane13_strm0_ready       ),
            .mgr2__std__lane13_strm0_cntl            ( mgr2__std__lane13_strm0_cntl        ),
            .mgr2__std__lane13_strm0_data            ( mgr2__std__lane13_strm0_data        ),
            .mgr2__std__lane13_strm0_data_valid      ( mgr2__std__lane13_strm0_data_valid  ),

            .std__mgr2__lane13_strm1_ready           ( std__mgr2__lane13_strm1_ready       ),
            .mgr2__std__lane13_strm1_cntl            ( mgr2__std__lane13_strm1_cntl        ),
            .mgr2__std__lane13_strm1_data            ( mgr2__std__lane13_strm1_data        ),
            .mgr2__std__lane13_strm1_data_valid      ( mgr2__std__lane13_strm1_data_valid  ),

            .std__mgr2__lane14_strm0_ready           ( std__mgr2__lane14_strm0_ready       ),
            .mgr2__std__lane14_strm0_cntl            ( mgr2__std__lane14_strm0_cntl        ),
            .mgr2__std__lane14_strm0_data            ( mgr2__std__lane14_strm0_data        ),
            .mgr2__std__lane14_strm0_data_valid      ( mgr2__std__lane14_strm0_data_valid  ),

            .std__mgr2__lane14_strm1_ready           ( std__mgr2__lane14_strm1_ready       ),
            .mgr2__std__lane14_strm1_cntl            ( mgr2__std__lane14_strm1_cntl        ),
            .mgr2__std__lane14_strm1_data            ( mgr2__std__lane14_strm1_data        ),
            .mgr2__std__lane14_strm1_data_valid      ( mgr2__std__lane14_strm1_data_valid  ),

            .std__mgr2__lane15_strm0_ready           ( std__mgr2__lane15_strm0_ready       ),
            .mgr2__std__lane15_strm0_cntl            ( mgr2__std__lane15_strm0_cntl        ),
            .mgr2__std__lane15_strm0_data            ( mgr2__std__lane15_strm0_data        ),
            .mgr2__std__lane15_strm0_data_valid      ( mgr2__std__lane15_strm0_data_valid  ),

            .std__mgr2__lane15_strm1_ready           ( std__mgr2__lane15_strm1_ready       ),
            .mgr2__std__lane15_strm1_cntl            ( mgr2__std__lane15_strm1_cntl        ),
            .mgr2__std__lane15_strm1_data            ( mgr2__std__lane15_strm1_data        ),
            .mgr2__std__lane15_strm1_data_valid      ( mgr2__std__lane15_strm1_data_valid  ),

            .std__mgr2__lane16_strm0_ready           ( std__mgr2__lane16_strm0_ready       ),
            .mgr2__std__lane16_strm0_cntl            ( mgr2__std__lane16_strm0_cntl        ),
            .mgr2__std__lane16_strm0_data            ( mgr2__std__lane16_strm0_data        ),
            .mgr2__std__lane16_strm0_data_valid      ( mgr2__std__lane16_strm0_data_valid  ),

            .std__mgr2__lane16_strm1_ready           ( std__mgr2__lane16_strm1_ready       ),
            .mgr2__std__lane16_strm1_cntl            ( mgr2__std__lane16_strm1_cntl        ),
            .mgr2__std__lane16_strm1_data            ( mgr2__std__lane16_strm1_data        ),
            .mgr2__std__lane16_strm1_data_valid      ( mgr2__std__lane16_strm1_data_valid  ),

            .std__mgr2__lane17_strm0_ready           ( std__mgr2__lane17_strm0_ready       ),
            .mgr2__std__lane17_strm0_cntl            ( mgr2__std__lane17_strm0_cntl        ),
            .mgr2__std__lane17_strm0_data            ( mgr2__std__lane17_strm0_data        ),
            .mgr2__std__lane17_strm0_data_valid      ( mgr2__std__lane17_strm0_data_valid  ),

            .std__mgr2__lane17_strm1_ready           ( std__mgr2__lane17_strm1_ready       ),
            .mgr2__std__lane17_strm1_cntl            ( mgr2__std__lane17_strm1_cntl        ),
            .mgr2__std__lane17_strm1_data            ( mgr2__std__lane17_strm1_data        ),
            .mgr2__std__lane17_strm1_data_valid      ( mgr2__std__lane17_strm1_data_valid  ),

            .std__mgr2__lane18_strm0_ready           ( std__mgr2__lane18_strm0_ready       ),
            .mgr2__std__lane18_strm0_cntl            ( mgr2__std__lane18_strm0_cntl        ),
            .mgr2__std__lane18_strm0_data            ( mgr2__std__lane18_strm0_data        ),
            .mgr2__std__lane18_strm0_data_valid      ( mgr2__std__lane18_strm0_data_valid  ),

            .std__mgr2__lane18_strm1_ready           ( std__mgr2__lane18_strm1_ready       ),
            .mgr2__std__lane18_strm1_cntl            ( mgr2__std__lane18_strm1_cntl        ),
            .mgr2__std__lane18_strm1_data            ( mgr2__std__lane18_strm1_data        ),
            .mgr2__std__lane18_strm1_data_valid      ( mgr2__std__lane18_strm1_data_valid  ),

            .std__mgr2__lane19_strm0_ready           ( std__mgr2__lane19_strm0_ready       ),
            .mgr2__std__lane19_strm0_cntl            ( mgr2__std__lane19_strm0_cntl        ),
            .mgr2__std__lane19_strm0_data            ( mgr2__std__lane19_strm0_data        ),
            .mgr2__std__lane19_strm0_data_valid      ( mgr2__std__lane19_strm0_data_valid  ),

            .std__mgr2__lane19_strm1_ready           ( std__mgr2__lane19_strm1_ready       ),
            .mgr2__std__lane19_strm1_cntl            ( mgr2__std__lane19_strm1_cntl        ),
            .mgr2__std__lane19_strm1_data            ( mgr2__std__lane19_strm1_data        ),
            .mgr2__std__lane19_strm1_data_valid      ( mgr2__std__lane19_strm1_data_valid  ),

            .std__mgr2__lane20_strm0_ready           ( std__mgr2__lane20_strm0_ready       ),
            .mgr2__std__lane20_strm0_cntl            ( mgr2__std__lane20_strm0_cntl        ),
            .mgr2__std__lane20_strm0_data            ( mgr2__std__lane20_strm0_data        ),
            .mgr2__std__lane20_strm0_data_valid      ( mgr2__std__lane20_strm0_data_valid  ),

            .std__mgr2__lane20_strm1_ready           ( std__mgr2__lane20_strm1_ready       ),
            .mgr2__std__lane20_strm1_cntl            ( mgr2__std__lane20_strm1_cntl        ),
            .mgr2__std__lane20_strm1_data            ( mgr2__std__lane20_strm1_data        ),
            .mgr2__std__lane20_strm1_data_valid      ( mgr2__std__lane20_strm1_data_valid  ),

            .std__mgr2__lane21_strm0_ready           ( std__mgr2__lane21_strm0_ready       ),
            .mgr2__std__lane21_strm0_cntl            ( mgr2__std__lane21_strm0_cntl        ),
            .mgr2__std__lane21_strm0_data            ( mgr2__std__lane21_strm0_data        ),
            .mgr2__std__lane21_strm0_data_valid      ( mgr2__std__lane21_strm0_data_valid  ),

            .std__mgr2__lane21_strm1_ready           ( std__mgr2__lane21_strm1_ready       ),
            .mgr2__std__lane21_strm1_cntl            ( mgr2__std__lane21_strm1_cntl        ),
            .mgr2__std__lane21_strm1_data            ( mgr2__std__lane21_strm1_data        ),
            .mgr2__std__lane21_strm1_data_valid      ( mgr2__std__lane21_strm1_data_valid  ),

            .std__mgr2__lane22_strm0_ready           ( std__mgr2__lane22_strm0_ready       ),
            .mgr2__std__lane22_strm0_cntl            ( mgr2__std__lane22_strm0_cntl        ),
            .mgr2__std__lane22_strm0_data            ( mgr2__std__lane22_strm0_data        ),
            .mgr2__std__lane22_strm0_data_valid      ( mgr2__std__lane22_strm0_data_valid  ),

            .std__mgr2__lane22_strm1_ready           ( std__mgr2__lane22_strm1_ready       ),
            .mgr2__std__lane22_strm1_cntl            ( mgr2__std__lane22_strm1_cntl        ),
            .mgr2__std__lane22_strm1_data            ( mgr2__std__lane22_strm1_data        ),
            .mgr2__std__lane22_strm1_data_valid      ( mgr2__std__lane22_strm1_data_valid  ),

            .std__mgr2__lane23_strm0_ready           ( std__mgr2__lane23_strm0_ready       ),
            .mgr2__std__lane23_strm0_cntl            ( mgr2__std__lane23_strm0_cntl        ),
            .mgr2__std__lane23_strm0_data            ( mgr2__std__lane23_strm0_data        ),
            .mgr2__std__lane23_strm0_data_valid      ( mgr2__std__lane23_strm0_data_valid  ),

            .std__mgr2__lane23_strm1_ready           ( std__mgr2__lane23_strm1_ready       ),
            .mgr2__std__lane23_strm1_cntl            ( mgr2__std__lane23_strm1_cntl        ),
            .mgr2__std__lane23_strm1_data            ( mgr2__std__lane23_strm1_data        ),
            .mgr2__std__lane23_strm1_data_valid      ( mgr2__std__lane23_strm1_data_valid  ),

            .std__mgr2__lane24_strm0_ready           ( std__mgr2__lane24_strm0_ready       ),
            .mgr2__std__lane24_strm0_cntl            ( mgr2__std__lane24_strm0_cntl        ),
            .mgr2__std__lane24_strm0_data            ( mgr2__std__lane24_strm0_data        ),
            .mgr2__std__lane24_strm0_data_valid      ( mgr2__std__lane24_strm0_data_valid  ),

            .std__mgr2__lane24_strm1_ready           ( std__mgr2__lane24_strm1_ready       ),
            .mgr2__std__lane24_strm1_cntl            ( mgr2__std__lane24_strm1_cntl        ),
            .mgr2__std__lane24_strm1_data            ( mgr2__std__lane24_strm1_data        ),
            .mgr2__std__lane24_strm1_data_valid      ( mgr2__std__lane24_strm1_data_valid  ),

            .std__mgr2__lane25_strm0_ready           ( std__mgr2__lane25_strm0_ready       ),
            .mgr2__std__lane25_strm0_cntl            ( mgr2__std__lane25_strm0_cntl        ),
            .mgr2__std__lane25_strm0_data            ( mgr2__std__lane25_strm0_data        ),
            .mgr2__std__lane25_strm0_data_valid      ( mgr2__std__lane25_strm0_data_valid  ),

            .std__mgr2__lane25_strm1_ready           ( std__mgr2__lane25_strm1_ready       ),
            .mgr2__std__lane25_strm1_cntl            ( mgr2__std__lane25_strm1_cntl        ),
            .mgr2__std__lane25_strm1_data            ( mgr2__std__lane25_strm1_data        ),
            .mgr2__std__lane25_strm1_data_valid      ( mgr2__std__lane25_strm1_data_valid  ),

            .std__mgr2__lane26_strm0_ready           ( std__mgr2__lane26_strm0_ready       ),
            .mgr2__std__lane26_strm0_cntl            ( mgr2__std__lane26_strm0_cntl        ),
            .mgr2__std__lane26_strm0_data            ( mgr2__std__lane26_strm0_data        ),
            .mgr2__std__lane26_strm0_data_valid      ( mgr2__std__lane26_strm0_data_valid  ),

            .std__mgr2__lane26_strm1_ready           ( std__mgr2__lane26_strm1_ready       ),
            .mgr2__std__lane26_strm1_cntl            ( mgr2__std__lane26_strm1_cntl        ),
            .mgr2__std__lane26_strm1_data            ( mgr2__std__lane26_strm1_data        ),
            .mgr2__std__lane26_strm1_data_valid      ( mgr2__std__lane26_strm1_data_valid  ),

            .std__mgr2__lane27_strm0_ready           ( std__mgr2__lane27_strm0_ready       ),
            .mgr2__std__lane27_strm0_cntl            ( mgr2__std__lane27_strm0_cntl        ),
            .mgr2__std__lane27_strm0_data            ( mgr2__std__lane27_strm0_data        ),
            .mgr2__std__lane27_strm0_data_valid      ( mgr2__std__lane27_strm0_data_valid  ),

            .std__mgr2__lane27_strm1_ready           ( std__mgr2__lane27_strm1_ready       ),
            .mgr2__std__lane27_strm1_cntl            ( mgr2__std__lane27_strm1_cntl        ),
            .mgr2__std__lane27_strm1_data            ( mgr2__std__lane27_strm1_data        ),
            .mgr2__std__lane27_strm1_data_valid      ( mgr2__std__lane27_strm1_data_valid  ),

            .std__mgr2__lane28_strm0_ready           ( std__mgr2__lane28_strm0_ready       ),
            .mgr2__std__lane28_strm0_cntl            ( mgr2__std__lane28_strm0_cntl        ),
            .mgr2__std__lane28_strm0_data            ( mgr2__std__lane28_strm0_data        ),
            .mgr2__std__lane28_strm0_data_valid      ( mgr2__std__lane28_strm0_data_valid  ),

            .std__mgr2__lane28_strm1_ready           ( std__mgr2__lane28_strm1_ready       ),
            .mgr2__std__lane28_strm1_cntl            ( mgr2__std__lane28_strm1_cntl        ),
            .mgr2__std__lane28_strm1_data            ( mgr2__std__lane28_strm1_data        ),
            .mgr2__std__lane28_strm1_data_valid      ( mgr2__std__lane28_strm1_data_valid  ),

            .std__mgr2__lane29_strm0_ready           ( std__mgr2__lane29_strm0_ready       ),
            .mgr2__std__lane29_strm0_cntl            ( mgr2__std__lane29_strm0_cntl        ),
            .mgr2__std__lane29_strm0_data            ( mgr2__std__lane29_strm0_data        ),
            .mgr2__std__lane29_strm0_data_valid      ( mgr2__std__lane29_strm0_data_valid  ),

            .std__mgr2__lane29_strm1_ready           ( std__mgr2__lane29_strm1_ready       ),
            .mgr2__std__lane29_strm1_cntl            ( mgr2__std__lane29_strm1_cntl        ),
            .mgr2__std__lane29_strm1_data            ( mgr2__std__lane29_strm1_data        ),
            .mgr2__std__lane29_strm1_data_valid      ( mgr2__std__lane29_strm1_data_valid  ),

            .std__mgr2__lane30_strm0_ready           ( std__mgr2__lane30_strm0_ready       ),
            .mgr2__std__lane30_strm0_cntl            ( mgr2__std__lane30_strm0_cntl        ),
            .mgr2__std__lane30_strm0_data            ( mgr2__std__lane30_strm0_data        ),
            .mgr2__std__lane30_strm0_data_valid      ( mgr2__std__lane30_strm0_data_valid  ),

            .std__mgr2__lane30_strm1_ready           ( std__mgr2__lane30_strm1_ready       ),
            .mgr2__std__lane30_strm1_cntl            ( mgr2__std__lane30_strm1_cntl        ),
            .mgr2__std__lane30_strm1_data            ( mgr2__std__lane30_strm1_data        ),
            .mgr2__std__lane30_strm1_data_valid      ( mgr2__std__lane30_strm1_data_valid  ),

            .std__mgr2__lane31_strm0_ready           ( std__mgr2__lane31_strm0_ready       ),
            .mgr2__std__lane31_strm0_cntl            ( mgr2__std__lane31_strm0_cntl        ),
            .mgr2__std__lane31_strm0_data            ( mgr2__std__lane31_strm0_data        ),
            .mgr2__std__lane31_strm0_data_valid      ( mgr2__std__lane31_strm0_data_valid  ),

            .std__mgr2__lane31_strm1_ready           ( std__mgr2__lane31_strm1_ready       ),
            .mgr2__std__lane31_strm1_cntl            ( mgr2__std__lane31_strm1_cntl        ),
            .mgr2__std__lane31_strm1_data            ( mgr2__std__lane31_strm1_data        ),
            .mgr2__std__lane31_strm1_data_valid      ( mgr2__std__lane31_strm1_data_valid  ),

            .std__mgr3__lane0_strm0_ready           ( std__mgr3__lane0_strm0_ready       ),
            .mgr3__std__lane0_strm0_cntl            ( mgr3__std__lane0_strm0_cntl        ),
            .mgr3__std__lane0_strm0_data            ( mgr3__std__lane0_strm0_data        ),
            .mgr3__std__lane0_strm0_data_valid      ( mgr3__std__lane0_strm0_data_valid  ),

            .std__mgr3__lane0_strm1_ready           ( std__mgr3__lane0_strm1_ready       ),
            .mgr3__std__lane0_strm1_cntl            ( mgr3__std__lane0_strm1_cntl        ),
            .mgr3__std__lane0_strm1_data            ( mgr3__std__lane0_strm1_data        ),
            .mgr3__std__lane0_strm1_data_valid      ( mgr3__std__lane0_strm1_data_valid  ),

            .std__mgr3__lane1_strm0_ready           ( std__mgr3__lane1_strm0_ready       ),
            .mgr3__std__lane1_strm0_cntl            ( mgr3__std__lane1_strm0_cntl        ),
            .mgr3__std__lane1_strm0_data            ( mgr3__std__lane1_strm0_data        ),
            .mgr3__std__lane1_strm0_data_valid      ( mgr3__std__lane1_strm0_data_valid  ),

            .std__mgr3__lane1_strm1_ready           ( std__mgr3__lane1_strm1_ready       ),
            .mgr3__std__lane1_strm1_cntl            ( mgr3__std__lane1_strm1_cntl        ),
            .mgr3__std__lane1_strm1_data            ( mgr3__std__lane1_strm1_data        ),
            .mgr3__std__lane1_strm1_data_valid      ( mgr3__std__lane1_strm1_data_valid  ),

            .std__mgr3__lane2_strm0_ready           ( std__mgr3__lane2_strm0_ready       ),
            .mgr3__std__lane2_strm0_cntl            ( mgr3__std__lane2_strm0_cntl        ),
            .mgr3__std__lane2_strm0_data            ( mgr3__std__lane2_strm0_data        ),
            .mgr3__std__lane2_strm0_data_valid      ( mgr3__std__lane2_strm0_data_valid  ),

            .std__mgr3__lane2_strm1_ready           ( std__mgr3__lane2_strm1_ready       ),
            .mgr3__std__lane2_strm1_cntl            ( mgr3__std__lane2_strm1_cntl        ),
            .mgr3__std__lane2_strm1_data            ( mgr3__std__lane2_strm1_data        ),
            .mgr3__std__lane2_strm1_data_valid      ( mgr3__std__lane2_strm1_data_valid  ),

            .std__mgr3__lane3_strm0_ready           ( std__mgr3__lane3_strm0_ready       ),
            .mgr3__std__lane3_strm0_cntl            ( mgr3__std__lane3_strm0_cntl        ),
            .mgr3__std__lane3_strm0_data            ( mgr3__std__lane3_strm0_data        ),
            .mgr3__std__lane3_strm0_data_valid      ( mgr3__std__lane3_strm0_data_valid  ),

            .std__mgr3__lane3_strm1_ready           ( std__mgr3__lane3_strm1_ready       ),
            .mgr3__std__lane3_strm1_cntl            ( mgr3__std__lane3_strm1_cntl        ),
            .mgr3__std__lane3_strm1_data            ( mgr3__std__lane3_strm1_data        ),
            .mgr3__std__lane3_strm1_data_valid      ( mgr3__std__lane3_strm1_data_valid  ),

            .std__mgr3__lane4_strm0_ready           ( std__mgr3__lane4_strm0_ready       ),
            .mgr3__std__lane4_strm0_cntl            ( mgr3__std__lane4_strm0_cntl        ),
            .mgr3__std__lane4_strm0_data            ( mgr3__std__lane4_strm0_data        ),
            .mgr3__std__lane4_strm0_data_valid      ( mgr3__std__lane4_strm0_data_valid  ),

            .std__mgr3__lane4_strm1_ready           ( std__mgr3__lane4_strm1_ready       ),
            .mgr3__std__lane4_strm1_cntl            ( mgr3__std__lane4_strm1_cntl        ),
            .mgr3__std__lane4_strm1_data            ( mgr3__std__lane4_strm1_data        ),
            .mgr3__std__lane4_strm1_data_valid      ( mgr3__std__lane4_strm1_data_valid  ),

            .std__mgr3__lane5_strm0_ready           ( std__mgr3__lane5_strm0_ready       ),
            .mgr3__std__lane5_strm0_cntl            ( mgr3__std__lane5_strm0_cntl        ),
            .mgr3__std__lane5_strm0_data            ( mgr3__std__lane5_strm0_data        ),
            .mgr3__std__lane5_strm0_data_valid      ( mgr3__std__lane5_strm0_data_valid  ),

            .std__mgr3__lane5_strm1_ready           ( std__mgr3__lane5_strm1_ready       ),
            .mgr3__std__lane5_strm1_cntl            ( mgr3__std__lane5_strm1_cntl        ),
            .mgr3__std__lane5_strm1_data            ( mgr3__std__lane5_strm1_data        ),
            .mgr3__std__lane5_strm1_data_valid      ( mgr3__std__lane5_strm1_data_valid  ),

            .std__mgr3__lane6_strm0_ready           ( std__mgr3__lane6_strm0_ready       ),
            .mgr3__std__lane6_strm0_cntl            ( mgr3__std__lane6_strm0_cntl        ),
            .mgr3__std__lane6_strm0_data            ( mgr3__std__lane6_strm0_data        ),
            .mgr3__std__lane6_strm0_data_valid      ( mgr3__std__lane6_strm0_data_valid  ),

            .std__mgr3__lane6_strm1_ready           ( std__mgr3__lane6_strm1_ready       ),
            .mgr3__std__lane6_strm1_cntl            ( mgr3__std__lane6_strm1_cntl        ),
            .mgr3__std__lane6_strm1_data            ( mgr3__std__lane6_strm1_data        ),
            .mgr3__std__lane6_strm1_data_valid      ( mgr3__std__lane6_strm1_data_valid  ),

            .std__mgr3__lane7_strm0_ready           ( std__mgr3__lane7_strm0_ready       ),
            .mgr3__std__lane7_strm0_cntl            ( mgr3__std__lane7_strm0_cntl        ),
            .mgr3__std__lane7_strm0_data            ( mgr3__std__lane7_strm0_data        ),
            .mgr3__std__lane7_strm0_data_valid      ( mgr3__std__lane7_strm0_data_valid  ),

            .std__mgr3__lane7_strm1_ready           ( std__mgr3__lane7_strm1_ready       ),
            .mgr3__std__lane7_strm1_cntl            ( mgr3__std__lane7_strm1_cntl        ),
            .mgr3__std__lane7_strm1_data            ( mgr3__std__lane7_strm1_data        ),
            .mgr3__std__lane7_strm1_data_valid      ( mgr3__std__lane7_strm1_data_valid  ),

            .std__mgr3__lane8_strm0_ready           ( std__mgr3__lane8_strm0_ready       ),
            .mgr3__std__lane8_strm0_cntl            ( mgr3__std__lane8_strm0_cntl        ),
            .mgr3__std__lane8_strm0_data            ( mgr3__std__lane8_strm0_data        ),
            .mgr3__std__lane8_strm0_data_valid      ( mgr3__std__lane8_strm0_data_valid  ),

            .std__mgr3__lane8_strm1_ready           ( std__mgr3__lane8_strm1_ready       ),
            .mgr3__std__lane8_strm1_cntl            ( mgr3__std__lane8_strm1_cntl        ),
            .mgr3__std__lane8_strm1_data            ( mgr3__std__lane8_strm1_data        ),
            .mgr3__std__lane8_strm1_data_valid      ( mgr3__std__lane8_strm1_data_valid  ),

            .std__mgr3__lane9_strm0_ready           ( std__mgr3__lane9_strm0_ready       ),
            .mgr3__std__lane9_strm0_cntl            ( mgr3__std__lane9_strm0_cntl        ),
            .mgr3__std__lane9_strm0_data            ( mgr3__std__lane9_strm0_data        ),
            .mgr3__std__lane9_strm0_data_valid      ( mgr3__std__lane9_strm0_data_valid  ),

            .std__mgr3__lane9_strm1_ready           ( std__mgr3__lane9_strm1_ready       ),
            .mgr3__std__lane9_strm1_cntl            ( mgr3__std__lane9_strm1_cntl        ),
            .mgr3__std__lane9_strm1_data            ( mgr3__std__lane9_strm1_data        ),
            .mgr3__std__lane9_strm1_data_valid      ( mgr3__std__lane9_strm1_data_valid  ),

            .std__mgr3__lane10_strm0_ready           ( std__mgr3__lane10_strm0_ready       ),
            .mgr3__std__lane10_strm0_cntl            ( mgr3__std__lane10_strm0_cntl        ),
            .mgr3__std__lane10_strm0_data            ( mgr3__std__lane10_strm0_data        ),
            .mgr3__std__lane10_strm0_data_valid      ( mgr3__std__lane10_strm0_data_valid  ),

            .std__mgr3__lane10_strm1_ready           ( std__mgr3__lane10_strm1_ready       ),
            .mgr3__std__lane10_strm1_cntl            ( mgr3__std__lane10_strm1_cntl        ),
            .mgr3__std__lane10_strm1_data            ( mgr3__std__lane10_strm1_data        ),
            .mgr3__std__lane10_strm1_data_valid      ( mgr3__std__lane10_strm1_data_valid  ),

            .std__mgr3__lane11_strm0_ready           ( std__mgr3__lane11_strm0_ready       ),
            .mgr3__std__lane11_strm0_cntl            ( mgr3__std__lane11_strm0_cntl        ),
            .mgr3__std__lane11_strm0_data            ( mgr3__std__lane11_strm0_data        ),
            .mgr3__std__lane11_strm0_data_valid      ( mgr3__std__lane11_strm0_data_valid  ),

            .std__mgr3__lane11_strm1_ready           ( std__mgr3__lane11_strm1_ready       ),
            .mgr3__std__lane11_strm1_cntl            ( mgr3__std__lane11_strm1_cntl        ),
            .mgr3__std__lane11_strm1_data            ( mgr3__std__lane11_strm1_data        ),
            .mgr3__std__lane11_strm1_data_valid      ( mgr3__std__lane11_strm1_data_valid  ),

            .std__mgr3__lane12_strm0_ready           ( std__mgr3__lane12_strm0_ready       ),
            .mgr3__std__lane12_strm0_cntl            ( mgr3__std__lane12_strm0_cntl        ),
            .mgr3__std__lane12_strm0_data            ( mgr3__std__lane12_strm0_data        ),
            .mgr3__std__lane12_strm0_data_valid      ( mgr3__std__lane12_strm0_data_valid  ),

            .std__mgr3__lane12_strm1_ready           ( std__mgr3__lane12_strm1_ready       ),
            .mgr3__std__lane12_strm1_cntl            ( mgr3__std__lane12_strm1_cntl        ),
            .mgr3__std__lane12_strm1_data            ( mgr3__std__lane12_strm1_data        ),
            .mgr3__std__lane12_strm1_data_valid      ( mgr3__std__lane12_strm1_data_valid  ),

            .std__mgr3__lane13_strm0_ready           ( std__mgr3__lane13_strm0_ready       ),
            .mgr3__std__lane13_strm0_cntl            ( mgr3__std__lane13_strm0_cntl        ),
            .mgr3__std__lane13_strm0_data            ( mgr3__std__lane13_strm0_data        ),
            .mgr3__std__lane13_strm0_data_valid      ( mgr3__std__lane13_strm0_data_valid  ),

            .std__mgr3__lane13_strm1_ready           ( std__mgr3__lane13_strm1_ready       ),
            .mgr3__std__lane13_strm1_cntl            ( mgr3__std__lane13_strm1_cntl        ),
            .mgr3__std__lane13_strm1_data            ( mgr3__std__lane13_strm1_data        ),
            .mgr3__std__lane13_strm1_data_valid      ( mgr3__std__lane13_strm1_data_valid  ),

            .std__mgr3__lane14_strm0_ready           ( std__mgr3__lane14_strm0_ready       ),
            .mgr3__std__lane14_strm0_cntl            ( mgr3__std__lane14_strm0_cntl        ),
            .mgr3__std__lane14_strm0_data            ( mgr3__std__lane14_strm0_data        ),
            .mgr3__std__lane14_strm0_data_valid      ( mgr3__std__lane14_strm0_data_valid  ),

            .std__mgr3__lane14_strm1_ready           ( std__mgr3__lane14_strm1_ready       ),
            .mgr3__std__lane14_strm1_cntl            ( mgr3__std__lane14_strm1_cntl        ),
            .mgr3__std__lane14_strm1_data            ( mgr3__std__lane14_strm1_data        ),
            .mgr3__std__lane14_strm1_data_valid      ( mgr3__std__lane14_strm1_data_valid  ),

            .std__mgr3__lane15_strm0_ready           ( std__mgr3__lane15_strm0_ready       ),
            .mgr3__std__lane15_strm0_cntl            ( mgr3__std__lane15_strm0_cntl        ),
            .mgr3__std__lane15_strm0_data            ( mgr3__std__lane15_strm0_data        ),
            .mgr3__std__lane15_strm0_data_valid      ( mgr3__std__lane15_strm0_data_valid  ),

            .std__mgr3__lane15_strm1_ready           ( std__mgr3__lane15_strm1_ready       ),
            .mgr3__std__lane15_strm1_cntl            ( mgr3__std__lane15_strm1_cntl        ),
            .mgr3__std__lane15_strm1_data            ( mgr3__std__lane15_strm1_data        ),
            .mgr3__std__lane15_strm1_data_valid      ( mgr3__std__lane15_strm1_data_valid  ),

            .std__mgr3__lane16_strm0_ready           ( std__mgr3__lane16_strm0_ready       ),
            .mgr3__std__lane16_strm0_cntl            ( mgr3__std__lane16_strm0_cntl        ),
            .mgr3__std__lane16_strm0_data            ( mgr3__std__lane16_strm0_data        ),
            .mgr3__std__lane16_strm0_data_valid      ( mgr3__std__lane16_strm0_data_valid  ),

            .std__mgr3__lane16_strm1_ready           ( std__mgr3__lane16_strm1_ready       ),
            .mgr3__std__lane16_strm1_cntl            ( mgr3__std__lane16_strm1_cntl        ),
            .mgr3__std__lane16_strm1_data            ( mgr3__std__lane16_strm1_data        ),
            .mgr3__std__lane16_strm1_data_valid      ( mgr3__std__lane16_strm1_data_valid  ),

            .std__mgr3__lane17_strm0_ready           ( std__mgr3__lane17_strm0_ready       ),
            .mgr3__std__lane17_strm0_cntl            ( mgr3__std__lane17_strm0_cntl        ),
            .mgr3__std__lane17_strm0_data            ( mgr3__std__lane17_strm0_data        ),
            .mgr3__std__lane17_strm0_data_valid      ( mgr3__std__lane17_strm0_data_valid  ),

            .std__mgr3__lane17_strm1_ready           ( std__mgr3__lane17_strm1_ready       ),
            .mgr3__std__lane17_strm1_cntl            ( mgr3__std__lane17_strm1_cntl        ),
            .mgr3__std__lane17_strm1_data            ( mgr3__std__lane17_strm1_data        ),
            .mgr3__std__lane17_strm1_data_valid      ( mgr3__std__lane17_strm1_data_valid  ),

            .std__mgr3__lane18_strm0_ready           ( std__mgr3__lane18_strm0_ready       ),
            .mgr3__std__lane18_strm0_cntl            ( mgr3__std__lane18_strm0_cntl        ),
            .mgr3__std__lane18_strm0_data            ( mgr3__std__lane18_strm0_data        ),
            .mgr3__std__lane18_strm0_data_valid      ( mgr3__std__lane18_strm0_data_valid  ),

            .std__mgr3__lane18_strm1_ready           ( std__mgr3__lane18_strm1_ready       ),
            .mgr3__std__lane18_strm1_cntl            ( mgr3__std__lane18_strm1_cntl        ),
            .mgr3__std__lane18_strm1_data            ( mgr3__std__lane18_strm1_data        ),
            .mgr3__std__lane18_strm1_data_valid      ( mgr3__std__lane18_strm1_data_valid  ),

            .std__mgr3__lane19_strm0_ready           ( std__mgr3__lane19_strm0_ready       ),
            .mgr3__std__lane19_strm0_cntl            ( mgr3__std__lane19_strm0_cntl        ),
            .mgr3__std__lane19_strm0_data            ( mgr3__std__lane19_strm0_data        ),
            .mgr3__std__lane19_strm0_data_valid      ( mgr3__std__lane19_strm0_data_valid  ),

            .std__mgr3__lane19_strm1_ready           ( std__mgr3__lane19_strm1_ready       ),
            .mgr3__std__lane19_strm1_cntl            ( mgr3__std__lane19_strm1_cntl        ),
            .mgr3__std__lane19_strm1_data            ( mgr3__std__lane19_strm1_data        ),
            .mgr3__std__lane19_strm1_data_valid      ( mgr3__std__lane19_strm1_data_valid  ),

            .std__mgr3__lane20_strm0_ready           ( std__mgr3__lane20_strm0_ready       ),
            .mgr3__std__lane20_strm0_cntl            ( mgr3__std__lane20_strm0_cntl        ),
            .mgr3__std__lane20_strm0_data            ( mgr3__std__lane20_strm0_data        ),
            .mgr3__std__lane20_strm0_data_valid      ( mgr3__std__lane20_strm0_data_valid  ),

            .std__mgr3__lane20_strm1_ready           ( std__mgr3__lane20_strm1_ready       ),
            .mgr3__std__lane20_strm1_cntl            ( mgr3__std__lane20_strm1_cntl        ),
            .mgr3__std__lane20_strm1_data            ( mgr3__std__lane20_strm1_data        ),
            .mgr3__std__lane20_strm1_data_valid      ( mgr3__std__lane20_strm1_data_valid  ),

            .std__mgr3__lane21_strm0_ready           ( std__mgr3__lane21_strm0_ready       ),
            .mgr3__std__lane21_strm0_cntl            ( mgr3__std__lane21_strm0_cntl        ),
            .mgr3__std__lane21_strm0_data            ( mgr3__std__lane21_strm0_data        ),
            .mgr3__std__lane21_strm0_data_valid      ( mgr3__std__lane21_strm0_data_valid  ),

            .std__mgr3__lane21_strm1_ready           ( std__mgr3__lane21_strm1_ready       ),
            .mgr3__std__lane21_strm1_cntl            ( mgr3__std__lane21_strm1_cntl        ),
            .mgr3__std__lane21_strm1_data            ( mgr3__std__lane21_strm1_data        ),
            .mgr3__std__lane21_strm1_data_valid      ( mgr3__std__lane21_strm1_data_valid  ),

            .std__mgr3__lane22_strm0_ready           ( std__mgr3__lane22_strm0_ready       ),
            .mgr3__std__lane22_strm0_cntl            ( mgr3__std__lane22_strm0_cntl        ),
            .mgr3__std__lane22_strm0_data            ( mgr3__std__lane22_strm0_data        ),
            .mgr3__std__lane22_strm0_data_valid      ( mgr3__std__lane22_strm0_data_valid  ),

            .std__mgr3__lane22_strm1_ready           ( std__mgr3__lane22_strm1_ready       ),
            .mgr3__std__lane22_strm1_cntl            ( mgr3__std__lane22_strm1_cntl        ),
            .mgr3__std__lane22_strm1_data            ( mgr3__std__lane22_strm1_data        ),
            .mgr3__std__lane22_strm1_data_valid      ( mgr3__std__lane22_strm1_data_valid  ),

            .std__mgr3__lane23_strm0_ready           ( std__mgr3__lane23_strm0_ready       ),
            .mgr3__std__lane23_strm0_cntl            ( mgr3__std__lane23_strm0_cntl        ),
            .mgr3__std__lane23_strm0_data            ( mgr3__std__lane23_strm0_data        ),
            .mgr3__std__lane23_strm0_data_valid      ( mgr3__std__lane23_strm0_data_valid  ),

            .std__mgr3__lane23_strm1_ready           ( std__mgr3__lane23_strm1_ready       ),
            .mgr3__std__lane23_strm1_cntl            ( mgr3__std__lane23_strm1_cntl        ),
            .mgr3__std__lane23_strm1_data            ( mgr3__std__lane23_strm1_data        ),
            .mgr3__std__lane23_strm1_data_valid      ( mgr3__std__lane23_strm1_data_valid  ),

            .std__mgr3__lane24_strm0_ready           ( std__mgr3__lane24_strm0_ready       ),
            .mgr3__std__lane24_strm0_cntl            ( mgr3__std__lane24_strm0_cntl        ),
            .mgr3__std__lane24_strm0_data            ( mgr3__std__lane24_strm0_data        ),
            .mgr3__std__lane24_strm0_data_valid      ( mgr3__std__lane24_strm0_data_valid  ),

            .std__mgr3__lane24_strm1_ready           ( std__mgr3__lane24_strm1_ready       ),
            .mgr3__std__lane24_strm1_cntl            ( mgr3__std__lane24_strm1_cntl        ),
            .mgr3__std__lane24_strm1_data            ( mgr3__std__lane24_strm1_data        ),
            .mgr3__std__lane24_strm1_data_valid      ( mgr3__std__lane24_strm1_data_valid  ),

            .std__mgr3__lane25_strm0_ready           ( std__mgr3__lane25_strm0_ready       ),
            .mgr3__std__lane25_strm0_cntl            ( mgr3__std__lane25_strm0_cntl        ),
            .mgr3__std__lane25_strm0_data            ( mgr3__std__lane25_strm0_data        ),
            .mgr3__std__lane25_strm0_data_valid      ( mgr3__std__lane25_strm0_data_valid  ),

            .std__mgr3__lane25_strm1_ready           ( std__mgr3__lane25_strm1_ready       ),
            .mgr3__std__lane25_strm1_cntl            ( mgr3__std__lane25_strm1_cntl        ),
            .mgr3__std__lane25_strm1_data            ( mgr3__std__lane25_strm1_data        ),
            .mgr3__std__lane25_strm1_data_valid      ( mgr3__std__lane25_strm1_data_valid  ),

            .std__mgr3__lane26_strm0_ready           ( std__mgr3__lane26_strm0_ready       ),
            .mgr3__std__lane26_strm0_cntl            ( mgr3__std__lane26_strm0_cntl        ),
            .mgr3__std__lane26_strm0_data            ( mgr3__std__lane26_strm0_data        ),
            .mgr3__std__lane26_strm0_data_valid      ( mgr3__std__lane26_strm0_data_valid  ),

            .std__mgr3__lane26_strm1_ready           ( std__mgr3__lane26_strm1_ready       ),
            .mgr3__std__lane26_strm1_cntl            ( mgr3__std__lane26_strm1_cntl        ),
            .mgr3__std__lane26_strm1_data            ( mgr3__std__lane26_strm1_data        ),
            .mgr3__std__lane26_strm1_data_valid      ( mgr3__std__lane26_strm1_data_valid  ),

            .std__mgr3__lane27_strm0_ready           ( std__mgr3__lane27_strm0_ready       ),
            .mgr3__std__lane27_strm0_cntl            ( mgr3__std__lane27_strm0_cntl        ),
            .mgr3__std__lane27_strm0_data            ( mgr3__std__lane27_strm0_data        ),
            .mgr3__std__lane27_strm0_data_valid      ( mgr3__std__lane27_strm0_data_valid  ),

            .std__mgr3__lane27_strm1_ready           ( std__mgr3__lane27_strm1_ready       ),
            .mgr3__std__lane27_strm1_cntl            ( mgr3__std__lane27_strm1_cntl        ),
            .mgr3__std__lane27_strm1_data            ( mgr3__std__lane27_strm1_data        ),
            .mgr3__std__lane27_strm1_data_valid      ( mgr3__std__lane27_strm1_data_valid  ),

            .std__mgr3__lane28_strm0_ready           ( std__mgr3__lane28_strm0_ready       ),
            .mgr3__std__lane28_strm0_cntl            ( mgr3__std__lane28_strm0_cntl        ),
            .mgr3__std__lane28_strm0_data            ( mgr3__std__lane28_strm0_data        ),
            .mgr3__std__lane28_strm0_data_valid      ( mgr3__std__lane28_strm0_data_valid  ),

            .std__mgr3__lane28_strm1_ready           ( std__mgr3__lane28_strm1_ready       ),
            .mgr3__std__lane28_strm1_cntl            ( mgr3__std__lane28_strm1_cntl        ),
            .mgr3__std__lane28_strm1_data            ( mgr3__std__lane28_strm1_data        ),
            .mgr3__std__lane28_strm1_data_valid      ( mgr3__std__lane28_strm1_data_valid  ),

            .std__mgr3__lane29_strm0_ready           ( std__mgr3__lane29_strm0_ready       ),
            .mgr3__std__lane29_strm0_cntl            ( mgr3__std__lane29_strm0_cntl        ),
            .mgr3__std__lane29_strm0_data            ( mgr3__std__lane29_strm0_data        ),
            .mgr3__std__lane29_strm0_data_valid      ( mgr3__std__lane29_strm0_data_valid  ),

            .std__mgr3__lane29_strm1_ready           ( std__mgr3__lane29_strm1_ready       ),
            .mgr3__std__lane29_strm1_cntl            ( mgr3__std__lane29_strm1_cntl        ),
            .mgr3__std__lane29_strm1_data            ( mgr3__std__lane29_strm1_data        ),
            .mgr3__std__lane29_strm1_data_valid      ( mgr3__std__lane29_strm1_data_valid  ),

            .std__mgr3__lane30_strm0_ready           ( std__mgr3__lane30_strm0_ready       ),
            .mgr3__std__lane30_strm0_cntl            ( mgr3__std__lane30_strm0_cntl        ),
            .mgr3__std__lane30_strm0_data            ( mgr3__std__lane30_strm0_data        ),
            .mgr3__std__lane30_strm0_data_valid      ( mgr3__std__lane30_strm0_data_valid  ),

            .std__mgr3__lane30_strm1_ready           ( std__mgr3__lane30_strm1_ready       ),
            .mgr3__std__lane30_strm1_cntl            ( mgr3__std__lane30_strm1_cntl        ),
            .mgr3__std__lane30_strm1_data            ( mgr3__std__lane30_strm1_data        ),
            .mgr3__std__lane30_strm1_data_valid      ( mgr3__std__lane30_strm1_data_valid  ),

            .std__mgr3__lane31_strm0_ready           ( std__mgr3__lane31_strm0_ready       ),
            .mgr3__std__lane31_strm0_cntl            ( mgr3__std__lane31_strm0_cntl        ),
            .mgr3__std__lane31_strm0_data            ( mgr3__std__lane31_strm0_data        ),
            .mgr3__std__lane31_strm0_data_valid      ( mgr3__std__lane31_strm0_data_valid  ),

            .std__mgr3__lane31_strm1_ready           ( std__mgr3__lane31_strm1_ready       ),
            .mgr3__std__lane31_strm1_cntl            ( mgr3__std__lane31_strm1_cntl        ),
            .mgr3__std__lane31_strm1_data            ( mgr3__std__lane31_strm1_data        ),
            .mgr3__std__lane31_strm1_data_valid      ( mgr3__std__lane31_strm1_data_valid  ),
