
            begin
              ldst_driver[0].run()  ;
            end
            begin
              mgr[0].run()  ;
            end
            begin
              oob_drv[0].run()  ;
            end
            begin
              up_check[0].run()  ;
            end
            begin
              gen[0][0].run()  ;
            end
            begin
              drv[0][0].run()  ;
            end
            begin
              mem_check[0][0].run()  ;
            end
            begin
              rf_driver[0][0].run()  ;
            end

            begin
              gen[0][1].run()  ;
            end
            begin
              drv[0][1].run()  ;
            end
            begin
              mem_check[0][1].run()  ;
            end
            begin
              rf_driver[0][1].run()  ;
            end

            begin
              gen[0][2].run()  ;
            end
            begin
              drv[0][2].run()  ;
            end
            begin
              mem_check[0][2].run()  ;
            end
            begin
              rf_driver[0][2].run()  ;
            end

            begin
              gen[0][3].run()  ;
            end
            begin
              drv[0][3].run()  ;
            end
            begin
              mem_check[0][3].run()  ;
            end
            begin
              rf_driver[0][3].run()  ;
            end

            begin
              gen[0][4].run()  ;
            end
            begin
              drv[0][4].run()  ;
            end
            begin
              mem_check[0][4].run()  ;
            end
            begin
              rf_driver[0][4].run()  ;
            end

            begin
              gen[0][5].run()  ;
            end
            begin
              drv[0][5].run()  ;
            end
            begin
              mem_check[0][5].run()  ;
            end
            begin
              rf_driver[0][5].run()  ;
            end

            begin
              gen[0][6].run()  ;
            end
            begin
              drv[0][6].run()  ;
            end
            begin
              mem_check[0][6].run()  ;
            end
            begin
              rf_driver[0][6].run()  ;
            end

            begin
              gen[0][7].run()  ;
            end
            begin
              drv[0][7].run()  ;
            end
            begin
              mem_check[0][7].run()  ;
            end
            begin
              rf_driver[0][7].run()  ;
            end

            begin
              gen[0][8].run()  ;
            end
            begin
              drv[0][8].run()  ;
            end
            begin
              mem_check[0][8].run()  ;
            end
            begin
              rf_driver[0][8].run()  ;
            end

            begin
              gen[0][9].run()  ;
            end
            begin
              drv[0][9].run()  ;
            end
            begin
              mem_check[0][9].run()  ;
            end
            begin
              rf_driver[0][9].run()  ;
            end

            begin
              gen[0][10].run()  ;
            end
            begin
              drv[0][10].run()  ;
            end
            begin
              mem_check[0][10].run()  ;
            end
            begin
              rf_driver[0][10].run()  ;
            end

            begin
              gen[0][11].run()  ;
            end
            begin
              drv[0][11].run()  ;
            end
            begin
              mem_check[0][11].run()  ;
            end
            begin
              rf_driver[0][11].run()  ;
            end

            begin
              gen[0][12].run()  ;
            end
            begin
              drv[0][12].run()  ;
            end
            begin
              mem_check[0][12].run()  ;
            end
            begin
              rf_driver[0][12].run()  ;
            end

            begin
              gen[0][13].run()  ;
            end
            begin
              drv[0][13].run()  ;
            end
            begin
              mem_check[0][13].run()  ;
            end
            begin
              rf_driver[0][13].run()  ;
            end

            begin
              gen[0][14].run()  ;
            end
            begin
              drv[0][14].run()  ;
            end
            begin
              mem_check[0][14].run()  ;
            end
            begin
              rf_driver[0][14].run()  ;
            end

            begin
              gen[0][15].run()  ;
            end
            begin
              drv[0][15].run()  ;
            end
            begin
              mem_check[0][15].run()  ;
            end
            begin
              rf_driver[0][15].run()  ;
            end

            begin
              gen[0][16].run()  ;
            end
            begin
              drv[0][16].run()  ;
            end
            begin
              mem_check[0][16].run()  ;
            end
            begin
              rf_driver[0][16].run()  ;
            end

            begin
              gen[0][17].run()  ;
            end
            begin
              drv[0][17].run()  ;
            end
            begin
              mem_check[0][17].run()  ;
            end
            begin
              rf_driver[0][17].run()  ;
            end

            begin
              gen[0][18].run()  ;
            end
            begin
              drv[0][18].run()  ;
            end
            begin
              mem_check[0][18].run()  ;
            end
            begin
              rf_driver[0][18].run()  ;
            end

            begin
              gen[0][19].run()  ;
            end
            begin
              drv[0][19].run()  ;
            end
            begin
              mem_check[0][19].run()  ;
            end
            begin
              rf_driver[0][19].run()  ;
            end

            begin
              gen[0][20].run()  ;
            end
            begin
              drv[0][20].run()  ;
            end
            begin
              mem_check[0][20].run()  ;
            end
            begin
              rf_driver[0][20].run()  ;
            end

            begin
              gen[0][21].run()  ;
            end
            begin
              drv[0][21].run()  ;
            end
            begin
              mem_check[0][21].run()  ;
            end
            begin
              rf_driver[0][21].run()  ;
            end

            begin
              gen[0][22].run()  ;
            end
            begin
              drv[0][22].run()  ;
            end
            begin
              mem_check[0][22].run()  ;
            end
            begin
              rf_driver[0][22].run()  ;
            end

            begin
              gen[0][23].run()  ;
            end
            begin
              drv[0][23].run()  ;
            end
            begin
              mem_check[0][23].run()  ;
            end
            begin
              rf_driver[0][23].run()  ;
            end

            begin
              gen[0][24].run()  ;
            end
            begin
              drv[0][24].run()  ;
            end
            begin
              mem_check[0][24].run()  ;
            end
            begin
              rf_driver[0][24].run()  ;
            end

            begin
              gen[0][25].run()  ;
            end
            begin
              drv[0][25].run()  ;
            end
            begin
              mem_check[0][25].run()  ;
            end
            begin
              rf_driver[0][25].run()  ;
            end

            begin
              gen[0][26].run()  ;
            end
            begin
              drv[0][26].run()  ;
            end
            begin
              mem_check[0][26].run()  ;
            end
            begin
              rf_driver[0][26].run()  ;
            end

            begin
              gen[0][27].run()  ;
            end
            begin
              drv[0][27].run()  ;
            end
            begin
              mem_check[0][27].run()  ;
            end
            begin
              rf_driver[0][27].run()  ;
            end

            begin
              gen[0][28].run()  ;
            end
            begin
              drv[0][28].run()  ;
            end
            begin
              mem_check[0][28].run()  ;
            end
            begin
              rf_driver[0][28].run()  ;
            end

            begin
              gen[0][29].run()  ;
            end
            begin
              drv[0][29].run()  ;
            end
            begin
              mem_check[0][29].run()  ;
            end
            begin
              rf_driver[0][29].run()  ;
            end

            begin
              gen[0][30].run()  ;
            end
            begin
              drv[0][30].run()  ;
            end
            begin
              mem_check[0][30].run()  ;
            end
            begin
              rf_driver[0][30].run()  ;
            end

            begin
              gen[0][31].run()  ;
            end
            begin
              drv[0][31].run()  ;
            end
            begin
              mem_check[0][31].run()  ;
            end
            begin
              rf_driver[0][31].run()  ;
            end

            begin
              ldst_driver[1].run()  ;
            end
            begin
              mgr[1].run()  ;
            end
            begin
              oob_drv[1].run()  ;
            end
            begin
              up_check[1].run()  ;
            end
            begin
              gen[1][0].run()  ;
            end
            begin
              drv[1][0].run()  ;
            end
            begin
              mem_check[1][0].run()  ;
            end
            begin
              rf_driver[1][0].run()  ;
            end

            begin
              gen[1][1].run()  ;
            end
            begin
              drv[1][1].run()  ;
            end
            begin
              mem_check[1][1].run()  ;
            end
            begin
              rf_driver[1][1].run()  ;
            end

            begin
              gen[1][2].run()  ;
            end
            begin
              drv[1][2].run()  ;
            end
            begin
              mem_check[1][2].run()  ;
            end
            begin
              rf_driver[1][2].run()  ;
            end

            begin
              gen[1][3].run()  ;
            end
            begin
              drv[1][3].run()  ;
            end
            begin
              mem_check[1][3].run()  ;
            end
            begin
              rf_driver[1][3].run()  ;
            end

            begin
              gen[1][4].run()  ;
            end
            begin
              drv[1][4].run()  ;
            end
            begin
              mem_check[1][4].run()  ;
            end
            begin
              rf_driver[1][4].run()  ;
            end

            begin
              gen[1][5].run()  ;
            end
            begin
              drv[1][5].run()  ;
            end
            begin
              mem_check[1][5].run()  ;
            end
            begin
              rf_driver[1][5].run()  ;
            end

            begin
              gen[1][6].run()  ;
            end
            begin
              drv[1][6].run()  ;
            end
            begin
              mem_check[1][6].run()  ;
            end
            begin
              rf_driver[1][6].run()  ;
            end

            begin
              gen[1][7].run()  ;
            end
            begin
              drv[1][7].run()  ;
            end
            begin
              mem_check[1][7].run()  ;
            end
            begin
              rf_driver[1][7].run()  ;
            end

            begin
              gen[1][8].run()  ;
            end
            begin
              drv[1][8].run()  ;
            end
            begin
              mem_check[1][8].run()  ;
            end
            begin
              rf_driver[1][8].run()  ;
            end

            begin
              gen[1][9].run()  ;
            end
            begin
              drv[1][9].run()  ;
            end
            begin
              mem_check[1][9].run()  ;
            end
            begin
              rf_driver[1][9].run()  ;
            end

            begin
              gen[1][10].run()  ;
            end
            begin
              drv[1][10].run()  ;
            end
            begin
              mem_check[1][10].run()  ;
            end
            begin
              rf_driver[1][10].run()  ;
            end

            begin
              gen[1][11].run()  ;
            end
            begin
              drv[1][11].run()  ;
            end
            begin
              mem_check[1][11].run()  ;
            end
            begin
              rf_driver[1][11].run()  ;
            end

            begin
              gen[1][12].run()  ;
            end
            begin
              drv[1][12].run()  ;
            end
            begin
              mem_check[1][12].run()  ;
            end
            begin
              rf_driver[1][12].run()  ;
            end

            begin
              gen[1][13].run()  ;
            end
            begin
              drv[1][13].run()  ;
            end
            begin
              mem_check[1][13].run()  ;
            end
            begin
              rf_driver[1][13].run()  ;
            end

            begin
              gen[1][14].run()  ;
            end
            begin
              drv[1][14].run()  ;
            end
            begin
              mem_check[1][14].run()  ;
            end
            begin
              rf_driver[1][14].run()  ;
            end

            begin
              gen[1][15].run()  ;
            end
            begin
              drv[1][15].run()  ;
            end
            begin
              mem_check[1][15].run()  ;
            end
            begin
              rf_driver[1][15].run()  ;
            end

            begin
              gen[1][16].run()  ;
            end
            begin
              drv[1][16].run()  ;
            end
            begin
              mem_check[1][16].run()  ;
            end
            begin
              rf_driver[1][16].run()  ;
            end

            begin
              gen[1][17].run()  ;
            end
            begin
              drv[1][17].run()  ;
            end
            begin
              mem_check[1][17].run()  ;
            end
            begin
              rf_driver[1][17].run()  ;
            end

            begin
              gen[1][18].run()  ;
            end
            begin
              drv[1][18].run()  ;
            end
            begin
              mem_check[1][18].run()  ;
            end
            begin
              rf_driver[1][18].run()  ;
            end

            begin
              gen[1][19].run()  ;
            end
            begin
              drv[1][19].run()  ;
            end
            begin
              mem_check[1][19].run()  ;
            end
            begin
              rf_driver[1][19].run()  ;
            end

            begin
              gen[1][20].run()  ;
            end
            begin
              drv[1][20].run()  ;
            end
            begin
              mem_check[1][20].run()  ;
            end
            begin
              rf_driver[1][20].run()  ;
            end

            begin
              gen[1][21].run()  ;
            end
            begin
              drv[1][21].run()  ;
            end
            begin
              mem_check[1][21].run()  ;
            end
            begin
              rf_driver[1][21].run()  ;
            end

            begin
              gen[1][22].run()  ;
            end
            begin
              drv[1][22].run()  ;
            end
            begin
              mem_check[1][22].run()  ;
            end
            begin
              rf_driver[1][22].run()  ;
            end

            begin
              gen[1][23].run()  ;
            end
            begin
              drv[1][23].run()  ;
            end
            begin
              mem_check[1][23].run()  ;
            end
            begin
              rf_driver[1][23].run()  ;
            end

            begin
              gen[1][24].run()  ;
            end
            begin
              drv[1][24].run()  ;
            end
            begin
              mem_check[1][24].run()  ;
            end
            begin
              rf_driver[1][24].run()  ;
            end

            begin
              gen[1][25].run()  ;
            end
            begin
              drv[1][25].run()  ;
            end
            begin
              mem_check[1][25].run()  ;
            end
            begin
              rf_driver[1][25].run()  ;
            end

            begin
              gen[1][26].run()  ;
            end
            begin
              drv[1][26].run()  ;
            end
            begin
              mem_check[1][26].run()  ;
            end
            begin
              rf_driver[1][26].run()  ;
            end

            begin
              gen[1][27].run()  ;
            end
            begin
              drv[1][27].run()  ;
            end
            begin
              mem_check[1][27].run()  ;
            end
            begin
              rf_driver[1][27].run()  ;
            end

            begin
              gen[1][28].run()  ;
            end
            begin
              drv[1][28].run()  ;
            end
            begin
              mem_check[1][28].run()  ;
            end
            begin
              rf_driver[1][28].run()  ;
            end

            begin
              gen[1][29].run()  ;
            end
            begin
              drv[1][29].run()  ;
            end
            begin
              mem_check[1][29].run()  ;
            end
            begin
              rf_driver[1][29].run()  ;
            end

            begin
              gen[1][30].run()  ;
            end
            begin
              drv[1][30].run()  ;
            end
            begin
              mem_check[1][30].run()  ;
            end
            begin
              rf_driver[1][30].run()  ;
            end

            begin
              gen[1][31].run()  ;
            end
            begin
              drv[1][31].run()  ;
            end
            begin
              mem_check[1][31].run()  ;
            end
            begin
              rf_driver[1][31].run()  ;
            end

            begin
              ldst_driver[2].run()  ;
            end
            begin
              mgr[2].run()  ;
            end
            begin
              oob_drv[2].run()  ;
            end
            begin
              up_check[2].run()  ;
            end
            begin
              gen[2][0].run()  ;
            end
            begin
              drv[2][0].run()  ;
            end
            begin
              mem_check[2][0].run()  ;
            end
            begin
              rf_driver[2][0].run()  ;
            end

            begin
              gen[2][1].run()  ;
            end
            begin
              drv[2][1].run()  ;
            end
            begin
              mem_check[2][1].run()  ;
            end
            begin
              rf_driver[2][1].run()  ;
            end

            begin
              gen[2][2].run()  ;
            end
            begin
              drv[2][2].run()  ;
            end
            begin
              mem_check[2][2].run()  ;
            end
            begin
              rf_driver[2][2].run()  ;
            end

            begin
              gen[2][3].run()  ;
            end
            begin
              drv[2][3].run()  ;
            end
            begin
              mem_check[2][3].run()  ;
            end
            begin
              rf_driver[2][3].run()  ;
            end

            begin
              gen[2][4].run()  ;
            end
            begin
              drv[2][4].run()  ;
            end
            begin
              mem_check[2][4].run()  ;
            end
            begin
              rf_driver[2][4].run()  ;
            end

            begin
              gen[2][5].run()  ;
            end
            begin
              drv[2][5].run()  ;
            end
            begin
              mem_check[2][5].run()  ;
            end
            begin
              rf_driver[2][5].run()  ;
            end

            begin
              gen[2][6].run()  ;
            end
            begin
              drv[2][6].run()  ;
            end
            begin
              mem_check[2][6].run()  ;
            end
            begin
              rf_driver[2][6].run()  ;
            end

            begin
              gen[2][7].run()  ;
            end
            begin
              drv[2][7].run()  ;
            end
            begin
              mem_check[2][7].run()  ;
            end
            begin
              rf_driver[2][7].run()  ;
            end

            begin
              gen[2][8].run()  ;
            end
            begin
              drv[2][8].run()  ;
            end
            begin
              mem_check[2][8].run()  ;
            end
            begin
              rf_driver[2][8].run()  ;
            end

            begin
              gen[2][9].run()  ;
            end
            begin
              drv[2][9].run()  ;
            end
            begin
              mem_check[2][9].run()  ;
            end
            begin
              rf_driver[2][9].run()  ;
            end

            begin
              gen[2][10].run()  ;
            end
            begin
              drv[2][10].run()  ;
            end
            begin
              mem_check[2][10].run()  ;
            end
            begin
              rf_driver[2][10].run()  ;
            end

            begin
              gen[2][11].run()  ;
            end
            begin
              drv[2][11].run()  ;
            end
            begin
              mem_check[2][11].run()  ;
            end
            begin
              rf_driver[2][11].run()  ;
            end

            begin
              gen[2][12].run()  ;
            end
            begin
              drv[2][12].run()  ;
            end
            begin
              mem_check[2][12].run()  ;
            end
            begin
              rf_driver[2][12].run()  ;
            end

            begin
              gen[2][13].run()  ;
            end
            begin
              drv[2][13].run()  ;
            end
            begin
              mem_check[2][13].run()  ;
            end
            begin
              rf_driver[2][13].run()  ;
            end

            begin
              gen[2][14].run()  ;
            end
            begin
              drv[2][14].run()  ;
            end
            begin
              mem_check[2][14].run()  ;
            end
            begin
              rf_driver[2][14].run()  ;
            end

            begin
              gen[2][15].run()  ;
            end
            begin
              drv[2][15].run()  ;
            end
            begin
              mem_check[2][15].run()  ;
            end
            begin
              rf_driver[2][15].run()  ;
            end

            begin
              gen[2][16].run()  ;
            end
            begin
              drv[2][16].run()  ;
            end
            begin
              mem_check[2][16].run()  ;
            end
            begin
              rf_driver[2][16].run()  ;
            end

            begin
              gen[2][17].run()  ;
            end
            begin
              drv[2][17].run()  ;
            end
            begin
              mem_check[2][17].run()  ;
            end
            begin
              rf_driver[2][17].run()  ;
            end

            begin
              gen[2][18].run()  ;
            end
            begin
              drv[2][18].run()  ;
            end
            begin
              mem_check[2][18].run()  ;
            end
            begin
              rf_driver[2][18].run()  ;
            end

            begin
              gen[2][19].run()  ;
            end
            begin
              drv[2][19].run()  ;
            end
            begin
              mem_check[2][19].run()  ;
            end
            begin
              rf_driver[2][19].run()  ;
            end

            begin
              gen[2][20].run()  ;
            end
            begin
              drv[2][20].run()  ;
            end
            begin
              mem_check[2][20].run()  ;
            end
            begin
              rf_driver[2][20].run()  ;
            end

            begin
              gen[2][21].run()  ;
            end
            begin
              drv[2][21].run()  ;
            end
            begin
              mem_check[2][21].run()  ;
            end
            begin
              rf_driver[2][21].run()  ;
            end

            begin
              gen[2][22].run()  ;
            end
            begin
              drv[2][22].run()  ;
            end
            begin
              mem_check[2][22].run()  ;
            end
            begin
              rf_driver[2][22].run()  ;
            end

            begin
              gen[2][23].run()  ;
            end
            begin
              drv[2][23].run()  ;
            end
            begin
              mem_check[2][23].run()  ;
            end
            begin
              rf_driver[2][23].run()  ;
            end

            begin
              gen[2][24].run()  ;
            end
            begin
              drv[2][24].run()  ;
            end
            begin
              mem_check[2][24].run()  ;
            end
            begin
              rf_driver[2][24].run()  ;
            end

            begin
              gen[2][25].run()  ;
            end
            begin
              drv[2][25].run()  ;
            end
            begin
              mem_check[2][25].run()  ;
            end
            begin
              rf_driver[2][25].run()  ;
            end

            begin
              gen[2][26].run()  ;
            end
            begin
              drv[2][26].run()  ;
            end
            begin
              mem_check[2][26].run()  ;
            end
            begin
              rf_driver[2][26].run()  ;
            end

            begin
              gen[2][27].run()  ;
            end
            begin
              drv[2][27].run()  ;
            end
            begin
              mem_check[2][27].run()  ;
            end
            begin
              rf_driver[2][27].run()  ;
            end

            begin
              gen[2][28].run()  ;
            end
            begin
              drv[2][28].run()  ;
            end
            begin
              mem_check[2][28].run()  ;
            end
            begin
              rf_driver[2][28].run()  ;
            end

            begin
              gen[2][29].run()  ;
            end
            begin
              drv[2][29].run()  ;
            end
            begin
              mem_check[2][29].run()  ;
            end
            begin
              rf_driver[2][29].run()  ;
            end

            begin
              gen[2][30].run()  ;
            end
            begin
              drv[2][30].run()  ;
            end
            begin
              mem_check[2][30].run()  ;
            end
            begin
              rf_driver[2][30].run()  ;
            end

            begin
              gen[2][31].run()  ;
            end
            begin
              drv[2][31].run()  ;
            end
            begin
              mem_check[2][31].run()  ;
            end
            begin
              rf_driver[2][31].run()  ;
            end

            begin
              ldst_driver[3].run()  ;
            end
            begin
              mgr[3].run()  ;
            end
            begin
              oob_drv[3].run()  ;
            end
            begin
              up_check[3].run()  ;
            end
            begin
              gen[3][0].run()  ;
            end
            begin
              drv[3][0].run()  ;
            end
            begin
              mem_check[3][0].run()  ;
            end
            begin
              rf_driver[3][0].run()  ;
            end

            begin
              gen[3][1].run()  ;
            end
            begin
              drv[3][1].run()  ;
            end
            begin
              mem_check[3][1].run()  ;
            end
            begin
              rf_driver[3][1].run()  ;
            end

            begin
              gen[3][2].run()  ;
            end
            begin
              drv[3][2].run()  ;
            end
            begin
              mem_check[3][2].run()  ;
            end
            begin
              rf_driver[3][2].run()  ;
            end

            begin
              gen[3][3].run()  ;
            end
            begin
              drv[3][3].run()  ;
            end
            begin
              mem_check[3][3].run()  ;
            end
            begin
              rf_driver[3][3].run()  ;
            end

            begin
              gen[3][4].run()  ;
            end
            begin
              drv[3][4].run()  ;
            end
            begin
              mem_check[3][4].run()  ;
            end
            begin
              rf_driver[3][4].run()  ;
            end

            begin
              gen[3][5].run()  ;
            end
            begin
              drv[3][5].run()  ;
            end
            begin
              mem_check[3][5].run()  ;
            end
            begin
              rf_driver[3][5].run()  ;
            end

            begin
              gen[3][6].run()  ;
            end
            begin
              drv[3][6].run()  ;
            end
            begin
              mem_check[3][6].run()  ;
            end
            begin
              rf_driver[3][6].run()  ;
            end

            begin
              gen[3][7].run()  ;
            end
            begin
              drv[3][7].run()  ;
            end
            begin
              mem_check[3][7].run()  ;
            end
            begin
              rf_driver[3][7].run()  ;
            end

            begin
              gen[3][8].run()  ;
            end
            begin
              drv[3][8].run()  ;
            end
            begin
              mem_check[3][8].run()  ;
            end
            begin
              rf_driver[3][8].run()  ;
            end

            begin
              gen[3][9].run()  ;
            end
            begin
              drv[3][9].run()  ;
            end
            begin
              mem_check[3][9].run()  ;
            end
            begin
              rf_driver[3][9].run()  ;
            end

            begin
              gen[3][10].run()  ;
            end
            begin
              drv[3][10].run()  ;
            end
            begin
              mem_check[3][10].run()  ;
            end
            begin
              rf_driver[3][10].run()  ;
            end

            begin
              gen[3][11].run()  ;
            end
            begin
              drv[3][11].run()  ;
            end
            begin
              mem_check[3][11].run()  ;
            end
            begin
              rf_driver[3][11].run()  ;
            end

            begin
              gen[3][12].run()  ;
            end
            begin
              drv[3][12].run()  ;
            end
            begin
              mem_check[3][12].run()  ;
            end
            begin
              rf_driver[3][12].run()  ;
            end

            begin
              gen[3][13].run()  ;
            end
            begin
              drv[3][13].run()  ;
            end
            begin
              mem_check[3][13].run()  ;
            end
            begin
              rf_driver[3][13].run()  ;
            end

            begin
              gen[3][14].run()  ;
            end
            begin
              drv[3][14].run()  ;
            end
            begin
              mem_check[3][14].run()  ;
            end
            begin
              rf_driver[3][14].run()  ;
            end

            begin
              gen[3][15].run()  ;
            end
            begin
              drv[3][15].run()  ;
            end
            begin
              mem_check[3][15].run()  ;
            end
            begin
              rf_driver[3][15].run()  ;
            end

            begin
              gen[3][16].run()  ;
            end
            begin
              drv[3][16].run()  ;
            end
            begin
              mem_check[3][16].run()  ;
            end
            begin
              rf_driver[3][16].run()  ;
            end

            begin
              gen[3][17].run()  ;
            end
            begin
              drv[3][17].run()  ;
            end
            begin
              mem_check[3][17].run()  ;
            end
            begin
              rf_driver[3][17].run()  ;
            end

            begin
              gen[3][18].run()  ;
            end
            begin
              drv[3][18].run()  ;
            end
            begin
              mem_check[3][18].run()  ;
            end
            begin
              rf_driver[3][18].run()  ;
            end

            begin
              gen[3][19].run()  ;
            end
            begin
              drv[3][19].run()  ;
            end
            begin
              mem_check[3][19].run()  ;
            end
            begin
              rf_driver[3][19].run()  ;
            end

            begin
              gen[3][20].run()  ;
            end
            begin
              drv[3][20].run()  ;
            end
            begin
              mem_check[3][20].run()  ;
            end
            begin
              rf_driver[3][20].run()  ;
            end

            begin
              gen[3][21].run()  ;
            end
            begin
              drv[3][21].run()  ;
            end
            begin
              mem_check[3][21].run()  ;
            end
            begin
              rf_driver[3][21].run()  ;
            end

            begin
              gen[3][22].run()  ;
            end
            begin
              drv[3][22].run()  ;
            end
            begin
              mem_check[3][22].run()  ;
            end
            begin
              rf_driver[3][22].run()  ;
            end

            begin
              gen[3][23].run()  ;
            end
            begin
              drv[3][23].run()  ;
            end
            begin
              mem_check[3][23].run()  ;
            end
            begin
              rf_driver[3][23].run()  ;
            end

            begin
              gen[3][24].run()  ;
            end
            begin
              drv[3][24].run()  ;
            end
            begin
              mem_check[3][24].run()  ;
            end
            begin
              rf_driver[3][24].run()  ;
            end

            begin
              gen[3][25].run()  ;
            end
            begin
              drv[3][25].run()  ;
            end
            begin
              mem_check[3][25].run()  ;
            end
            begin
              rf_driver[3][25].run()  ;
            end

            begin
              gen[3][26].run()  ;
            end
            begin
              drv[3][26].run()  ;
            end
            begin
              mem_check[3][26].run()  ;
            end
            begin
              rf_driver[3][26].run()  ;
            end

            begin
              gen[3][27].run()  ;
            end
            begin
              drv[3][27].run()  ;
            end
            begin
              mem_check[3][27].run()  ;
            end
            begin
              rf_driver[3][27].run()  ;
            end

            begin
              gen[3][28].run()  ;
            end
            begin
              drv[3][28].run()  ;
            end
            begin
              mem_check[3][28].run()  ;
            end
            begin
              rf_driver[3][28].run()  ;
            end

            begin
              gen[3][29].run()  ;
            end
            begin
              drv[3][29].run()  ;
            end
            begin
              mem_check[3][29].run()  ;
            end
            begin
              rf_driver[3][29].run()  ;
            end

            begin
              gen[3][30].run()  ;
            end
            begin
              drv[3][30].run()  ;
            end
            begin
              mem_check[3][30].run()  ;
            end
            begin
              rf_driver[3][30].run()  ;
            end

            begin
              gen[3][31].run()  ;
            end
            begin
              drv[3][31].run()  ;
            end
            begin
              mem_check[3][31].run()  ;
            end
            begin
              rf_driver[3][31].run()  ;
            end

            begin
              ldst_driver[4].run()  ;
            end
            begin
              mgr[4].run()  ;
            end
            begin
              oob_drv[4].run()  ;
            end
            begin
              up_check[4].run()  ;
            end
            begin
              gen[4][0].run()  ;
            end
            begin
              drv[4][0].run()  ;
            end
            begin
              mem_check[4][0].run()  ;
            end
            begin
              rf_driver[4][0].run()  ;
            end

            begin
              gen[4][1].run()  ;
            end
            begin
              drv[4][1].run()  ;
            end
            begin
              mem_check[4][1].run()  ;
            end
            begin
              rf_driver[4][1].run()  ;
            end

            begin
              gen[4][2].run()  ;
            end
            begin
              drv[4][2].run()  ;
            end
            begin
              mem_check[4][2].run()  ;
            end
            begin
              rf_driver[4][2].run()  ;
            end

            begin
              gen[4][3].run()  ;
            end
            begin
              drv[4][3].run()  ;
            end
            begin
              mem_check[4][3].run()  ;
            end
            begin
              rf_driver[4][3].run()  ;
            end

            begin
              gen[4][4].run()  ;
            end
            begin
              drv[4][4].run()  ;
            end
            begin
              mem_check[4][4].run()  ;
            end
            begin
              rf_driver[4][4].run()  ;
            end

            begin
              gen[4][5].run()  ;
            end
            begin
              drv[4][5].run()  ;
            end
            begin
              mem_check[4][5].run()  ;
            end
            begin
              rf_driver[4][5].run()  ;
            end

            begin
              gen[4][6].run()  ;
            end
            begin
              drv[4][6].run()  ;
            end
            begin
              mem_check[4][6].run()  ;
            end
            begin
              rf_driver[4][6].run()  ;
            end

            begin
              gen[4][7].run()  ;
            end
            begin
              drv[4][7].run()  ;
            end
            begin
              mem_check[4][7].run()  ;
            end
            begin
              rf_driver[4][7].run()  ;
            end

            begin
              gen[4][8].run()  ;
            end
            begin
              drv[4][8].run()  ;
            end
            begin
              mem_check[4][8].run()  ;
            end
            begin
              rf_driver[4][8].run()  ;
            end

            begin
              gen[4][9].run()  ;
            end
            begin
              drv[4][9].run()  ;
            end
            begin
              mem_check[4][9].run()  ;
            end
            begin
              rf_driver[4][9].run()  ;
            end

            begin
              gen[4][10].run()  ;
            end
            begin
              drv[4][10].run()  ;
            end
            begin
              mem_check[4][10].run()  ;
            end
            begin
              rf_driver[4][10].run()  ;
            end

            begin
              gen[4][11].run()  ;
            end
            begin
              drv[4][11].run()  ;
            end
            begin
              mem_check[4][11].run()  ;
            end
            begin
              rf_driver[4][11].run()  ;
            end

            begin
              gen[4][12].run()  ;
            end
            begin
              drv[4][12].run()  ;
            end
            begin
              mem_check[4][12].run()  ;
            end
            begin
              rf_driver[4][12].run()  ;
            end

            begin
              gen[4][13].run()  ;
            end
            begin
              drv[4][13].run()  ;
            end
            begin
              mem_check[4][13].run()  ;
            end
            begin
              rf_driver[4][13].run()  ;
            end

            begin
              gen[4][14].run()  ;
            end
            begin
              drv[4][14].run()  ;
            end
            begin
              mem_check[4][14].run()  ;
            end
            begin
              rf_driver[4][14].run()  ;
            end

            begin
              gen[4][15].run()  ;
            end
            begin
              drv[4][15].run()  ;
            end
            begin
              mem_check[4][15].run()  ;
            end
            begin
              rf_driver[4][15].run()  ;
            end

            begin
              gen[4][16].run()  ;
            end
            begin
              drv[4][16].run()  ;
            end
            begin
              mem_check[4][16].run()  ;
            end
            begin
              rf_driver[4][16].run()  ;
            end

            begin
              gen[4][17].run()  ;
            end
            begin
              drv[4][17].run()  ;
            end
            begin
              mem_check[4][17].run()  ;
            end
            begin
              rf_driver[4][17].run()  ;
            end

            begin
              gen[4][18].run()  ;
            end
            begin
              drv[4][18].run()  ;
            end
            begin
              mem_check[4][18].run()  ;
            end
            begin
              rf_driver[4][18].run()  ;
            end

            begin
              gen[4][19].run()  ;
            end
            begin
              drv[4][19].run()  ;
            end
            begin
              mem_check[4][19].run()  ;
            end
            begin
              rf_driver[4][19].run()  ;
            end

            begin
              gen[4][20].run()  ;
            end
            begin
              drv[4][20].run()  ;
            end
            begin
              mem_check[4][20].run()  ;
            end
            begin
              rf_driver[4][20].run()  ;
            end

            begin
              gen[4][21].run()  ;
            end
            begin
              drv[4][21].run()  ;
            end
            begin
              mem_check[4][21].run()  ;
            end
            begin
              rf_driver[4][21].run()  ;
            end

            begin
              gen[4][22].run()  ;
            end
            begin
              drv[4][22].run()  ;
            end
            begin
              mem_check[4][22].run()  ;
            end
            begin
              rf_driver[4][22].run()  ;
            end

            begin
              gen[4][23].run()  ;
            end
            begin
              drv[4][23].run()  ;
            end
            begin
              mem_check[4][23].run()  ;
            end
            begin
              rf_driver[4][23].run()  ;
            end

            begin
              gen[4][24].run()  ;
            end
            begin
              drv[4][24].run()  ;
            end
            begin
              mem_check[4][24].run()  ;
            end
            begin
              rf_driver[4][24].run()  ;
            end

            begin
              gen[4][25].run()  ;
            end
            begin
              drv[4][25].run()  ;
            end
            begin
              mem_check[4][25].run()  ;
            end
            begin
              rf_driver[4][25].run()  ;
            end

            begin
              gen[4][26].run()  ;
            end
            begin
              drv[4][26].run()  ;
            end
            begin
              mem_check[4][26].run()  ;
            end
            begin
              rf_driver[4][26].run()  ;
            end

            begin
              gen[4][27].run()  ;
            end
            begin
              drv[4][27].run()  ;
            end
            begin
              mem_check[4][27].run()  ;
            end
            begin
              rf_driver[4][27].run()  ;
            end

            begin
              gen[4][28].run()  ;
            end
            begin
              drv[4][28].run()  ;
            end
            begin
              mem_check[4][28].run()  ;
            end
            begin
              rf_driver[4][28].run()  ;
            end

            begin
              gen[4][29].run()  ;
            end
            begin
              drv[4][29].run()  ;
            end
            begin
              mem_check[4][29].run()  ;
            end
            begin
              rf_driver[4][29].run()  ;
            end

            begin
              gen[4][30].run()  ;
            end
            begin
              drv[4][30].run()  ;
            end
            begin
              mem_check[4][30].run()  ;
            end
            begin
              rf_driver[4][30].run()  ;
            end

            begin
              gen[4][31].run()  ;
            end
            begin
              drv[4][31].run()  ;
            end
            begin
              mem_check[4][31].run()  ;
            end
            begin
              rf_driver[4][31].run()  ;
            end

            begin
              ldst_driver[5].run()  ;
            end
            begin
              mgr[5].run()  ;
            end
            begin
              oob_drv[5].run()  ;
            end
            begin
              up_check[5].run()  ;
            end
            begin
              gen[5][0].run()  ;
            end
            begin
              drv[5][0].run()  ;
            end
            begin
              mem_check[5][0].run()  ;
            end
            begin
              rf_driver[5][0].run()  ;
            end

            begin
              gen[5][1].run()  ;
            end
            begin
              drv[5][1].run()  ;
            end
            begin
              mem_check[5][1].run()  ;
            end
            begin
              rf_driver[5][1].run()  ;
            end

            begin
              gen[5][2].run()  ;
            end
            begin
              drv[5][2].run()  ;
            end
            begin
              mem_check[5][2].run()  ;
            end
            begin
              rf_driver[5][2].run()  ;
            end

            begin
              gen[5][3].run()  ;
            end
            begin
              drv[5][3].run()  ;
            end
            begin
              mem_check[5][3].run()  ;
            end
            begin
              rf_driver[5][3].run()  ;
            end

            begin
              gen[5][4].run()  ;
            end
            begin
              drv[5][4].run()  ;
            end
            begin
              mem_check[5][4].run()  ;
            end
            begin
              rf_driver[5][4].run()  ;
            end

            begin
              gen[5][5].run()  ;
            end
            begin
              drv[5][5].run()  ;
            end
            begin
              mem_check[5][5].run()  ;
            end
            begin
              rf_driver[5][5].run()  ;
            end

            begin
              gen[5][6].run()  ;
            end
            begin
              drv[5][6].run()  ;
            end
            begin
              mem_check[5][6].run()  ;
            end
            begin
              rf_driver[5][6].run()  ;
            end

            begin
              gen[5][7].run()  ;
            end
            begin
              drv[5][7].run()  ;
            end
            begin
              mem_check[5][7].run()  ;
            end
            begin
              rf_driver[5][7].run()  ;
            end

            begin
              gen[5][8].run()  ;
            end
            begin
              drv[5][8].run()  ;
            end
            begin
              mem_check[5][8].run()  ;
            end
            begin
              rf_driver[5][8].run()  ;
            end

            begin
              gen[5][9].run()  ;
            end
            begin
              drv[5][9].run()  ;
            end
            begin
              mem_check[5][9].run()  ;
            end
            begin
              rf_driver[5][9].run()  ;
            end

            begin
              gen[5][10].run()  ;
            end
            begin
              drv[5][10].run()  ;
            end
            begin
              mem_check[5][10].run()  ;
            end
            begin
              rf_driver[5][10].run()  ;
            end

            begin
              gen[5][11].run()  ;
            end
            begin
              drv[5][11].run()  ;
            end
            begin
              mem_check[5][11].run()  ;
            end
            begin
              rf_driver[5][11].run()  ;
            end

            begin
              gen[5][12].run()  ;
            end
            begin
              drv[5][12].run()  ;
            end
            begin
              mem_check[5][12].run()  ;
            end
            begin
              rf_driver[5][12].run()  ;
            end

            begin
              gen[5][13].run()  ;
            end
            begin
              drv[5][13].run()  ;
            end
            begin
              mem_check[5][13].run()  ;
            end
            begin
              rf_driver[5][13].run()  ;
            end

            begin
              gen[5][14].run()  ;
            end
            begin
              drv[5][14].run()  ;
            end
            begin
              mem_check[5][14].run()  ;
            end
            begin
              rf_driver[5][14].run()  ;
            end

            begin
              gen[5][15].run()  ;
            end
            begin
              drv[5][15].run()  ;
            end
            begin
              mem_check[5][15].run()  ;
            end
            begin
              rf_driver[5][15].run()  ;
            end

            begin
              gen[5][16].run()  ;
            end
            begin
              drv[5][16].run()  ;
            end
            begin
              mem_check[5][16].run()  ;
            end
            begin
              rf_driver[5][16].run()  ;
            end

            begin
              gen[5][17].run()  ;
            end
            begin
              drv[5][17].run()  ;
            end
            begin
              mem_check[5][17].run()  ;
            end
            begin
              rf_driver[5][17].run()  ;
            end

            begin
              gen[5][18].run()  ;
            end
            begin
              drv[5][18].run()  ;
            end
            begin
              mem_check[5][18].run()  ;
            end
            begin
              rf_driver[5][18].run()  ;
            end

            begin
              gen[5][19].run()  ;
            end
            begin
              drv[5][19].run()  ;
            end
            begin
              mem_check[5][19].run()  ;
            end
            begin
              rf_driver[5][19].run()  ;
            end

            begin
              gen[5][20].run()  ;
            end
            begin
              drv[5][20].run()  ;
            end
            begin
              mem_check[5][20].run()  ;
            end
            begin
              rf_driver[5][20].run()  ;
            end

            begin
              gen[5][21].run()  ;
            end
            begin
              drv[5][21].run()  ;
            end
            begin
              mem_check[5][21].run()  ;
            end
            begin
              rf_driver[5][21].run()  ;
            end

            begin
              gen[5][22].run()  ;
            end
            begin
              drv[5][22].run()  ;
            end
            begin
              mem_check[5][22].run()  ;
            end
            begin
              rf_driver[5][22].run()  ;
            end

            begin
              gen[5][23].run()  ;
            end
            begin
              drv[5][23].run()  ;
            end
            begin
              mem_check[5][23].run()  ;
            end
            begin
              rf_driver[5][23].run()  ;
            end

            begin
              gen[5][24].run()  ;
            end
            begin
              drv[5][24].run()  ;
            end
            begin
              mem_check[5][24].run()  ;
            end
            begin
              rf_driver[5][24].run()  ;
            end

            begin
              gen[5][25].run()  ;
            end
            begin
              drv[5][25].run()  ;
            end
            begin
              mem_check[5][25].run()  ;
            end
            begin
              rf_driver[5][25].run()  ;
            end

            begin
              gen[5][26].run()  ;
            end
            begin
              drv[5][26].run()  ;
            end
            begin
              mem_check[5][26].run()  ;
            end
            begin
              rf_driver[5][26].run()  ;
            end

            begin
              gen[5][27].run()  ;
            end
            begin
              drv[5][27].run()  ;
            end
            begin
              mem_check[5][27].run()  ;
            end
            begin
              rf_driver[5][27].run()  ;
            end

            begin
              gen[5][28].run()  ;
            end
            begin
              drv[5][28].run()  ;
            end
            begin
              mem_check[5][28].run()  ;
            end
            begin
              rf_driver[5][28].run()  ;
            end

            begin
              gen[5][29].run()  ;
            end
            begin
              drv[5][29].run()  ;
            end
            begin
              mem_check[5][29].run()  ;
            end
            begin
              rf_driver[5][29].run()  ;
            end

            begin
              gen[5][30].run()  ;
            end
            begin
              drv[5][30].run()  ;
            end
            begin
              mem_check[5][30].run()  ;
            end
            begin
              rf_driver[5][30].run()  ;
            end

            begin
              gen[5][31].run()  ;
            end
            begin
              drv[5][31].run()  ;
            end
            begin
              mem_check[5][31].run()  ;
            end
            begin
              rf_driver[5][31].run()  ;
            end

            begin
              ldst_driver[6].run()  ;
            end
            begin
              mgr[6].run()  ;
            end
            begin
              oob_drv[6].run()  ;
            end
            begin
              up_check[6].run()  ;
            end
            begin
              gen[6][0].run()  ;
            end
            begin
              drv[6][0].run()  ;
            end
            begin
              mem_check[6][0].run()  ;
            end
            begin
              rf_driver[6][0].run()  ;
            end

            begin
              gen[6][1].run()  ;
            end
            begin
              drv[6][1].run()  ;
            end
            begin
              mem_check[6][1].run()  ;
            end
            begin
              rf_driver[6][1].run()  ;
            end

            begin
              gen[6][2].run()  ;
            end
            begin
              drv[6][2].run()  ;
            end
            begin
              mem_check[6][2].run()  ;
            end
            begin
              rf_driver[6][2].run()  ;
            end

            begin
              gen[6][3].run()  ;
            end
            begin
              drv[6][3].run()  ;
            end
            begin
              mem_check[6][3].run()  ;
            end
            begin
              rf_driver[6][3].run()  ;
            end

            begin
              gen[6][4].run()  ;
            end
            begin
              drv[6][4].run()  ;
            end
            begin
              mem_check[6][4].run()  ;
            end
            begin
              rf_driver[6][4].run()  ;
            end

            begin
              gen[6][5].run()  ;
            end
            begin
              drv[6][5].run()  ;
            end
            begin
              mem_check[6][5].run()  ;
            end
            begin
              rf_driver[6][5].run()  ;
            end

            begin
              gen[6][6].run()  ;
            end
            begin
              drv[6][6].run()  ;
            end
            begin
              mem_check[6][6].run()  ;
            end
            begin
              rf_driver[6][6].run()  ;
            end

            begin
              gen[6][7].run()  ;
            end
            begin
              drv[6][7].run()  ;
            end
            begin
              mem_check[6][7].run()  ;
            end
            begin
              rf_driver[6][7].run()  ;
            end

            begin
              gen[6][8].run()  ;
            end
            begin
              drv[6][8].run()  ;
            end
            begin
              mem_check[6][8].run()  ;
            end
            begin
              rf_driver[6][8].run()  ;
            end

            begin
              gen[6][9].run()  ;
            end
            begin
              drv[6][9].run()  ;
            end
            begin
              mem_check[6][9].run()  ;
            end
            begin
              rf_driver[6][9].run()  ;
            end

            begin
              gen[6][10].run()  ;
            end
            begin
              drv[6][10].run()  ;
            end
            begin
              mem_check[6][10].run()  ;
            end
            begin
              rf_driver[6][10].run()  ;
            end

            begin
              gen[6][11].run()  ;
            end
            begin
              drv[6][11].run()  ;
            end
            begin
              mem_check[6][11].run()  ;
            end
            begin
              rf_driver[6][11].run()  ;
            end

            begin
              gen[6][12].run()  ;
            end
            begin
              drv[6][12].run()  ;
            end
            begin
              mem_check[6][12].run()  ;
            end
            begin
              rf_driver[6][12].run()  ;
            end

            begin
              gen[6][13].run()  ;
            end
            begin
              drv[6][13].run()  ;
            end
            begin
              mem_check[6][13].run()  ;
            end
            begin
              rf_driver[6][13].run()  ;
            end

            begin
              gen[6][14].run()  ;
            end
            begin
              drv[6][14].run()  ;
            end
            begin
              mem_check[6][14].run()  ;
            end
            begin
              rf_driver[6][14].run()  ;
            end

            begin
              gen[6][15].run()  ;
            end
            begin
              drv[6][15].run()  ;
            end
            begin
              mem_check[6][15].run()  ;
            end
            begin
              rf_driver[6][15].run()  ;
            end

            begin
              gen[6][16].run()  ;
            end
            begin
              drv[6][16].run()  ;
            end
            begin
              mem_check[6][16].run()  ;
            end
            begin
              rf_driver[6][16].run()  ;
            end

            begin
              gen[6][17].run()  ;
            end
            begin
              drv[6][17].run()  ;
            end
            begin
              mem_check[6][17].run()  ;
            end
            begin
              rf_driver[6][17].run()  ;
            end

            begin
              gen[6][18].run()  ;
            end
            begin
              drv[6][18].run()  ;
            end
            begin
              mem_check[6][18].run()  ;
            end
            begin
              rf_driver[6][18].run()  ;
            end

            begin
              gen[6][19].run()  ;
            end
            begin
              drv[6][19].run()  ;
            end
            begin
              mem_check[6][19].run()  ;
            end
            begin
              rf_driver[6][19].run()  ;
            end

            begin
              gen[6][20].run()  ;
            end
            begin
              drv[6][20].run()  ;
            end
            begin
              mem_check[6][20].run()  ;
            end
            begin
              rf_driver[6][20].run()  ;
            end

            begin
              gen[6][21].run()  ;
            end
            begin
              drv[6][21].run()  ;
            end
            begin
              mem_check[6][21].run()  ;
            end
            begin
              rf_driver[6][21].run()  ;
            end

            begin
              gen[6][22].run()  ;
            end
            begin
              drv[6][22].run()  ;
            end
            begin
              mem_check[6][22].run()  ;
            end
            begin
              rf_driver[6][22].run()  ;
            end

            begin
              gen[6][23].run()  ;
            end
            begin
              drv[6][23].run()  ;
            end
            begin
              mem_check[6][23].run()  ;
            end
            begin
              rf_driver[6][23].run()  ;
            end

            begin
              gen[6][24].run()  ;
            end
            begin
              drv[6][24].run()  ;
            end
            begin
              mem_check[6][24].run()  ;
            end
            begin
              rf_driver[6][24].run()  ;
            end

            begin
              gen[6][25].run()  ;
            end
            begin
              drv[6][25].run()  ;
            end
            begin
              mem_check[6][25].run()  ;
            end
            begin
              rf_driver[6][25].run()  ;
            end

            begin
              gen[6][26].run()  ;
            end
            begin
              drv[6][26].run()  ;
            end
            begin
              mem_check[6][26].run()  ;
            end
            begin
              rf_driver[6][26].run()  ;
            end

            begin
              gen[6][27].run()  ;
            end
            begin
              drv[6][27].run()  ;
            end
            begin
              mem_check[6][27].run()  ;
            end
            begin
              rf_driver[6][27].run()  ;
            end

            begin
              gen[6][28].run()  ;
            end
            begin
              drv[6][28].run()  ;
            end
            begin
              mem_check[6][28].run()  ;
            end
            begin
              rf_driver[6][28].run()  ;
            end

            begin
              gen[6][29].run()  ;
            end
            begin
              drv[6][29].run()  ;
            end
            begin
              mem_check[6][29].run()  ;
            end
            begin
              rf_driver[6][29].run()  ;
            end

            begin
              gen[6][30].run()  ;
            end
            begin
              drv[6][30].run()  ;
            end
            begin
              mem_check[6][30].run()  ;
            end
            begin
              rf_driver[6][30].run()  ;
            end

            begin
              gen[6][31].run()  ;
            end
            begin
              drv[6][31].run()  ;
            end
            begin
              mem_check[6][31].run()  ;
            end
            begin
              rf_driver[6][31].run()  ;
            end

            begin
              ldst_driver[7].run()  ;
            end
            begin
              mgr[7].run()  ;
            end
            begin
              oob_drv[7].run()  ;
            end
            begin
              up_check[7].run()  ;
            end
            begin
              gen[7][0].run()  ;
            end
            begin
              drv[7][0].run()  ;
            end
            begin
              mem_check[7][0].run()  ;
            end
            begin
              rf_driver[7][0].run()  ;
            end

            begin
              gen[7][1].run()  ;
            end
            begin
              drv[7][1].run()  ;
            end
            begin
              mem_check[7][1].run()  ;
            end
            begin
              rf_driver[7][1].run()  ;
            end

            begin
              gen[7][2].run()  ;
            end
            begin
              drv[7][2].run()  ;
            end
            begin
              mem_check[7][2].run()  ;
            end
            begin
              rf_driver[7][2].run()  ;
            end

            begin
              gen[7][3].run()  ;
            end
            begin
              drv[7][3].run()  ;
            end
            begin
              mem_check[7][3].run()  ;
            end
            begin
              rf_driver[7][3].run()  ;
            end

            begin
              gen[7][4].run()  ;
            end
            begin
              drv[7][4].run()  ;
            end
            begin
              mem_check[7][4].run()  ;
            end
            begin
              rf_driver[7][4].run()  ;
            end

            begin
              gen[7][5].run()  ;
            end
            begin
              drv[7][5].run()  ;
            end
            begin
              mem_check[7][5].run()  ;
            end
            begin
              rf_driver[7][5].run()  ;
            end

            begin
              gen[7][6].run()  ;
            end
            begin
              drv[7][6].run()  ;
            end
            begin
              mem_check[7][6].run()  ;
            end
            begin
              rf_driver[7][6].run()  ;
            end

            begin
              gen[7][7].run()  ;
            end
            begin
              drv[7][7].run()  ;
            end
            begin
              mem_check[7][7].run()  ;
            end
            begin
              rf_driver[7][7].run()  ;
            end

            begin
              gen[7][8].run()  ;
            end
            begin
              drv[7][8].run()  ;
            end
            begin
              mem_check[7][8].run()  ;
            end
            begin
              rf_driver[7][8].run()  ;
            end

            begin
              gen[7][9].run()  ;
            end
            begin
              drv[7][9].run()  ;
            end
            begin
              mem_check[7][9].run()  ;
            end
            begin
              rf_driver[7][9].run()  ;
            end

            begin
              gen[7][10].run()  ;
            end
            begin
              drv[7][10].run()  ;
            end
            begin
              mem_check[7][10].run()  ;
            end
            begin
              rf_driver[7][10].run()  ;
            end

            begin
              gen[7][11].run()  ;
            end
            begin
              drv[7][11].run()  ;
            end
            begin
              mem_check[7][11].run()  ;
            end
            begin
              rf_driver[7][11].run()  ;
            end

            begin
              gen[7][12].run()  ;
            end
            begin
              drv[7][12].run()  ;
            end
            begin
              mem_check[7][12].run()  ;
            end
            begin
              rf_driver[7][12].run()  ;
            end

            begin
              gen[7][13].run()  ;
            end
            begin
              drv[7][13].run()  ;
            end
            begin
              mem_check[7][13].run()  ;
            end
            begin
              rf_driver[7][13].run()  ;
            end

            begin
              gen[7][14].run()  ;
            end
            begin
              drv[7][14].run()  ;
            end
            begin
              mem_check[7][14].run()  ;
            end
            begin
              rf_driver[7][14].run()  ;
            end

            begin
              gen[7][15].run()  ;
            end
            begin
              drv[7][15].run()  ;
            end
            begin
              mem_check[7][15].run()  ;
            end
            begin
              rf_driver[7][15].run()  ;
            end

            begin
              gen[7][16].run()  ;
            end
            begin
              drv[7][16].run()  ;
            end
            begin
              mem_check[7][16].run()  ;
            end
            begin
              rf_driver[7][16].run()  ;
            end

            begin
              gen[7][17].run()  ;
            end
            begin
              drv[7][17].run()  ;
            end
            begin
              mem_check[7][17].run()  ;
            end
            begin
              rf_driver[7][17].run()  ;
            end

            begin
              gen[7][18].run()  ;
            end
            begin
              drv[7][18].run()  ;
            end
            begin
              mem_check[7][18].run()  ;
            end
            begin
              rf_driver[7][18].run()  ;
            end

            begin
              gen[7][19].run()  ;
            end
            begin
              drv[7][19].run()  ;
            end
            begin
              mem_check[7][19].run()  ;
            end
            begin
              rf_driver[7][19].run()  ;
            end

            begin
              gen[7][20].run()  ;
            end
            begin
              drv[7][20].run()  ;
            end
            begin
              mem_check[7][20].run()  ;
            end
            begin
              rf_driver[7][20].run()  ;
            end

            begin
              gen[7][21].run()  ;
            end
            begin
              drv[7][21].run()  ;
            end
            begin
              mem_check[7][21].run()  ;
            end
            begin
              rf_driver[7][21].run()  ;
            end

            begin
              gen[7][22].run()  ;
            end
            begin
              drv[7][22].run()  ;
            end
            begin
              mem_check[7][22].run()  ;
            end
            begin
              rf_driver[7][22].run()  ;
            end

            begin
              gen[7][23].run()  ;
            end
            begin
              drv[7][23].run()  ;
            end
            begin
              mem_check[7][23].run()  ;
            end
            begin
              rf_driver[7][23].run()  ;
            end

            begin
              gen[7][24].run()  ;
            end
            begin
              drv[7][24].run()  ;
            end
            begin
              mem_check[7][24].run()  ;
            end
            begin
              rf_driver[7][24].run()  ;
            end

            begin
              gen[7][25].run()  ;
            end
            begin
              drv[7][25].run()  ;
            end
            begin
              mem_check[7][25].run()  ;
            end
            begin
              rf_driver[7][25].run()  ;
            end

            begin
              gen[7][26].run()  ;
            end
            begin
              drv[7][26].run()  ;
            end
            begin
              mem_check[7][26].run()  ;
            end
            begin
              rf_driver[7][26].run()  ;
            end

            begin
              gen[7][27].run()  ;
            end
            begin
              drv[7][27].run()  ;
            end
            begin
              mem_check[7][27].run()  ;
            end
            begin
              rf_driver[7][27].run()  ;
            end

            begin
              gen[7][28].run()  ;
            end
            begin
              drv[7][28].run()  ;
            end
            begin
              mem_check[7][28].run()  ;
            end
            begin
              rf_driver[7][28].run()  ;
            end

            begin
              gen[7][29].run()  ;
            end
            begin
              drv[7][29].run()  ;
            end
            begin
              mem_check[7][29].run()  ;
            end
            begin
              rf_driver[7][29].run()  ;
            end

            begin
              gen[7][30].run()  ;
            end
            begin
              drv[7][30].run()  ;
            end
            begin
              mem_check[7][30].run()  ;
            end
            begin
              rf_driver[7][30].run()  ;
            end

            begin
              gen[7][31].run()  ;
            end
            begin
              drv[7][31].run()  ;
            end
            begin
              mem_check[7][31].run()  ;
            end
            begin
              rf_driver[7][31].run()  ;
            end

            begin
              ldst_driver[8].run()  ;
            end
            begin
              mgr[8].run()  ;
            end
            begin
              oob_drv[8].run()  ;
            end
            begin
              up_check[8].run()  ;
            end
            begin
              gen[8][0].run()  ;
            end
            begin
              drv[8][0].run()  ;
            end
            begin
              mem_check[8][0].run()  ;
            end
            begin
              rf_driver[8][0].run()  ;
            end

            begin
              gen[8][1].run()  ;
            end
            begin
              drv[8][1].run()  ;
            end
            begin
              mem_check[8][1].run()  ;
            end
            begin
              rf_driver[8][1].run()  ;
            end

            begin
              gen[8][2].run()  ;
            end
            begin
              drv[8][2].run()  ;
            end
            begin
              mem_check[8][2].run()  ;
            end
            begin
              rf_driver[8][2].run()  ;
            end

            begin
              gen[8][3].run()  ;
            end
            begin
              drv[8][3].run()  ;
            end
            begin
              mem_check[8][3].run()  ;
            end
            begin
              rf_driver[8][3].run()  ;
            end

            begin
              gen[8][4].run()  ;
            end
            begin
              drv[8][4].run()  ;
            end
            begin
              mem_check[8][4].run()  ;
            end
            begin
              rf_driver[8][4].run()  ;
            end

            begin
              gen[8][5].run()  ;
            end
            begin
              drv[8][5].run()  ;
            end
            begin
              mem_check[8][5].run()  ;
            end
            begin
              rf_driver[8][5].run()  ;
            end

            begin
              gen[8][6].run()  ;
            end
            begin
              drv[8][6].run()  ;
            end
            begin
              mem_check[8][6].run()  ;
            end
            begin
              rf_driver[8][6].run()  ;
            end

            begin
              gen[8][7].run()  ;
            end
            begin
              drv[8][7].run()  ;
            end
            begin
              mem_check[8][7].run()  ;
            end
            begin
              rf_driver[8][7].run()  ;
            end

            begin
              gen[8][8].run()  ;
            end
            begin
              drv[8][8].run()  ;
            end
            begin
              mem_check[8][8].run()  ;
            end
            begin
              rf_driver[8][8].run()  ;
            end

            begin
              gen[8][9].run()  ;
            end
            begin
              drv[8][9].run()  ;
            end
            begin
              mem_check[8][9].run()  ;
            end
            begin
              rf_driver[8][9].run()  ;
            end

            begin
              gen[8][10].run()  ;
            end
            begin
              drv[8][10].run()  ;
            end
            begin
              mem_check[8][10].run()  ;
            end
            begin
              rf_driver[8][10].run()  ;
            end

            begin
              gen[8][11].run()  ;
            end
            begin
              drv[8][11].run()  ;
            end
            begin
              mem_check[8][11].run()  ;
            end
            begin
              rf_driver[8][11].run()  ;
            end

            begin
              gen[8][12].run()  ;
            end
            begin
              drv[8][12].run()  ;
            end
            begin
              mem_check[8][12].run()  ;
            end
            begin
              rf_driver[8][12].run()  ;
            end

            begin
              gen[8][13].run()  ;
            end
            begin
              drv[8][13].run()  ;
            end
            begin
              mem_check[8][13].run()  ;
            end
            begin
              rf_driver[8][13].run()  ;
            end

            begin
              gen[8][14].run()  ;
            end
            begin
              drv[8][14].run()  ;
            end
            begin
              mem_check[8][14].run()  ;
            end
            begin
              rf_driver[8][14].run()  ;
            end

            begin
              gen[8][15].run()  ;
            end
            begin
              drv[8][15].run()  ;
            end
            begin
              mem_check[8][15].run()  ;
            end
            begin
              rf_driver[8][15].run()  ;
            end

            begin
              gen[8][16].run()  ;
            end
            begin
              drv[8][16].run()  ;
            end
            begin
              mem_check[8][16].run()  ;
            end
            begin
              rf_driver[8][16].run()  ;
            end

            begin
              gen[8][17].run()  ;
            end
            begin
              drv[8][17].run()  ;
            end
            begin
              mem_check[8][17].run()  ;
            end
            begin
              rf_driver[8][17].run()  ;
            end

            begin
              gen[8][18].run()  ;
            end
            begin
              drv[8][18].run()  ;
            end
            begin
              mem_check[8][18].run()  ;
            end
            begin
              rf_driver[8][18].run()  ;
            end

            begin
              gen[8][19].run()  ;
            end
            begin
              drv[8][19].run()  ;
            end
            begin
              mem_check[8][19].run()  ;
            end
            begin
              rf_driver[8][19].run()  ;
            end

            begin
              gen[8][20].run()  ;
            end
            begin
              drv[8][20].run()  ;
            end
            begin
              mem_check[8][20].run()  ;
            end
            begin
              rf_driver[8][20].run()  ;
            end

            begin
              gen[8][21].run()  ;
            end
            begin
              drv[8][21].run()  ;
            end
            begin
              mem_check[8][21].run()  ;
            end
            begin
              rf_driver[8][21].run()  ;
            end

            begin
              gen[8][22].run()  ;
            end
            begin
              drv[8][22].run()  ;
            end
            begin
              mem_check[8][22].run()  ;
            end
            begin
              rf_driver[8][22].run()  ;
            end

            begin
              gen[8][23].run()  ;
            end
            begin
              drv[8][23].run()  ;
            end
            begin
              mem_check[8][23].run()  ;
            end
            begin
              rf_driver[8][23].run()  ;
            end

            begin
              gen[8][24].run()  ;
            end
            begin
              drv[8][24].run()  ;
            end
            begin
              mem_check[8][24].run()  ;
            end
            begin
              rf_driver[8][24].run()  ;
            end

            begin
              gen[8][25].run()  ;
            end
            begin
              drv[8][25].run()  ;
            end
            begin
              mem_check[8][25].run()  ;
            end
            begin
              rf_driver[8][25].run()  ;
            end

            begin
              gen[8][26].run()  ;
            end
            begin
              drv[8][26].run()  ;
            end
            begin
              mem_check[8][26].run()  ;
            end
            begin
              rf_driver[8][26].run()  ;
            end

            begin
              gen[8][27].run()  ;
            end
            begin
              drv[8][27].run()  ;
            end
            begin
              mem_check[8][27].run()  ;
            end
            begin
              rf_driver[8][27].run()  ;
            end

            begin
              gen[8][28].run()  ;
            end
            begin
              drv[8][28].run()  ;
            end
            begin
              mem_check[8][28].run()  ;
            end
            begin
              rf_driver[8][28].run()  ;
            end

            begin
              gen[8][29].run()  ;
            end
            begin
              drv[8][29].run()  ;
            end
            begin
              mem_check[8][29].run()  ;
            end
            begin
              rf_driver[8][29].run()  ;
            end

            begin
              gen[8][30].run()  ;
            end
            begin
              drv[8][30].run()  ;
            end
            begin
              mem_check[8][30].run()  ;
            end
            begin
              rf_driver[8][30].run()  ;
            end

            begin
              gen[8][31].run()  ;
            end
            begin
              drv[8][31].run()  ;
            end
            begin
              mem_check[8][31].run()  ;
            end
            begin
              rf_driver[8][31].run()  ;
            end

            begin
              ldst_driver[9].run()  ;
            end
            begin
              mgr[9].run()  ;
            end
            begin
              oob_drv[9].run()  ;
            end
            begin
              up_check[9].run()  ;
            end
            begin
              gen[9][0].run()  ;
            end
            begin
              drv[9][0].run()  ;
            end
            begin
              mem_check[9][0].run()  ;
            end
            begin
              rf_driver[9][0].run()  ;
            end

            begin
              gen[9][1].run()  ;
            end
            begin
              drv[9][1].run()  ;
            end
            begin
              mem_check[9][1].run()  ;
            end
            begin
              rf_driver[9][1].run()  ;
            end

            begin
              gen[9][2].run()  ;
            end
            begin
              drv[9][2].run()  ;
            end
            begin
              mem_check[9][2].run()  ;
            end
            begin
              rf_driver[9][2].run()  ;
            end

            begin
              gen[9][3].run()  ;
            end
            begin
              drv[9][3].run()  ;
            end
            begin
              mem_check[9][3].run()  ;
            end
            begin
              rf_driver[9][3].run()  ;
            end

            begin
              gen[9][4].run()  ;
            end
            begin
              drv[9][4].run()  ;
            end
            begin
              mem_check[9][4].run()  ;
            end
            begin
              rf_driver[9][4].run()  ;
            end

            begin
              gen[9][5].run()  ;
            end
            begin
              drv[9][5].run()  ;
            end
            begin
              mem_check[9][5].run()  ;
            end
            begin
              rf_driver[9][5].run()  ;
            end

            begin
              gen[9][6].run()  ;
            end
            begin
              drv[9][6].run()  ;
            end
            begin
              mem_check[9][6].run()  ;
            end
            begin
              rf_driver[9][6].run()  ;
            end

            begin
              gen[9][7].run()  ;
            end
            begin
              drv[9][7].run()  ;
            end
            begin
              mem_check[9][7].run()  ;
            end
            begin
              rf_driver[9][7].run()  ;
            end

            begin
              gen[9][8].run()  ;
            end
            begin
              drv[9][8].run()  ;
            end
            begin
              mem_check[9][8].run()  ;
            end
            begin
              rf_driver[9][8].run()  ;
            end

            begin
              gen[9][9].run()  ;
            end
            begin
              drv[9][9].run()  ;
            end
            begin
              mem_check[9][9].run()  ;
            end
            begin
              rf_driver[9][9].run()  ;
            end

            begin
              gen[9][10].run()  ;
            end
            begin
              drv[9][10].run()  ;
            end
            begin
              mem_check[9][10].run()  ;
            end
            begin
              rf_driver[9][10].run()  ;
            end

            begin
              gen[9][11].run()  ;
            end
            begin
              drv[9][11].run()  ;
            end
            begin
              mem_check[9][11].run()  ;
            end
            begin
              rf_driver[9][11].run()  ;
            end

            begin
              gen[9][12].run()  ;
            end
            begin
              drv[9][12].run()  ;
            end
            begin
              mem_check[9][12].run()  ;
            end
            begin
              rf_driver[9][12].run()  ;
            end

            begin
              gen[9][13].run()  ;
            end
            begin
              drv[9][13].run()  ;
            end
            begin
              mem_check[9][13].run()  ;
            end
            begin
              rf_driver[9][13].run()  ;
            end

            begin
              gen[9][14].run()  ;
            end
            begin
              drv[9][14].run()  ;
            end
            begin
              mem_check[9][14].run()  ;
            end
            begin
              rf_driver[9][14].run()  ;
            end

            begin
              gen[9][15].run()  ;
            end
            begin
              drv[9][15].run()  ;
            end
            begin
              mem_check[9][15].run()  ;
            end
            begin
              rf_driver[9][15].run()  ;
            end

            begin
              gen[9][16].run()  ;
            end
            begin
              drv[9][16].run()  ;
            end
            begin
              mem_check[9][16].run()  ;
            end
            begin
              rf_driver[9][16].run()  ;
            end

            begin
              gen[9][17].run()  ;
            end
            begin
              drv[9][17].run()  ;
            end
            begin
              mem_check[9][17].run()  ;
            end
            begin
              rf_driver[9][17].run()  ;
            end

            begin
              gen[9][18].run()  ;
            end
            begin
              drv[9][18].run()  ;
            end
            begin
              mem_check[9][18].run()  ;
            end
            begin
              rf_driver[9][18].run()  ;
            end

            begin
              gen[9][19].run()  ;
            end
            begin
              drv[9][19].run()  ;
            end
            begin
              mem_check[9][19].run()  ;
            end
            begin
              rf_driver[9][19].run()  ;
            end

            begin
              gen[9][20].run()  ;
            end
            begin
              drv[9][20].run()  ;
            end
            begin
              mem_check[9][20].run()  ;
            end
            begin
              rf_driver[9][20].run()  ;
            end

            begin
              gen[9][21].run()  ;
            end
            begin
              drv[9][21].run()  ;
            end
            begin
              mem_check[9][21].run()  ;
            end
            begin
              rf_driver[9][21].run()  ;
            end

            begin
              gen[9][22].run()  ;
            end
            begin
              drv[9][22].run()  ;
            end
            begin
              mem_check[9][22].run()  ;
            end
            begin
              rf_driver[9][22].run()  ;
            end

            begin
              gen[9][23].run()  ;
            end
            begin
              drv[9][23].run()  ;
            end
            begin
              mem_check[9][23].run()  ;
            end
            begin
              rf_driver[9][23].run()  ;
            end

            begin
              gen[9][24].run()  ;
            end
            begin
              drv[9][24].run()  ;
            end
            begin
              mem_check[9][24].run()  ;
            end
            begin
              rf_driver[9][24].run()  ;
            end

            begin
              gen[9][25].run()  ;
            end
            begin
              drv[9][25].run()  ;
            end
            begin
              mem_check[9][25].run()  ;
            end
            begin
              rf_driver[9][25].run()  ;
            end

            begin
              gen[9][26].run()  ;
            end
            begin
              drv[9][26].run()  ;
            end
            begin
              mem_check[9][26].run()  ;
            end
            begin
              rf_driver[9][26].run()  ;
            end

            begin
              gen[9][27].run()  ;
            end
            begin
              drv[9][27].run()  ;
            end
            begin
              mem_check[9][27].run()  ;
            end
            begin
              rf_driver[9][27].run()  ;
            end

            begin
              gen[9][28].run()  ;
            end
            begin
              drv[9][28].run()  ;
            end
            begin
              mem_check[9][28].run()  ;
            end
            begin
              rf_driver[9][28].run()  ;
            end

            begin
              gen[9][29].run()  ;
            end
            begin
              drv[9][29].run()  ;
            end
            begin
              mem_check[9][29].run()  ;
            end
            begin
              rf_driver[9][29].run()  ;
            end

            begin
              gen[9][30].run()  ;
            end
            begin
              drv[9][30].run()  ;
            end
            begin
              mem_check[9][30].run()  ;
            end
            begin
              rf_driver[9][30].run()  ;
            end

            begin
              gen[9][31].run()  ;
            end
            begin
              drv[9][31].run()  ;
            end
            begin
              mem_check[9][31].run()  ;
            end
            begin
              rf_driver[9][31].run()  ;
            end

            begin
              ldst_driver[10].run()  ;
            end
            begin
              mgr[10].run()  ;
            end
            begin
              oob_drv[10].run()  ;
            end
            begin
              up_check[10].run()  ;
            end
            begin
              gen[10][0].run()  ;
            end
            begin
              drv[10][0].run()  ;
            end
            begin
              mem_check[10][0].run()  ;
            end
            begin
              rf_driver[10][0].run()  ;
            end

            begin
              gen[10][1].run()  ;
            end
            begin
              drv[10][1].run()  ;
            end
            begin
              mem_check[10][1].run()  ;
            end
            begin
              rf_driver[10][1].run()  ;
            end

            begin
              gen[10][2].run()  ;
            end
            begin
              drv[10][2].run()  ;
            end
            begin
              mem_check[10][2].run()  ;
            end
            begin
              rf_driver[10][2].run()  ;
            end

            begin
              gen[10][3].run()  ;
            end
            begin
              drv[10][3].run()  ;
            end
            begin
              mem_check[10][3].run()  ;
            end
            begin
              rf_driver[10][3].run()  ;
            end

            begin
              gen[10][4].run()  ;
            end
            begin
              drv[10][4].run()  ;
            end
            begin
              mem_check[10][4].run()  ;
            end
            begin
              rf_driver[10][4].run()  ;
            end

            begin
              gen[10][5].run()  ;
            end
            begin
              drv[10][5].run()  ;
            end
            begin
              mem_check[10][5].run()  ;
            end
            begin
              rf_driver[10][5].run()  ;
            end

            begin
              gen[10][6].run()  ;
            end
            begin
              drv[10][6].run()  ;
            end
            begin
              mem_check[10][6].run()  ;
            end
            begin
              rf_driver[10][6].run()  ;
            end

            begin
              gen[10][7].run()  ;
            end
            begin
              drv[10][7].run()  ;
            end
            begin
              mem_check[10][7].run()  ;
            end
            begin
              rf_driver[10][7].run()  ;
            end

            begin
              gen[10][8].run()  ;
            end
            begin
              drv[10][8].run()  ;
            end
            begin
              mem_check[10][8].run()  ;
            end
            begin
              rf_driver[10][8].run()  ;
            end

            begin
              gen[10][9].run()  ;
            end
            begin
              drv[10][9].run()  ;
            end
            begin
              mem_check[10][9].run()  ;
            end
            begin
              rf_driver[10][9].run()  ;
            end

            begin
              gen[10][10].run()  ;
            end
            begin
              drv[10][10].run()  ;
            end
            begin
              mem_check[10][10].run()  ;
            end
            begin
              rf_driver[10][10].run()  ;
            end

            begin
              gen[10][11].run()  ;
            end
            begin
              drv[10][11].run()  ;
            end
            begin
              mem_check[10][11].run()  ;
            end
            begin
              rf_driver[10][11].run()  ;
            end

            begin
              gen[10][12].run()  ;
            end
            begin
              drv[10][12].run()  ;
            end
            begin
              mem_check[10][12].run()  ;
            end
            begin
              rf_driver[10][12].run()  ;
            end

            begin
              gen[10][13].run()  ;
            end
            begin
              drv[10][13].run()  ;
            end
            begin
              mem_check[10][13].run()  ;
            end
            begin
              rf_driver[10][13].run()  ;
            end

            begin
              gen[10][14].run()  ;
            end
            begin
              drv[10][14].run()  ;
            end
            begin
              mem_check[10][14].run()  ;
            end
            begin
              rf_driver[10][14].run()  ;
            end

            begin
              gen[10][15].run()  ;
            end
            begin
              drv[10][15].run()  ;
            end
            begin
              mem_check[10][15].run()  ;
            end
            begin
              rf_driver[10][15].run()  ;
            end

            begin
              gen[10][16].run()  ;
            end
            begin
              drv[10][16].run()  ;
            end
            begin
              mem_check[10][16].run()  ;
            end
            begin
              rf_driver[10][16].run()  ;
            end

            begin
              gen[10][17].run()  ;
            end
            begin
              drv[10][17].run()  ;
            end
            begin
              mem_check[10][17].run()  ;
            end
            begin
              rf_driver[10][17].run()  ;
            end

            begin
              gen[10][18].run()  ;
            end
            begin
              drv[10][18].run()  ;
            end
            begin
              mem_check[10][18].run()  ;
            end
            begin
              rf_driver[10][18].run()  ;
            end

            begin
              gen[10][19].run()  ;
            end
            begin
              drv[10][19].run()  ;
            end
            begin
              mem_check[10][19].run()  ;
            end
            begin
              rf_driver[10][19].run()  ;
            end

            begin
              gen[10][20].run()  ;
            end
            begin
              drv[10][20].run()  ;
            end
            begin
              mem_check[10][20].run()  ;
            end
            begin
              rf_driver[10][20].run()  ;
            end

            begin
              gen[10][21].run()  ;
            end
            begin
              drv[10][21].run()  ;
            end
            begin
              mem_check[10][21].run()  ;
            end
            begin
              rf_driver[10][21].run()  ;
            end

            begin
              gen[10][22].run()  ;
            end
            begin
              drv[10][22].run()  ;
            end
            begin
              mem_check[10][22].run()  ;
            end
            begin
              rf_driver[10][22].run()  ;
            end

            begin
              gen[10][23].run()  ;
            end
            begin
              drv[10][23].run()  ;
            end
            begin
              mem_check[10][23].run()  ;
            end
            begin
              rf_driver[10][23].run()  ;
            end

            begin
              gen[10][24].run()  ;
            end
            begin
              drv[10][24].run()  ;
            end
            begin
              mem_check[10][24].run()  ;
            end
            begin
              rf_driver[10][24].run()  ;
            end

            begin
              gen[10][25].run()  ;
            end
            begin
              drv[10][25].run()  ;
            end
            begin
              mem_check[10][25].run()  ;
            end
            begin
              rf_driver[10][25].run()  ;
            end

            begin
              gen[10][26].run()  ;
            end
            begin
              drv[10][26].run()  ;
            end
            begin
              mem_check[10][26].run()  ;
            end
            begin
              rf_driver[10][26].run()  ;
            end

            begin
              gen[10][27].run()  ;
            end
            begin
              drv[10][27].run()  ;
            end
            begin
              mem_check[10][27].run()  ;
            end
            begin
              rf_driver[10][27].run()  ;
            end

            begin
              gen[10][28].run()  ;
            end
            begin
              drv[10][28].run()  ;
            end
            begin
              mem_check[10][28].run()  ;
            end
            begin
              rf_driver[10][28].run()  ;
            end

            begin
              gen[10][29].run()  ;
            end
            begin
              drv[10][29].run()  ;
            end
            begin
              mem_check[10][29].run()  ;
            end
            begin
              rf_driver[10][29].run()  ;
            end

            begin
              gen[10][30].run()  ;
            end
            begin
              drv[10][30].run()  ;
            end
            begin
              mem_check[10][30].run()  ;
            end
            begin
              rf_driver[10][30].run()  ;
            end

            begin
              gen[10][31].run()  ;
            end
            begin
              drv[10][31].run()  ;
            end
            begin
              mem_check[10][31].run()  ;
            end
            begin
              rf_driver[10][31].run()  ;
            end

            begin
              ldst_driver[11].run()  ;
            end
            begin
              mgr[11].run()  ;
            end
            begin
              oob_drv[11].run()  ;
            end
            begin
              up_check[11].run()  ;
            end
            begin
              gen[11][0].run()  ;
            end
            begin
              drv[11][0].run()  ;
            end
            begin
              mem_check[11][0].run()  ;
            end
            begin
              rf_driver[11][0].run()  ;
            end

            begin
              gen[11][1].run()  ;
            end
            begin
              drv[11][1].run()  ;
            end
            begin
              mem_check[11][1].run()  ;
            end
            begin
              rf_driver[11][1].run()  ;
            end

            begin
              gen[11][2].run()  ;
            end
            begin
              drv[11][2].run()  ;
            end
            begin
              mem_check[11][2].run()  ;
            end
            begin
              rf_driver[11][2].run()  ;
            end

            begin
              gen[11][3].run()  ;
            end
            begin
              drv[11][3].run()  ;
            end
            begin
              mem_check[11][3].run()  ;
            end
            begin
              rf_driver[11][3].run()  ;
            end

            begin
              gen[11][4].run()  ;
            end
            begin
              drv[11][4].run()  ;
            end
            begin
              mem_check[11][4].run()  ;
            end
            begin
              rf_driver[11][4].run()  ;
            end

            begin
              gen[11][5].run()  ;
            end
            begin
              drv[11][5].run()  ;
            end
            begin
              mem_check[11][5].run()  ;
            end
            begin
              rf_driver[11][5].run()  ;
            end

            begin
              gen[11][6].run()  ;
            end
            begin
              drv[11][6].run()  ;
            end
            begin
              mem_check[11][6].run()  ;
            end
            begin
              rf_driver[11][6].run()  ;
            end

            begin
              gen[11][7].run()  ;
            end
            begin
              drv[11][7].run()  ;
            end
            begin
              mem_check[11][7].run()  ;
            end
            begin
              rf_driver[11][7].run()  ;
            end

            begin
              gen[11][8].run()  ;
            end
            begin
              drv[11][8].run()  ;
            end
            begin
              mem_check[11][8].run()  ;
            end
            begin
              rf_driver[11][8].run()  ;
            end

            begin
              gen[11][9].run()  ;
            end
            begin
              drv[11][9].run()  ;
            end
            begin
              mem_check[11][9].run()  ;
            end
            begin
              rf_driver[11][9].run()  ;
            end

            begin
              gen[11][10].run()  ;
            end
            begin
              drv[11][10].run()  ;
            end
            begin
              mem_check[11][10].run()  ;
            end
            begin
              rf_driver[11][10].run()  ;
            end

            begin
              gen[11][11].run()  ;
            end
            begin
              drv[11][11].run()  ;
            end
            begin
              mem_check[11][11].run()  ;
            end
            begin
              rf_driver[11][11].run()  ;
            end

            begin
              gen[11][12].run()  ;
            end
            begin
              drv[11][12].run()  ;
            end
            begin
              mem_check[11][12].run()  ;
            end
            begin
              rf_driver[11][12].run()  ;
            end

            begin
              gen[11][13].run()  ;
            end
            begin
              drv[11][13].run()  ;
            end
            begin
              mem_check[11][13].run()  ;
            end
            begin
              rf_driver[11][13].run()  ;
            end

            begin
              gen[11][14].run()  ;
            end
            begin
              drv[11][14].run()  ;
            end
            begin
              mem_check[11][14].run()  ;
            end
            begin
              rf_driver[11][14].run()  ;
            end

            begin
              gen[11][15].run()  ;
            end
            begin
              drv[11][15].run()  ;
            end
            begin
              mem_check[11][15].run()  ;
            end
            begin
              rf_driver[11][15].run()  ;
            end

            begin
              gen[11][16].run()  ;
            end
            begin
              drv[11][16].run()  ;
            end
            begin
              mem_check[11][16].run()  ;
            end
            begin
              rf_driver[11][16].run()  ;
            end

            begin
              gen[11][17].run()  ;
            end
            begin
              drv[11][17].run()  ;
            end
            begin
              mem_check[11][17].run()  ;
            end
            begin
              rf_driver[11][17].run()  ;
            end

            begin
              gen[11][18].run()  ;
            end
            begin
              drv[11][18].run()  ;
            end
            begin
              mem_check[11][18].run()  ;
            end
            begin
              rf_driver[11][18].run()  ;
            end

            begin
              gen[11][19].run()  ;
            end
            begin
              drv[11][19].run()  ;
            end
            begin
              mem_check[11][19].run()  ;
            end
            begin
              rf_driver[11][19].run()  ;
            end

            begin
              gen[11][20].run()  ;
            end
            begin
              drv[11][20].run()  ;
            end
            begin
              mem_check[11][20].run()  ;
            end
            begin
              rf_driver[11][20].run()  ;
            end

            begin
              gen[11][21].run()  ;
            end
            begin
              drv[11][21].run()  ;
            end
            begin
              mem_check[11][21].run()  ;
            end
            begin
              rf_driver[11][21].run()  ;
            end

            begin
              gen[11][22].run()  ;
            end
            begin
              drv[11][22].run()  ;
            end
            begin
              mem_check[11][22].run()  ;
            end
            begin
              rf_driver[11][22].run()  ;
            end

            begin
              gen[11][23].run()  ;
            end
            begin
              drv[11][23].run()  ;
            end
            begin
              mem_check[11][23].run()  ;
            end
            begin
              rf_driver[11][23].run()  ;
            end

            begin
              gen[11][24].run()  ;
            end
            begin
              drv[11][24].run()  ;
            end
            begin
              mem_check[11][24].run()  ;
            end
            begin
              rf_driver[11][24].run()  ;
            end

            begin
              gen[11][25].run()  ;
            end
            begin
              drv[11][25].run()  ;
            end
            begin
              mem_check[11][25].run()  ;
            end
            begin
              rf_driver[11][25].run()  ;
            end

            begin
              gen[11][26].run()  ;
            end
            begin
              drv[11][26].run()  ;
            end
            begin
              mem_check[11][26].run()  ;
            end
            begin
              rf_driver[11][26].run()  ;
            end

            begin
              gen[11][27].run()  ;
            end
            begin
              drv[11][27].run()  ;
            end
            begin
              mem_check[11][27].run()  ;
            end
            begin
              rf_driver[11][27].run()  ;
            end

            begin
              gen[11][28].run()  ;
            end
            begin
              drv[11][28].run()  ;
            end
            begin
              mem_check[11][28].run()  ;
            end
            begin
              rf_driver[11][28].run()  ;
            end

            begin
              gen[11][29].run()  ;
            end
            begin
              drv[11][29].run()  ;
            end
            begin
              mem_check[11][29].run()  ;
            end
            begin
              rf_driver[11][29].run()  ;
            end

            begin
              gen[11][30].run()  ;
            end
            begin
              drv[11][30].run()  ;
            end
            begin
              mem_check[11][30].run()  ;
            end
            begin
              rf_driver[11][30].run()  ;
            end

            begin
              gen[11][31].run()  ;
            end
            begin
              drv[11][31].run()  ;
            end
            begin
              mem_check[11][31].run()  ;
            end
            begin
              rf_driver[11][31].run()  ;
            end

            begin
              ldst_driver[12].run()  ;
            end
            begin
              mgr[12].run()  ;
            end
            begin
              oob_drv[12].run()  ;
            end
            begin
              up_check[12].run()  ;
            end
            begin
              gen[12][0].run()  ;
            end
            begin
              drv[12][0].run()  ;
            end
            begin
              mem_check[12][0].run()  ;
            end
            begin
              rf_driver[12][0].run()  ;
            end

            begin
              gen[12][1].run()  ;
            end
            begin
              drv[12][1].run()  ;
            end
            begin
              mem_check[12][1].run()  ;
            end
            begin
              rf_driver[12][1].run()  ;
            end

            begin
              gen[12][2].run()  ;
            end
            begin
              drv[12][2].run()  ;
            end
            begin
              mem_check[12][2].run()  ;
            end
            begin
              rf_driver[12][2].run()  ;
            end

            begin
              gen[12][3].run()  ;
            end
            begin
              drv[12][3].run()  ;
            end
            begin
              mem_check[12][3].run()  ;
            end
            begin
              rf_driver[12][3].run()  ;
            end

            begin
              gen[12][4].run()  ;
            end
            begin
              drv[12][4].run()  ;
            end
            begin
              mem_check[12][4].run()  ;
            end
            begin
              rf_driver[12][4].run()  ;
            end

            begin
              gen[12][5].run()  ;
            end
            begin
              drv[12][5].run()  ;
            end
            begin
              mem_check[12][5].run()  ;
            end
            begin
              rf_driver[12][5].run()  ;
            end

            begin
              gen[12][6].run()  ;
            end
            begin
              drv[12][6].run()  ;
            end
            begin
              mem_check[12][6].run()  ;
            end
            begin
              rf_driver[12][6].run()  ;
            end

            begin
              gen[12][7].run()  ;
            end
            begin
              drv[12][7].run()  ;
            end
            begin
              mem_check[12][7].run()  ;
            end
            begin
              rf_driver[12][7].run()  ;
            end

            begin
              gen[12][8].run()  ;
            end
            begin
              drv[12][8].run()  ;
            end
            begin
              mem_check[12][8].run()  ;
            end
            begin
              rf_driver[12][8].run()  ;
            end

            begin
              gen[12][9].run()  ;
            end
            begin
              drv[12][9].run()  ;
            end
            begin
              mem_check[12][9].run()  ;
            end
            begin
              rf_driver[12][9].run()  ;
            end

            begin
              gen[12][10].run()  ;
            end
            begin
              drv[12][10].run()  ;
            end
            begin
              mem_check[12][10].run()  ;
            end
            begin
              rf_driver[12][10].run()  ;
            end

            begin
              gen[12][11].run()  ;
            end
            begin
              drv[12][11].run()  ;
            end
            begin
              mem_check[12][11].run()  ;
            end
            begin
              rf_driver[12][11].run()  ;
            end

            begin
              gen[12][12].run()  ;
            end
            begin
              drv[12][12].run()  ;
            end
            begin
              mem_check[12][12].run()  ;
            end
            begin
              rf_driver[12][12].run()  ;
            end

            begin
              gen[12][13].run()  ;
            end
            begin
              drv[12][13].run()  ;
            end
            begin
              mem_check[12][13].run()  ;
            end
            begin
              rf_driver[12][13].run()  ;
            end

            begin
              gen[12][14].run()  ;
            end
            begin
              drv[12][14].run()  ;
            end
            begin
              mem_check[12][14].run()  ;
            end
            begin
              rf_driver[12][14].run()  ;
            end

            begin
              gen[12][15].run()  ;
            end
            begin
              drv[12][15].run()  ;
            end
            begin
              mem_check[12][15].run()  ;
            end
            begin
              rf_driver[12][15].run()  ;
            end

            begin
              gen[12][16].run()  ;
            end
            begin
              drv[12][16].run()  ;
            end
            begin
              mem_check[12][16].run()  ;
            end
            begin
              rf_driver[12][16].run()  ;
            end

            begin
              gen[12][17].run()  ;
            end
            begin
              drv[12][17].run()  ;
            end
            begin
              mem_check[12][17].run()  ;
            end
            begin
              rf_driver[12][17].run()  ;
            end

            begin
              gen[12][18].run()  ;
            end
            begin
              drv[12][18].run()  ;
            end
            begin
              mem_check[12][18].run()  ;
            end
            begin
              rf_driver[12][18].run()  ;
            end

            begin
              gen[12][19].run()  ;
            end
            begin
              drv[12][19].run()  ;
            end
            begin
              mem_check[12][19].run()  ;
            end
            begin
              rf_driver[12][19].run()  ;
            end

            begin
              gen[12][20].run()  ;
            end
            begin
              drv[12][20].run()  ;
            end
            begin
              mem_check[12][20].run()  ;
            end
            begin
              rf_driver[12][20].run()  ;
            end

            begin
              gen[12][21].run()  ;
            end
            begin
              drv[12][21].run()  ;
            end
            begin
              mem_check[12][21].run()  ;
            end
            begin
              rf_driver[12][21].run()  ;
            end

            begin
              gen[12][22].run()  ;
            end
            begin
              drv[12][22].run()  ;
            end
            begin
              mem_check[12][22].run()  ;
            end
            begin
              rf_driver[12][22].run()  ;
            end

            begin
              gen[12][23].run()  ;
            end
            begin
              drv[12][23].run()  ;
            end
            begin
              mem_check[12][23].run()  ;
            end
            begin
              rf_driver[12][23].run()  ;
            end

            begin
              gen[12][24].run()  ;
            end
            begin
              drv[12][24].run()  ;
            end
            begin
              mem_check[12][24].run()  ;
            end
            begin
              rf_driver[12][24].run()  ;
            end

            begin
              gen[12][25].run()  ;
            end
            begin
              drv[12][25].run()  ;
            end
            begin
              mem_check[12][25].run()  ;
            end
            begin
              rf_driver[12][25].run()  ;
            end

            begin
              gen[12][26].run()  ;
            end
            begin
              drv[12][26].run()  ;
            end
            begin
              mem_check[12][26].run()  ;
            end
            begin
              rf_driver[12][26].run()  ;
            end

            begin
              gen[12][27].run()  ;
            end
            begin
              drv[12][27].run()  ;
            end
            begin
              mem_check[12][27].run()  ;
            end
            begin
              rf_driver[12][27].run()  ;
            end

            begin
              gen[12][28].run()  ;
            end
            begin
              drv[12][28].run()  ;
            end
            begin
              mem_check[12][28].run()  ;
            end
            begin
              rf_driver[12][28].run()  ;
            end

            begin
              gen[12][29].run()  ;
            end
            begin
              drv[12][29].run()  ;
            end
            begin
              mem_check[12][29].run()  ;
            end
            begin
              rf_driver[12][29].run()  ;
            end

            begin
              gen[12][30].run()  ;
            end
            begin
              drv[12][30].run()  ;
            end
            begin
              mem_check[12][30].run()  ;
            end
            begin
              rf_driver[12][30].run()  ;
            end

            begin
              gen[12][31].run()  ;
            end
            begin
              drv[12][31].run()  ;
            end
            begin
              mem_check[12][31].run()  ;
            end
            begin
              rf_driver[12][31].run()  ;
            end

            begin
              ldst_driver[13].run()  ;
            end
            begin
              mgr[13].run()  ;
            end
            begin
              oob_drv[13].run()  ;
            end
            begin
              up_check[13].run()  ;
            end
            begin
              gen[13][0].run()  ;
            end
            begin
              drv[13][0].run()  ;
            end
            begin
              mem_check[13][0].run()  ;
            end
            begin
              rf_driver[13][0].run()  ;
            end

            begin
              gen[13][1].run()  ;
            end
            begin
              drv[13][1].run()  ;
            end
            begin
              mem_check[13][1].run()  ;
            end
            begin
              rf_driver[13][1].run()  ;
            end

            begin
              gen[13][2].run()  ;
            end
            begin
              drv[13][2].run()  ;
            end
            begin
              mem_check[13][2].run()  ;
            end
            begin
              rf_driver[13][2].run()  ;
            end

            begin
              gen[13][3].run()  ;
            end
            begin
              drv[13][3].run()  ;
            end
            begin
              mem_check[13][3].run()  ;
            end
            begin
              rf_driver[13][3].run()  ;
            end

            begin
              gen[13][4].run()  ;
            end
            begin
              drv[13][4].run()  ;
            end
            begin
              mem_check[13][4].run()  ;
            end
            begin
              rf_driver[13][4].run()  ;
            end

            begin
              gen[13][5].run()  ;
            end
            begin
              drv[13][5].run()  ;
            end
            begin
              mem_check[13][5].run()  ;
            end
            begin
              rf_driver[13][5].run()  ;
            end

            begin
              gen[13][6].run()  ;
            end
            begin
              drv[13][6].run()  ;
            end
            begin
              mem_check[13][6].run()  ;
            end
            begin
              rf_driver[13][6].run()  ;
            end

            begin
              gen[13][7].run()  ;
            end
            begin
              drv[13][7].run()  ;
            end
            begin
              mem_check[13][7].run()  ;
            end
            begin
              rf_driver[13][7].run()  ;
            end

            begin
              gen[13][8].run()  ;
            end
            begin
              drv[13][8].run()  ;
            end
            begin
              mem_check[13][8].run()  ;
            end
            begin
              rf_driver[13][8].run()  ;
            end

            begin
              gen[13][9].run()  ;
            end
            begin
              drv[13][9].run()  ;
            end
            begin
              mem_check[13][9].run()  ;
            end
            begin
              rf_driver[13][9].run()  ;
            end

            begin
              gen[13][10].run()  ;
            end
            begin
              drv[13][10].run()  ;
            end
            begin
              mem_check[13][10].run()  ;
            end
            begin
              rf_driver[13][10].run()  ;
            end

            begin
              gen[13][11].run()  ;
            end
            begin
              drv[13][11].run()  ;
            end
            begin
              mem_check[13][11].run()  ;
            end
            begin
              rf_driver[13][11].run()  ;
            end

            begin
              gen[13][12].run()  ;
            end
            begin
              drv[13][12].run()  ;
            end
            begin
              mem_check[13][12].run()  ;
            end
            begin
              rf_driver[13][12].run()  ;
            end

            begin
              gen[13][13].run()  ;
            end
            begin
              drv[13][13].run()  ;
            end
            begin
              mem_check[13][13].run()  ;
            end
            begin
              rf_driver[13][13].run()  ;
            end

            begin
              gen[13][14].run()  ;
            end
            begin
              drv[13][14].run()  ;
            end
            begin
              mem_check[13][14].run()  ;
            end
            begin
              rf_driver[13][14].run()  ;
            end

            begin
              gen[13][15].run()  ;
            end
            begin
              drv[13][15].run()  ;
            end
            begin
              mem_check[13][15].run()  ;
            end
            begin
              rf_driver[13][15].run()  ;
            end

            begin
              gen[13][16].run()  ;
            end
            begin
              drv[13][16].run()  ;
            end
            begin
              mem_check[13][16].run()  ;
            end
            begin
              rf_driver[13][16].run()  ;
            end

            begin
              gen[13][17].run()  ;
            end
            begin
              drv[13][17].run()  ;
            end
            begin
              mem_check[13][17].run()  ;
            end
            begin
              rf_driver[13][17].run()  ;
            end

            begin
              gen[13][18].run()  ;
            end
            begin
              drv[13][18].run()  ;
            end
            begin
              mem_check[13][18].run()  ;
            end
            begin
              rf_driver[13][18].run()  ;
            end

            begin
              gen[13][19].run()  ;
            end
            begin
              drv[13][19].run()  ;
            end
            begin
              mem_check[13][19].run()  ;
            end
            begin
              rf_driver[13][19].run()  ;
            end

            begin
              gen[13][20].run()  ;
            end
            begin
              drv[13][20].run()  ;
            end
            begin
              mem_check[13][20].run()  ;
            end
            begin
              rf_driver[13][20].run()  ;
            end

            begin
              gen[13][21].run()  ;
            end
            begin
              drv[13][21].run()  ;
            end
            begin
              mem_check[13][21].run()  ;
            end
            begin
              rf_driver[13][21].run()  ;
            end

            begin
              gen[13][22].run()  ;
            end
            begin
              drv[13][22].run()  ;
            end
            begin
              mem_check[13][22].run()  ;
            end
            begin
              rf_driver[13][22].run()  ;
            end

            begin
              gen[13][23].run()  ;
            end
            begin
              drv[13][23].run()  ;
            end
            begin
              mem_check[13][23].run()  ;
            end
            begin
              rf_driver[13][23].run()  ;
            end

            begin
              gen[13][24].run()  ;
            end
            begin
              drv[13][24].run()  ;
            end
            begin
              mem_check[13][24].run()  ;
            end
            begin
              rf_driver[13][24].run()  ;
            end

            begin
              gen[13][25].run()  ;
            end
            begin
              drv[13][25].run()  ;
            end
            begin
              mem_check[13][25].run()  ;
            end
            begin
              rf_driver[13][25].run()  ;
            end

            begin
              gen[13][26].run()  ;
            end
            begin
              drv[13][26].run()  ;
            end
            begin
              mem_check[13][26].run()  ;
            end
            begin
              rf_driver[13][26].run()  ;
            end

            begin
              gen[13][27].run()  ;
            end
            begin
              drv[13][27].run()  ;
            end
            begin
              mem_check[13][27].run()  ;
            end
            begin
              rf_driver[13][27].run()  ;
            end

            begin
              gen[13][28].run()  ;
            end
            begin
              drv[13][28].run()  ;
            end
            begin
              mem_check[13][28].run()  ;
            end
            begin
              rf_driver[13][28].run()  ;
            end

            begin
              gen[13][29].run()  ;
            end
            begin
              drv[13][29].run()  ;
            end
            begin
              mem_check[13][29].run()  ;
            end
            begin
              rf_driver[13][29].run()  ;
            end

            begin
              gen[13][30].run()  ;
            end
            begin
              drv[13][30].run()  ;
            end
            begin
              mem_check[13][30].run()  ;
            end
            begin
              rf_driver[13][30].run()  ;
            end

            begin
              gen[13][31].run()  ;
            end
            begin
              drv[13][31].run()  ;
            end
            begin
              mem_check[13][31].run()  ;
            end
            begin
              rf_driver[13][31].run()  ;
            end

            begin
              ldst_driver[14].run()  ;
            end
            begin
              mgr[14].run()  ;
            end
            begin
              oob_drv[14].run()  ;
            end
            begin
              up_check[14].run()  ;
            end
            begin
              gen[14][0].run()  ;
            end
            begin
              drv[14][0].run()  ;
            end
            begin
              mem_check[14][0].run()  ;
            end
            begin
              rf_driver[14][0].run()  ;
            end

            begin
              gen[14][1].run()  ;
            end
            begin
              drv[14][1].run()  ;
            end
            begin
              mem_check[14][1].run()  ;
            end
            begin
              rf_driver[14][1].run()  ;
            end

            begin
              gen[14][2].run()  ;
            end
            begin
              drv[14][2].run()  ;
            end
            begin
              mem_check[14][2].run()  ;
            end
            begin
              rf_driver[14][2].run()  ;
            end

            begin
              gen[14][3].run()  ;
            end
            begin
              drv[14][3].run()  ;
            end
            begin
              mem_check[14][3].run()  ;
            end
            begin
              rf_driver[14][3].run()  ;
            end

            begin
              gen[14][4].run()  ;
            end
            begin
              drv[14][4].run()  ;
            end
            begin
              mem_check[14][4].run()  ;
            end
            begin
              rf_driver[14][4].run()  ;
            end

            begin
              gen[14][5].run()  ;
            end
            begin
              drv[14][5].run()  ;
            end
            begin
              mem_check[14][5].run()  ;
            end
            begin
              rf_driver[14][5].run()  ;
            end

            begin
              gen[14][6].run()  ;
            end
            begin
              drv[14][6].run()  ;
            end
            begin
              mem_check[14][6].run()  ;
            end
            begin
              rf_driver[14][6].run()  ;
            end

            begin
              gen[14][7].run()  ;
            end
            begin
              drv[14][7].run()  ;
            end
            begin
              mem_check[14][7].run()  ;
            end
            begin
              rf_driver[14][7].run()  ;
            end

            begin
              gen[14][8].run()  ;
            end
            begin
              drv[14][8].run()  ;
            end
            begin
              mem_check[14][8].run()  ;
            end
            begin
              rf_driver[14][8].run()  ;
            end

            begin
              gen[14][9].run()  ;
            end
            begin
              drv[14][9].run()  ;
            end
            begin
              mem_check[14][9].run()  ;
            end
            begin
              rf_driver[14][9].run()  ;
            end

            begin
              gen[14][10].run()  ;
            end
            begin
              drv[14][10].run()  ;
            end
            begin
              mem_check[14][10].run()  ;
            end
            begin
              rf_driver[14][10].run()  ;
            end

            begin
              gen[14][11].run()  ;
            end
            begin
              drv[14][11].run()  ;
            end
            begin
              mem_check[14][11].run()  ;
            end
            begin
              rf_driver[14][11].run()  ;
            end

            begin
              gen[14][12].run()  ;
            end
            begin
              drv[14][12].run()  ;
            end
            begin
              mem_check[14][12].run()  ;
            end
            begin
              rf_driver[14][12].run()  ;
            end

            begin
              gen[14][13].run()  ;
            end
            begin
              drv[14][13].run()  ;
            end
            begin
              mem_check[14][13].run()  ;
            end
            begin
              rf_driver[14][13].run()  ;
            end

            begin
              gen[14][14].run()  ;
            end
            begin
              drv[14][14].run()  ;
            end
            begin
              mem_check[14][14].run()  ;
            end
            begin
              rf_driver[14][14].run()  ;
            end

            begin
              gen[14][15].run()  ;
            end
            begin
              drv[14][15].run()  ;
            end
            begin
              mem_check[14][15].run()  ;
            end
            begin
              rf_driver[14][15].run()  ;
            end

            begin
              gen[14][16].run()  ;
            end
            begin
              drv[14][16].run()  ;
            end
            begin
              mem_check[14][16].run()  ;
            end
            begin
              rf_driver[14][16].run()  ;
            end

            begin
              gen[14][17].run()  ;
            end
            begin
              drv[14][17].run()  ;
            end
            begin
              mem_check[14][17].run()  ;
            end
            begin
              rf_driver[14][17].run()  ;
            end

            begin
              gen[14][18].run()  ;
            end
            begin
              drv[14][18].run()  ;
            end
            begin
              mem_check[14][18].run()  ;
            end
            begin
              rf_driver[14][18].run()  ;
            end

            begin
              gen[14][19].run()  ;
            end
            begin
              drv[14][19].run()  ;
            end
            begin
              mem_check[14][19].run()  ;
            end
            begin
              rf_driver[14][19].run()  ;
            end

            begin
              gen[14][20].run()  ;
            end
            begin
              drv[14][20].run()  ;
            end
            begin
              mem_check[14][20].run()  ;
            end
            begin
              rf_driver[14][20].run()  ;
            end

            begin
              gen[14][21].run()  ;
            end
            begin
              drv[14][21].run()  ;
            end
            begin
              mem_check[14][21].run()  ;
            end
            begin
              rf_driver[14][21].run()  ;
            end

            begin
              gen[14][22].run()  ;
            end
            begin
              drv[14][22].run()  ;
            end
            begin
              mem_check[14][22].run()  ;
            end
            begin
              rf_driver[14][22].run()  ;
            end

            begin
              gen[14][23].run()  ;
            end
            begin
              drv[14][23].run()  ;
            end
            begin
              mem_check[14][23].run()  ;
            end
            begin
              rf_driver[14][23].run()  ;
            end

            begin
              gen[14][24].run()  ;
            end
            begin
              drv[14][24].run()  ;
            end
            begin
              mem_check[14][24].run()  ;
            end
            begin
              rf_driver[14][24].run()  ;
            end

            begin
              gen[14][25].run()  ;
            end
            begin
              drv[14][25].run()  ;
            end
            begin
              mem_check[14][25].run()  ;
            end
            begin
              rf_driver[14][25].run()  ;
            end

            begin
              gen[14][26].run()  ;
            end
            begin
              drv[14][26].run()  ;
            end
            begin
              mem_check[14][26].run()  ;
            end
            begin
              rf_driver[14][26].run()  ;
            end

            begin
              gen[14][27].run()  ;
            end
            begin
              drv[14][27].run()  ;
            end
            begin
              mem_check[14][27].run()  ;
            end
            begin
              rf_driver[14][27].run()  ;
            end

            begin
              gen[14][28].run()  ;
            end
            begin
              drv[14][28].run()  ;
            end
            begin
              mem_check[14][28].run()  ;
            end
            begin
              rf_driver[14][28].run()  ;
            end

            begin
              gen[14][29].run()  ;
            end
            begin
              drv[14][29].run()  ;
            end
            begin
              mem_check[14][29].run()  ;
            end
            begin
              rf_driver[14][29].run()  ;
            end

            begin
              gen[14][30].run()  ;
            end
            begin
              drv[14][30].run()  ;
            end
            begin
              mem_check[14][30].run()  ;
            end
            begin
              rf_driver[14][30].run()  ;
            end

            begin
              gen[14][31].run()  ;
            end
            begin
              drv[14][31].run()  ;
            end
            begin
              mem_check[14][31].run()  ;
            end
            begin
              rf_driver[14][31].run()  ;
            end

            begin
              ldst_driver[15].run()  ;
            end
            begin
              mgr[15].run()  ;
            end
            begin
              oob_drv[15].run()  ;
            end
            begin
              up_check[15].run()  ;
            end
            begin
              gen[15][0].run()  ;
            end
            begin
              drv[15][0].run()  ;
            end
            begin
              mem_check[15][0].run()  ;
            end
            begin
              rf_driver[15][0].run()  ;
            end

            begin
              gen[15][1].run()  ;
            end
            begin
              drv[15][1].run()  ;
            end
            begin
              mem_check[15][1].run()  ;
            end
            begin
              rf_driver[15][1].run()  ;
            end

            begin
              gen[15][2].run()  ;
            end
            begin
              drv[15][2].run()  ;
            end
            begin
              mem_check[15][2].run()  ;
            end
            begin
              rf_driver[15][2].run()  ;
            end

            begin
              gen[15][3].run()  ;
            end
            begin
              drv[15][3].run()  ;
            end
            begin
              mem_check[15][3].run()  ;
            end
            begin
              rf_driver[15][3].run()  ;
            end

            begin
              gen[15][4].run()  ;
            end
            begin
              drv[15][4].run()  ;
            end
            begin
              mem_check[15][4].run()  ;
            end
            begin
              rf_driver[15][4].run()  ;
            end

            begin
              gen[15][5].run()  ;
            end
            begin
              drv[15][5].run()  ;
            end
            begin
              mem_check[15][5].run()  ;
            end
            begin
              rf_driver[15][5].run()  ;
            end

            begin
              gen[15][6].run()  ;
            end
            begin
              drv[15][6].run()  ;
            end
            begin
              mem_check[15][6].run()  ;
            end
            begin
              rf_driver[15][6].run()  ;
            end

            begin
              gen[15][7].run()  ;
            end
            begin
              drv[15][7].run()  ;
            end
            begin
              mem_check[15][7].run()  ;
            end
            begin
              rf_driver[15][7].run()  ;
            end

            begin
              gen[15][8].run()  ;
            end
            begin
              drv[15][8].run()  ;
            end
            begin
              mem_check[15][8].run()  ;
            end
            begin
              rf_driver[15][8].run()  ;
            end

            begin
              gen[15][9].run()  ;
            end
            begin
              drv[15][9].run()  ;
            end
            begin
              mem_check[15][9].run()  ;
            end
            begin
              rf_driver[15][9].run()  ;
            end

            begin
              gen[15][10].run()  ;
            end
            begin
              drv[15][10].run()  ;
            end
            begin
              mem_check[15][10].run()  ;
            end
            begin
              rf_driver[15][10].run()  ;
            end

            begin
              gen[15][11].run()  ;
            end
            begin
              drv[15][11].run()  ;
            end
            begin
              mem_check[15][11].run()  ;
            end
            begin
              rf_driver[15][11].run()  ;
            end

            begin
              gen[15][12].run()  ;
            end
            begin
              drv[15][12].run()  ;
            end
            begin
              mem_check[15][12].run()  ;
            end
            begin
              rf_driver[15][12].run()  ;
            end

            begin
              gen[15][13].run()  ;
            end
            begin
              drv[15][13].run()  ;
            end
            begin
              mem_check[15][13].run()  ;
            end
            begin
              rf_driver[15][13].run()  ;
            end

            begin
              gen[15][14].run()  ;
            end
            begin
              drv[15][14].run()  ;
            end
            begin
              mem_check[15][14].run()  ;
            end
            begin
              rf_driver[15][14].run()  ;
            end

            begin
              gen[15][15].run()  ;
            end
            begin
              drv[15][15].run()  ;
            end
            begin
              mem_check[15][15].run()  ;
            end
            begin
              rf_driver[15][15].run()  ;
            end

            begin
              gen[15][16].run()  ;
            end
            begin
              drv[15][16].run()  ;
            end
            begin
              mem_check[15][16].run()  ;
            end
            begin
              rf_driver[15][16].run()  ;
            end

            begin
              gen[15][17].run()  ;
            end
            begin
              drv[15][17].run()  ;
            end
            begin
              mem_check[15][17].run()  ;
            end
            begin
              rf_driver[15][17].run()  ;
            end

            begin
              gen[15][18].run()  ;
            end
            begin
              drv[15][18].run()  ;
            end
            begin
              mem_check[15][18].run()  ;
            end
            begin
              rf_driver[15][18].run()  ;
            end

            begin
              gen[15][19].run()  ;
            end
            begin
              drv[15][19].run()  ;
            end
            begin
              mem_check[15][19].run()  ;
            end
            begin
              rf_driver[15][19].run()  ;
            end

            begin
              gen[15][20].run()  ;
            end
            begin
              drv[15][20].run()  ;
            end
            begin
              mem_check[15][20].run()  ;
            end
            begin
              rf_driver[15][20].run()  ;
            end

            begin
              gen[15][21].run()  ;
            end
            begin
              drv[15][21].run()  ;
            end
            begin
              mem_check[15][21].run()  ;
            end
            begin
              rf_driver[15][21].run()  ;
            end

            begin
              gen[15][22].run()  ;
            end
            begin
              drv[15][22].run()  ;
            end
            begin
              mem_check[15][22].run()  ;
            end
            begin
              rf_driver[15][22].run()  ;
            end

            begin
              gen[15][23].run()  ;
            end
            begin
              drv[15][23].run()  ;
            end
            begin
              mem_check[15][23].run()  ;
            end
            begin
              rf_driver[15][23].run()  ;
            end

            begin
              gen[15][24].run()  ;
            end
            begin
              drv[15][24].run()  ;
            end
            begin
              mem_check[15][24].run()  ;
            end
            begin
              rf_driver[15][24].run()  ;
            end

            begin
              gen[15][25].run()  ;
            end
            begin
              drv[15][25].run()  ;
            end
            begin
              mem_check[15][25].run()  ;
            end
            begin
              rf_driver[15][25].run()  ;
            end

            begin
              gen[15][26].run()  ;
            end
            begin
              drv[15][26].run()  ;
            end
            begin
              mem_check[15][26].run()  ;
            end
            begin
              rf_driver[15][26].run()  ;
            end

            begin
              gen[15][27].run()  ;
            end
            begin
              drv[15][27].run()  ;
            end
            begin
              mem_check[15][27].run()  ;
            end
            begin
              rf_driver[15][27].run()  ;
            end

            begin
              gen[15][28].run()  ;
            end
            begin
              drv[15][28].run()  ;
            end
            begin
              mem_check[15][28].run()  ;
            end
            begin
              rf_driver[15][28].run()  ;
            end

            begin
              gen[15][29].run()  ;
            end
            begin
              drv[15][29].run()  ;
            end
            begin
              mem_check[15][29].run()  ;
            end
            begin
              rf_driver[15][29].run()  ;
            end

            begin
              gen[15][30].run()  ;
            end
            begin
              drv[15][30].run()  ;
            end
            begin
              mem_check[15][30].run()  ;
            end
            begin
              rf_driver[15][30].run()  ;
            end

            begin
              gen[15][31].run()  ;
            end
            begin
              drv[15][31].run()  ;
            end
            begin
              mem_check[15][31].run()  ;
            end
            begin
              rf_driver[15][31].run()  ;
            end

            begin
              ldst_driver[16].run()  ;
            end
            begin
              mgr[16].run()  ;
            end
            begin
              oob_drv[16].run()  ;
            end
            begin
              up_check[16].run()  ;
            end
            begin
              gen[16][0].run()  ;
            end
            begin
              drv[16][0].run()  ;
            end
            begin
              mem_check[16][0].run()  ;
            end
            begin
              rf_driver[16][0].run()  ;
            end

            begin
              gen[16][1].run()  ;
            end
            begin
              drv[16][1].run()  ;
            end
            begin
              mem_check[16][1].run()  ;
            end
            begin
              rf_driver[16][1].run()  ;
            end

            begin
              gen[16][2].run()  ;
            end
            begin
              drv[16][2].run()  ;
            end
            begin
              mem_check[16][2].run()  ;
            end
            begin
              rf_driver[16][2].run()  ;
            end

            begin
              gen[16][3].run()  ;
            end
            begin
              drv[16][3].run()  ;
            end
            begin
              mem_check[16][3].run()  ;
            end
            begin
              rf_driver[16][3].run()  ;
            end

            begin
              gen[16][4].run()  ;
            end
            begin
              drv[16][4].run()  ;
            end
            begin
              mem_check[16][4].run()  ;
            end
            begin
              rf_driver[16][4].run()  ;
            end

            begin
              gen[16][5].run()  ;
            end
            begin
              drv[16][5].run()  ;
            end
            begin
              mem_check[16][5].run()  ;
            end
            begin
              rf_driver[16][5].run()  ;
            end

            begin
              gen[16][6].run()  ;
            end
            begin
              drv[16][6].run()  ;
            end
            begin
              mem_check[16][6].run()  ;
            end
            begin
              rf_driver[16][6].run()  ;
            end

            begin
              gen[16][7].run()  ;
            end
            begin
              drv[16][7].run()  ;
            end
            begin
              mem_check[16][7].run()  ;
            end
            begin
              rf_driver[16][7].run()  ;
            end

            begin
              gen[16][8].run()  ;
            end
            begin
              drv[16][8].run()  ;
            end
            begin
              mem_check[16][8].run()  ;
            end
            begin
              rf_driver[16][8].run()  ;
            end

            begin
              gen[16][9].run()  ;
            end
            begin
              drv[16][9].run()  ;
            end
            begin
              mem_check[16][9].run()  ;
            end
            begin
              rf_driver[16][9].run()  ;
            end

            begin
              gen[16][10].run()  ;
            end
            begin
              drv[16][10].run()  ;
            end
            begin
              mem_check[16][10].run()  ;
            end
            begin
              rf_driver[16][10].run()  ;
            end

            begin
              gen[16][11].run()  ;
            end
            begin
              drv[16][11].run()  ;
            end
            begin
              mem_check[16][11].run()  ;
            end
            begin
              rf_driver[16][11].run()  ;
            end

            begin
              gen[16][12].run()  ;
            end
            begin
              drv[16][12].run()  ;
            end
            begin
              mem_check[16][12].run()  ;
            end
            begin
              rf_driver[16][12].run()  ;
            end

            begin
              gen[16][13].run()  ;
            end
            begin
              drv[16][13].run()  ;
            end
            begin
              mem_check[16][13].run()  ;
            end
            begin
              rf_driver[16][13].run()  ;
            end

            begin
              gen[16][14].run()  ;
            end
            begin
              drv[16][14].run()  ;
            end
            begin
              mem_check[16][14].run()  ;
            end
            begin
              rf_driver[16][14].run()  ;
            end

            begin
              gen[16][15].run()  ;
            end
            begin
              drv[16][15].run()  ;
            end
            begin
              mem_check[16][15].run()  ;
            end
            begin
              rf_driver[16][15].run()  ;
            end

            begin
              gen[16][16].run()  ;
            end
            begin
              drv[16][16].run()  ;
            end
            begin
              mem_check[16][16].run()  ;
            end
            begin
              rf_driver[16][16].run()  ;
            end

            begin
              gen[16][17].run()  ;
            end
            begin
              drv[16][17].run()  ;
            end
            begin
              mem_check[16][17].run()  ;
            end
            begin
              rf_driver[16][17].run()  ;
            end

            begin
              gen[16][18].run()  ;
            end
            begin
              drv[16][18].run()  ;
            end
            begin
              mem_check[16][18].run()  ;
            end
            begin
              rf_driver[16][18].run()  ;
            end

            begin
              gen[16][19].run()  ;
            end
            begin
              drv[16][19].run()  ;
            end
            begin
              mem_check[16][19].run()  ;
            end
            begin
              rf_driver[16][19].run()  ;
            end

            begin
              gen[16][20].run()  ;
            end
            begin
              drv[16][20].run()  ;
            end
            begin
              mem_check[16][20].run()  ;
            end
            begin
              rf_driver[16][20].run()  ;
            end

            begin
              gen[16][21].run()  ;
            end
            begin
              drv[16][21].run()  ;
            end
            begin
              mem_check[16][21].run()  ;
            end
            begin
              rf_driver[16][21].run()  ;
            end

            begin
              gen[16][22].run()  ;
            end
            begin
              drv[16][22].run()  ;
            end
            begin
              mem_check[16][22].run()  ;
            end
            begin
              rf_driver[16][22].run()  ;
            end

            begin
              gen[16][23].run()  ;
            end
            begin
              drv[16][23].run()  ;
            end
            begin
              mem_check[16][23].run()  ;
            end
            begin
              rf_driver[16][23].run()  ;
            end

            begin
              gen[16][24].run()  ;
            end
            begin
              drv[16][24].run()  ;
            end
            begin
              mem_check[16][24].run()  ;
            end
            begin
              rf_driver[16][24].run()  ;
            end

            begin
              gen[16][25].run()  ;
            end
            begin
              drv[16][25].run()  ;
            end
            begin
              mem_check[16][25].run()  ;
            end
            begin
              rf_driver[16][25].run()  ;
            end

            begin
              gen[16][26].run()  ;
            end
            begin
              drv[16][26].run()  ;
            end
            begin
              mem_check[16][26].run()  ;
            end
            begin
              rf_driver[16][26].run()  ;
            end

            begin
              gen[16][27].run()  ;
            end
            begin
              drv[16][27].run()  ;
            end
            begin
              mem_check[16][27].run()  ;
            end
            begin
              rf_driver[16][27].run()  ;
            end

            begin
              gen[16][28].run()  ;
            end
            begin
              drv[16][28].run()  ;
            end
            begin
              mem_check[16][28].run()  ;
            end
            begin
              rf_driver[16][28].run()  ;
            end

            begin
              gen[16][29].run()  ;
            end
            begin
              drv[16][29].run()  ;
            end
            begin
              mem_check[16][29].run()  ;
            end
            begin
              rf_driver[16][29].run()  ;
            end

            begin
              gen[16][30].run()  ;
            end
            begin
              drv[16][30].run()  ;
            end
            begin
              mem_check[16][30].run()  ;
            end
            begin
              rf_driver[16][30].run()  ;
            end

            begin
              gen[16][31].run()  ;
            end
            begin
              drv[16][31].run()  ;
            end
            begin
              mem_check[16][31].run()  ;
            end
            begin
              rf_driver[16][31].run()  ;
            end

            begin
              ldst_driver[17].run()  ;
            end
            begin
              mgr[17].run()  ;
            end
            begin
              oob_drv[17].run()  ;
            end
            begin
              up_check[17].run()  ;
            end
            begin
              gen[17][0].run()  ;
            end
            begin
              drv[17][0].run()  ;
            end
            begin
              mem_check[17][0].run()  ;
            end
            begin
              rf_driver[17][0].run()  ;
            end

            begin
              gen[17][1].run()  ;
            end
            begin
              drv[17][1].run()  ;
            end
            begin
              mem_check[17][1].run()  ;
            end
            begin
              rf_driver[17][1].run()  ;
            end

            begin
              gen[17][2].run()  ;
            end
            begin
              drv[17][2].run()  ;
            end
            begin
              mem_check[17][2].run()  ;
            end
            begin
              rf_driver[17][2].run()  ;
            end

            begin
              gen[17][3].run()  ;
            end
            begin
              drv[17][3].run()  ;
            end
            begin
              mem_check[17][3].run()  ;
            end
            begin
              rf_driver[17][3].run()  ;
            end

            begin
              gen[17][4].run()  ;
            end
            begin
              drv[17][4].run()  ;
            end
            begin
              mem_check[17][4].run()  ;
            end
            begin
              rf_driver[17][4].run()  ;
            end

            begin
              gen[17][5].run()  ;
            end
            begin
              drv[17][5].run()  ;
            end
            begin
              mem_check[17][5].run()  ;
            end
            begin
              rf_driver[17][5].run()  ;
            end

            begin
              gen[17][6].run()  ;
            end
            begin
              drv[17][6].run()  ;
            end
            begin
              mem_check[17][6].run()  ;
            end
            begin
              rf_driver[17][6].run()  ;
            end

            begin
              gen[17][7].run()  ;
            end
            begin
              drv[17][7].run()  ;
            end
            begin
              mem_check[17][7].run()  ;
            end
            begin
              rf_driver[17][7].run()  ;
            end

            begin
              gen[17][8].run()  ;
            end
            begin
              drv[17][8].run()  ;
            end
            begin
              mem_check[17][8].run()  ;
            end
            begin
              rf_driver[17][8].run()  ;
            end

            begin
              gen[17][9].run()  ;
            end
            begin
              drv[17][9].run()  ;
            end
            begin
              mem_check[17][9].run()  ;
            end
            begin
              rf_driver[17][9].run()  ;
            end

            begin
              gen[17][10].run()  ;
            end
            begin
              drv[17][10].run()  ;
            end
            begin
              mem_check[17][10].run()  ;
            end
            begin
              rf_driver[17][10].run()  ;
            end

            begin
              gen[17][11].run()  ;
            end
            begin
              drv[17][11].run()  ;
            end
            begin
              mem_check[17][11].run()  ;
            end
            begin
              rf_driver[17][11].run()  ;
            end

            begin
              gen[17][12].run()  ;
            end
            begin
              drv[17][12].run()  ;
            end
            begin
              mem_check[17][12].run()  ;
            end
            begin
              rf_driver[17][12].run()  ;
            end

            begin
              gen[17][13].run()  ;
            end
            begin
              drv[17][13].run()  ;
            end
            begin
              mem_check[17][13].run()  ;
            end
            begin
              rf_driver[17][13].run()  ;
            end

            begin
              gen[17][14].run()  ;
            end
            begin
              drv[17][14].run()  ;
            end
            begin
              mem_check[17][14].run()  ;
            end
            begin
              rf_driver[17][14].run()  ;
            end

            begin
              gen[17][15].run()  ;
            end
            begin
              drv[17][15].run()  ;
            end
            begin
              mem_check[17][15].run()  ;
            end
            begin
              rf_driver[17][15].run()  ;
            end

            begin
              gen[17][16].run()  ;
            end
            begin
              drv[17][16].run()  ;
            end
            begin
              mem_check[17][16].run()  ;
            end
            begin
              rf_driver[17][16].run()  ;
            end

            begin
              gen[17][17].run()  ;
            end
            begin
              drv[17][17].run()  ;
            end
            begin
              mem_check[17][17].run()  ;
            end
            begin
              rf_driver[17][17].run()  ;
            end

            begin
              gen[17][18].run()  ;
            end
            begin
              drv[17][18].run()  ;
            end
            begin
              mem_check[17][18].run()  ;
            end
            begin
              rf_driver[17][18].run()  ;
            end

            begin
              gen[17][19].run()  ;
            end
            begin
              drv[17][19].run()  ;
            end
            begin
              mem_check[17][19].run()  ;
            end
            begin
              rf_driver[17][19].run()  ;
            end

            begin
              gen[17][20].run()  ;
            end
            begin
              drv[17][20].run()  ;
            end
            begin
              mem_check[17][20].run()  ;
            end
            begin
              rf_driver[17][20].run()  ;
            end

            begin
              gen[17][21].run()  ;
            end
            begin
              drv[17][21].run()  ;
            end
            begin
              mem_check[17][21].run()  ;
            end
            begin
              rf_driver[17][21].run()  ;
            end

            begin
              gen[17][22].run()  ;
            end
            begin
              drv[17][22].run()  ;
            end
            begin
              mem_check[17][22].run()  ;
            end
            begin
              rf_driver[17][22].run()  ;
            end

            begin
              gen[17][23].run()  ;
            end
            begin
              drv[17][23].run()  ;
            end
            begin
              mem_check[17][23].run()  ;
            end
            begin
              rf_driver[17][23].run()  ;
            end

            begin
              gen[17][24].run()  ;
            end
            begin
              drv[17][24].run()  ;
            end
            begin
              mem_check[17][24].run()  ;
            end
            begin
              rf_driver[17][24].run()  ;
            end

            begin
              gen[17][25].run()  ;
            end
            begin
              drv[17][25].run()  ;
            end
            begin
              mem_check[17][25].run()  ;
            end
            begin
              rf_driver[17][25].run()  ;
            end

            begin
              gen[17][26].run()  ;
            end
            begin
              drv[17][26].run()  ;
            end
            begin
              mem_check[17][26].run()  ;
            end
            begin
              rf_driver[17][26].run()  ;
            end

            begin
              gen[17][27].run()  ;
            end
            begin
              drv[17][27].run()  ;
            end
            begin
              mem_check[17][27].run()  ;
            end
            begin
              rf_driver[17][27].run()  ;
            end

            begin
              gen[17][28].run()  ;
            end
            begin
              drv[17][28].run()  ;
            end
            begin
              mem_check[17][28].run()  ;
            end
            begin
              rf_driver[17][28].run()  ;
            end

            begin
              gen[17][29].run()  ;
            end
            begin
              drv[17][29].run()  ;
            end
            begin
              mem_check[17][29].run()  ;
            end
            begin
              rf_driver[17][29].run()  ;
            end

            begin
              gen[17][30].run()  ;
            end
            begin
              drv[17][30].run()  ;
            end
            begin
              mem_check[17][30].run()  ;
            end
            begin
              rf_driver[17][30].run()  ;
            end

            begin
              gen[17][31].run()  ;
            end
            begin
              drv[17][31].run()  ;
            end
            begin
              mem_check[17][31].run()  ;
            end
            begin
              rf_driver[17][31].run()  ;
            end

            begin
              ldst_driver[18].run()  ;
            end
            begin
              mgr[18].run()  ;
            end
            begin
              oob_drv[18].run()  ;
            end
            begin
              up_check[18].run()  ;
            end
            begin
              gen[18][0].run()  ;
            end
            begin
              drv[18][0].run()  ;
            end
            begin
              mem_check[18][0].run()  ;
            end
            begin
              rf_driver[18][0].run()  ;
            end

            begin
              gen[18][1].run()  ;
            end
            begin
              drv[18][1].run()  ;
            end
            begin
              mem_check[18][1].run()  ;
            end
            begin
              rf_driver[18][1].run()  ;
            end

            begin
              gen[18][2].run()  ;
            end
            begin
              drv[18][2].run()  ;
            end
            begin
              mem_check[18][2].run()  ;
            end
            begin
              rf_driver[18][2].run()  ;
            end

            begin
              gen[18][3].run()  ;
            end
            begin
              drv[18][3].run()  ;
            end
            begin
              mem_check[18][3].run()  ;
            end
            begin
              rf_driver[18][3].run()  ;
            end

            begin
              gen[18][4].run()  ;
            end
            begin
              drv[18][4].run()  ;
            end
            begin
              mem_check[18][4].run()  ;
            end
            begin
              rf_driver[18][4].run()  ;
            end

            begin
              gen[18][5].run()  ;
            end
            begin
              drv[18][5].run()  ;
            end
            begin
              mem_check[18][5].run()  ;
            end
            begin
              rf_driver[18][5].run()  ;
            end

            begin
              gen[18][6].run()  ;
            end
            begin
              drv[18][6].run()  ;
            end
            begin
              mem_check[18][6].run()  ;
            end
            begin
              rf_driver[18][6].run()  ;
            end

            begin
              gen[18][7].run()  ;
            end
            begin
              drv[18][7].run()  ;
            end
            begin
              mem_check[18][7].run()  ;
            end
            begin
              rf_driver[18][7].run()  ;
            end

            begin
              gen[18][8].run()  ;
            end
            begin
              drv[18][8].run()  ;
            end
            begin
              mem_check[18][8].run()  ;
            end
            begin
              rf_driver[18][8].run()  ;
            end

            begin
              gen[18][9].run()  ;
            end
            begin
              drv[18][9].run()  ;
            end
            begin
              mem_check[18][9].run()  ;
            end
            begin
              rf_driver[18][9].run()  ;
            end

            begin
              gen[18][10].run()  ;
            end
            begin
              drv[18][10].run()  ;
            end
            begin
              mem_check[18][10].run()  ;
            end
            begin
              rf_driver[18][10].run()  ;
            end

            begin
              gen[18][11].run()  ;
            end
            begin
              drv[18][11].run()  ;
            end
            begin
              mem_check[18][11].run()  ;
            end
            begin
              rf_driver[18][11].run()  ;
            end

            begin
              gen[18][12].run()  ;
            end
            begin
              drv[18][12].run()  ;
            end
            begin
              mem_check[18][12].run()  ;
            end
            begin
              rf_driver[18][12].run()  ;
            end

            begin
              gen[18][13].run()  ;
            end
            begin
              drv[18][13].run()  ;
            end
            begin
              mem_check[18][13].run()  ;
            end
            begin
              rf_driver[18][13].run()  ;
            end

            begin
              gen[18][14].run()  ;
            end
            begin
              drv[18][14].run()  ;
            end
            begin
              mem_check[18][14].run()  ;
            end
            begin
              rf_driver[18][14].run()  ;
            end

            begin
              gen[18][15].run()  ;
            end
            begin
              drv[18][15].run()  ;
            end
            begin
              mem_check[18][15].run()  ;
            end
            begin
              rf_driver[18][15].run()  ;
            end

            begin
              gen[18][16].run()  ;
            end
            begin
              drv[18][16].run()  ;
            end
            begin
              mem_check[18][16].run()  ;
            end
            begin
              rf_driver[18][16].run()  ;
            end

            begin
              gen[18][17].run()  ;
            end
            begin
              drv[18][17].run()  ;
            end
            begin
              mem_check[18][17].run()  ;
            end
            begin
              rf_driver[18][17].run()  ;
            end

            begin
              gen[18][18].run()  ;
            end
            begin
              drv[18][18].run()  ;
            end
            begin
              mem_check[18][18].run()  ;
            end
            begin
              rf_driver[18][18].run()  ;
            end

            begin
              gen[18][19].run()  ;
            end
            begin
              drv[18][19].run()  ;
            end
            begin
              mem_check[18][19].run()  ;
            end
            begin
              rf_driver[18][19].run()  ;
            end

            begin
              gen[18][20].run()  ;
            end
            begin
              drv[18][20].run()  ;
            end
            begin
              mem_check[18][20].run()  ;
            end
            begin
              rf_driver[18][20].run()  ;
            end

            begin
              gen[18][21].run()  ;
            end
            begin
              drv[18][21].run()  ;
            end
            begin
              mem_check[18][21].run()  ;
            end
            begin
              rf_driver[18][21].run()  ;
            end

            begin
              gen[18][22].run()  ;
            end
            begin
              drv[18][22].run()  ;
            end
            begin
              mem_check[18][22].run()  ;
            end
            begin
              rf_driver[18][22].run()  ;
            end

            begin
              gen[18][23].run()  ;
            end
            begin
              drv[18][23].run()  ;
            end
            begin
              mem_check[18][23].run()  ;
            end
            begin
              rf_driver[18][23].run()  ;
            end

            begin
              gen[18][24].run()  ;
            end
            begin
              drv[18][24].run()  ;
            end
            begin
              mem_check[18][24].run()  ;
            end
            begin
              rf_driver[18][24].run()  ;
            end

            begin
              gen[18][25].run()  ;
            end
            begin
              drv[18][25].run()  ;
            end
            begin
              mem_check[18][25].run()  ;
            end
            begin
              rf_driver[18][25].run()  ;
            end

            begin
              gen[18][26].run()  ;
            end
            begin
              drv[18][26].run()  ;
            end
            begin
              mem_check[18][26].run()  ;
            end
            begin
              rf_driver[18][26].run()  ;
            end

            begin
              gen[18][27].run()  ;
            end
            begin
              drv[18][27].run()  ;
            end
            begin
              mem_check[18][27].run()  ;
            end
            begin
              rf_driver[18][27].run()  ;
            end

            begin
              gen[18][28].run()  ;
            end
            begin
              drv[18][28].run()  ;
            end
            begin
              mem_check[18][28].run()  ;
            end
            begin
              rf_driver[18][28].run()  ;
            end

            begin
              gen[18][29].run()  ;
            end
            begin
              drv[18][29].run()  ;
            end
            begin
              mem_check[18][29].run()  ;
            end
            begin
              rf_driver[18][29].run()  ;
            end

            begin
              gen[18][30].run()  ;
            end
            begin
              drv[18][30].run()  ;
            end
            begin
              mem_check[18][30].run()  ;
            end
            begin
              rf_driver[18][30].run()  ;
            end

            begin
              gen[18][31].run()  ;
            end
            begin
              drv[18][31].run()  ;
            end
            begin
              mem_check[18][31].run()  ;
            end
            begin
              rf_driver[18][31].run()  ;
            end

            begin
              ldst_driver[19].run()  ;
            end
            begin
              mgr[19].run()  ;
            end
            begin
              oob_drv[19].run()  ;
            end
            begin
              up_check[19].run()  ;
            end
            begin
              gen[19][0].run()  ;
            end
            begin
              drv[19][0].run()  ;
            end
            begin
              mem_check[19][0].run()  ;
            end
            begin
              rf_driver[19][0].run()  ;
            end

            begin
              gen[19][1].run()  ;
            end
            begin
              drv[19][1].run()  ;
            end
            begin
              mem_check[19][1].run()  ;
            end
            begin
              rf_driver[19][1].run()  ;
            end

            begin
              gen[19][2].run()  ;
            end
            begin
              drv[19][2].run()  ;
            end
            begin
              mem_check[19][2].run()  ;
            end
            begin
              rf_driver[19][2].run()  ;
            end

            begin
              gen[19][3].run()  ;
            end
            begin
              drv[19][3].run()  ;
            end
            begin
              mem_check[19][3].run()  ;
            end
            begin
              rf_driver[19][3].run()  ;
            end

            begin
              gen[19][4].run()  ;
            end
            begin
              drv[19][4].run()  ;
            end
            begin
              mem_check[19][4].run()  ;
            end
            begin
              rf_driver[19][4].run()  ;
            end

            begin
              gen[19][5].run()  ;
            end
            begin
              drv[19][5].run()  ;
            end
            begin
              mem_check[19][5].run()  ;
            end
            begin
              rf_driver[19][5].run()  ;
            end

            begin
              gen[19][6].run()  ;
            end
            begin
              drv[19][6].run()  ;
            end
            begin
              mem_check[19][6].run()  ;
            end
            begin
              rf_driver[19][6].run()  ;
            end

            begin
              gen[19][7].run()  ;
            end
            begin
              drv[19][7].run()  ;
            end
            begin
              mem_check[19][7].run()  ;
            end
            begin
              rf_driver[19][7].run()  ;
            end

            begin
              gen[19][8].run()  ;
            end
            begin
              drv[19][8].run()  ;
            end
            begin
              mem_check[19][8].run()  ;
            end
            begin
              rf_driver[19][8].run()  ;
            end

            begin
              gen[19][9].run()  ;
            end
            begin
              drv[19][9].run()  ;
            end
            begin
              mem_check[19][9].run()  ;
            end
            begin
              rf_driver[19][9].run()  ;
            end

            begin
              gen[19][10].run()  ;
            end
            begin
              drv[19][10].run()  ;
            end
            begin
              mem_check[19][10].run()  ;
            end
            begin
              rf_driver[19][10].run()  ;
            end

            begin
              gen[19][11].run()  ;
            end
            begin
              drv[19][11].run()  ;
            end
            begin
              mem_check[19][11].run()  ;
            end
            begin
              rf_driver[19][11].run()  ;
            end

            begin
              gen[19][12].run()  ;
            end
            begin
              drv[19][12].run()  ;
            end
            begin
              mem_check[19][12].run()  ;
            end
            begin
              rf_driver[19][12].run()  ;
            end

            begin
              gen[19][13].run()  ;
            end
            begin
              drv[19][13].run()  ;
            end
            begin
              mem_check[19][13].run()  ;
            end
            begin
              rf_driver[19][13].run()  ;
            end

            begin
              gen[19][14].run()  ;
            end
            begin
              drv[19][14].run()  ;
            end
            begin
              mem_check[19][14].run()  ;
            end
            begin
              rf_driver[19][14].run()  ;
            end

            begin
              gen[19][15].run()  ;
            end
            begin
              drv[19][15].run()  ;
            end
            begin
              mem_check[19][15].run()  ;
            end
            begin
              rf_driver[19][15].run()  ;
            end

            begin
              gen[19][16].run()  ;
            end
            begin
              drv[19][16].run()  ;
            end
            begin
              mem_check[19][16].run()  ;
            end
            begin
              rf_driver[19][16].run()  ;
            end

            begin
              gen[19][17].run()  ;
            end
            begin
              drv[19][17].run()  ;
            end
            begin
              mem_check[19][17].run()  ;
            end
            begin
              rf_driver[19][17].run()  ;
            end

            begin
              gen[19][18].run()  ;
            end
            begin
              drv[19][18].run()  ;
            end
            begin
              mem_check[19][18].run()  ;
            end
            begin
              rf_driver[19][18].run()  ;
            end

            begin
              gen[19][19].run()  ;
            end
            begin
              drv[19][19].run()  ;
            end
            begin
              mem_check[19][19].run()  ;
            end
            begin
              rf_driver[19][19].run()  ;
            end

            begin
              gen[19][20].run()  ;
            end
            begin
              drv[19][20].run()  ;
            end
            begin
              mem_check[19][20].run()  ;
            end
            begin
              rf_driver[19][20].run()  ;
            end

            begin
              gen[19][21].run()  ;
            end
            begin
              drv[19][21].run()  ;
            end
            begin
              mem_check[19][21].run()  ;
            end
            begin
              rf_driver[19][21].run()  ;
            end

            begin
              gen[19][22].run()  ;
            end
            begin
              drv[19][22].run()  ;
            end
            begin
              mem_check[19][22].run()  ;
            end
            begin
              rf_driver[19][22].run()  ;
            end

            begin
              gen[19][23].run()  ;
            end
            begin
              drv[19][23].run()  ;
            end
            begin
              mem_check[19][23].run()  ;
            end
            begin
              rf_driver[19][23].run()  ;
            end

            begin
              gen[19][24].run()  ;
            end
            begin
              drv[19][24].run()  ;
            end
            begin
              mem_check[19][24].run()  ;
            end
            begin
              rf_driver[19][24].run()  ;
            end

            begin
              gen[19][25].run()  ;
            end
            begin
              drv[19][25].run()  ;
            end
            begin
              mem_check[19][25].run()  ;
            end
            begin
              rf_driver[19][25].run()  ;
            end

            begin
              gen[19][26].run()  ;
            end
            begin
              drv[19][26].run()  ;
            end
            begin
              mem_check[19][26].run()  ;
            end
            begin
              rf_driver[19][26].run()  ;
            end

            begin
              gen[19][27].run()  ;
            end
            begin
              drv[19][27].run()  ;
            end
            begin
              mem_check[19][27].run()  ;
            end
            begin
              rf_driver[19][27].run()  ;
            end

            begin
              gen[19][28].run()  ;
            end
            begin
              drv[19][28].run()  ;
            end
            begin
              mem_check[19][28].run()  ;
            end
            begin
              rf_driver[19][28].run()  ;
            end

            begin
              gen[19][29].run()  ;
            end
            begin
              drv[19][29].run()  ;
            end
            begin
              mem_check[19][29].run()  ;
            end
            begin
              rf_driver[19][29].run()  ;
            end

            begin
              gen[19][30].run()  ;
            end
            begin
              drv[19][30].run()  ;
            end
            begin
              mem_check[19][30].run()  ;
            end
            begin
              rf_driver[19][30].run()  ;
            end

            begin
              gen[19][31].run()  ;
            end
            begin
              drv[19][31].run()  ;
            end
            begin
              mem_check[19][31].run()  ;
            end
            begin
              rf_driver[19][31].run()  ;
            end

            begin
              ldst_driver[20].run()  ;
            end
            begin
              mgr[20].run()  ;
            end
            begin
              oob_drv[20].run()  ;
            end
            begin
              up_check[20].run()  ;
            end
            begin
              gen[20][0].run()  ;
            end
            begin
              drv[20][0].run()  ;
            end
            begin
              mem_check[20][0].run()  ;
            end
            begin
              rf_driver[20][0].run()  ;
            end

            begin
              gen[20][1].run()  ;
            end
            begin
              drv[20][1].run()  ;
            end
            begin
              mem_check[20][1].run()  ;
            end
            begin
              rf_driver[20][1].run()  ;
            end

            begin
              gen[20][2].run()  ;
            end
            begin
              drv[20][2].run()  ;
            end
            begin
              mem_check[20][2].run()  ;
            end
            begin
              rf_driver[20][2].run()  ;
            end

            begin
              gen[20][3].run()  ;
            end
            begin
              drv[20][3].run()  ;
            end
            begin
              mem_check[20][3].run()  ;
            end
            begin
              rf_driver[20][3].run()  ;
            end

            begin
              gen[20][4].run()  ;
            end
            begin
              drv[20][4].run()  ;
            end
            begin
              mem_check[20][4].run()  ;
            end
            begin
              rf_driver[20][4].run()  ;
            end

            begin
              gen[20][5].run()  ;
            end
            begin
              drv[20][5].run()  ;
            end
            begin
              mem_check[20][5].run()  ;
            end
            begin
              rf_driver[20][5].run()  ;
            end

            begin
              gen[20][6].run()  ;
            end
            begin
              drv[20][6].run()  ;
            end
            begin
              mem_check[20][6].run()  ;
            end
            begin
              rf_driver[20][6].run()  ;
            end

            begin
              gen[20][7].run()  ;
            end
            begin
              drv[20][7].run()  ;
            end
            begin
              mem_check[20][7].run()  ;
            end
            begin
              rf_driver[20][7].run()  ;
            end

            begin
              gen[20][8].run()  ;
            end
            begin
              drv[20][8].run()  ;
            end
            begin
              mem_check[20][8].run()  ;
            end
            begin
              rf_driver[20][8].run()  ;
            end

            begin
              gen[20][9].run()  ;
            end
            begin
              drv[20][9].run()  ;
            end
            begin
              mem_check[20][9].run()  ;
            end
            begin
              rf_driver[20][9].run()  ;
            end

            begin
              gen[20][10].run()  ;
            end
            begin
              drv[20][10].run()  ;
            end
            begin
              mem_check[20][10].run()  ;
            end
            begin
              rf_driver[20][10].run()  ;
            end

            begin
              gen[20][11].run()  ;
            end
            begin
              drv[20][11].run()  ;
            end
            begin
              mem_check[20][11].run()  ;
            end
            begin
              rf_driver[20][11].run()  ;
            end

            begin
              gen[20][12].run()  ;
            end
            begin
              drv[20][12].run()  ;
            end
            begin
              mem_check[20][12].run()  ;
            end
            begin
              rf_driver[20][12].run()  ;
            end

            begin
              gen[20][13].run()  ;
            end
            begin
              drv[20][13].run()  ;
            end
            begin
              mem_check[20][13].run()  ;
            end
            begin
              rf_driver[20][13].run()  ;
            end

            begin
              gen[20][14].run()  ;
            end
            begin
              drv[20][14].run()  ;
            end
            begin
              mem_check[20][14].run()  ;
            end
            begin
              rf_driver[20][14].run()  ;
            end

            begin
              gen[20][15].run()  ;
            end
            begin
              drv[20][15].run()  ;
            end
            begin
              mem_check[20][15].run()  ;
            end
            begin
              rf_driver[20][15].run()  ;
            end

            begin
              gen[20][16].run()  ;
            end
            begin
              drv[20][16].run()  ;
            end
            begin
              mem_check[20][16].run()  ;
            end
            begin
              rf_driver[20][16].run()  ;
            end

            begin
              gen[20][17].run()  ;
            end
            begin
              drv[20][17].run()  ;
            end
            begin
              mem_check[20][17].run()  ;
            end
            begin
              rf_driver[20][17].run()  ;
            end

            begin
              gen[20][18].run()  ;
            end
            begin
              drv[20][18].run()  ;
            end
            begin
              mem_check[20][18].run()  ;
            end
            begin
              rf_driver[20][18].run()  ;
            end

            begin
              gen[20][19].run()  ;
            end
            begin
              drv[20][19].run()  ;
            end
            begin
              mem_check[20][19].run()  ;
            end
            begin
              rf_driver[20][19].run()  ;
            end

            begin
              gen[20][20].run()  ;
            end
            begin
              drv[20][20].run()  ;
            end
            begin
              mem_check[20][20].run()  ;
            end
            begin
              rf_driver[20][20].run()  ;
            end

            begin
              gen[20][21].run()  ;
            end
            begin
              drv[20][21].run()  ;
            end
            begin
              mem_check[20][21].run()  ;
            end
            begin
              rf_driver[20][21].run()  ;
            end

            begin
              gen[20][22].run()  ;
            end
            begin
              drv[20][22].run()  ;
            end
            begin
              mem_check[20][22].run()  ;
            end
            begin
              rf_driver[20][22].run()  ;
            end

            begin
              gen[20][23].run()  ;
            end
            begin
              drv[20][23].run()  ;
            end
            begin
              mem_check[20][23].run()  ;
            end
            begin
              rf_driver[20][23].run()  ;
            end

            begin
              gen[20][24].run()  ;
            end
            begin
              drv[20][24].run()  ;
            end
            begin
              mem_check[20][24].run()  ;
            end
            begin
              rf_driver[20][24].run()  ;
            end

            begin
              gen[20][25].run()  ;
            end
            begin
              drv[20][25].run()  ;
            end
            begin
              mem_check[20][25].run()  ;
            end
            begin
              rf_driver[20][25].run()  ;
            end

            begin
              gen[20][26].run()  ;
            end
            begin
              drv[20][26].run()  ;
            end
            begin
              mem_check[20][26].run()  ;
            end
            begin
              rf_driver[20][26].run()  ;
            end

            begin
              gen[20][27].run()  ;
            end
            begin
              drv[20][27].run()  ;
            end
            begin
              mem_check[20][27].run()  ;
            end
            begin
              rf_driver[20][27].run()  ;
            end

            begin
              gen[20][28].run()  ;
            end
            begin
              drv[20][28].run()  ;
            end
            begin
              mem_check[20][28].run()  ;
            end
            begin
              rf_driver[20][28].run()  ;
            end

            begin
              gen[20][29].run()  ;
            end
            begin
              drv[20][29].run()  ;
            end
            begin
              mem_check[20][29].run()  ;
            end
            begin
              rf_driver[20][29].run()  ;
            end

            begin
              gen[20][30].run()  ;
            end
            begin
              drv[20][30].run()  ;
            end
            begin
              mem_check[20][30].run()  ;
            end
            begin
              rf_driver[20][30].run()  ;
            end

            begin
              gen[20][31].run()  ;
            end
            begin
              drv[20][31].run()  ;
            end
            begin
              mem_check[20][31].run()  ;
            end
            begin
              rf_driver[20][31].run()  ;
            end

            begin
              ldst_driver[21].run()  ;
            end
            begin
              mgr[21].run()  ;
            end
            begin
              oob_drv[21].run()  ;
            end
            begin
              up_check[21].run()  ;
            end
            begin
              gen[21][0].run()  ;
            end
            begin
              drv[21][0].run()  ;
            end
            begin
              mem_check[21][0].run()  ;
            end
            begin
              rf_driver[21][0].run()  ;
            end

            begin
              gen[21][1].run()  ;
            end
            begin
              drv[21][1].run()  ;
            end
            begin
              mem_check[21][1].run()  ;
            end
            begin
              rf_driver[21][1].run()  ;
            end

            begin
              gen[21][2].run()  ;
            end
            begin
              drv[21][2].run()  ;
            end
            begin
              mem_check[21][2].run()  ;
            end
            begin
              rf_driver[21][2].run()  ;
            end

            begin
              gen[21][3].run()  ;
            end
            begin
              drv[21][3].run()  ;
            end
            begin
              mem_check[21][3].run()  ;
            end
            begin
              rf_driver[21][3].run()  ;
            end

            begin
              gen[21][4].run()  ;
            end
            begin
              drv[21][4].run()  ;
            end
            begin
              mem_check[21][4].run()  ;
            end
            begin
              rf_driver[21][4].run()  ;
            end

            begin
              gen[21][5].run()  ;
            end
            begin
              drv[21][5].run()  ;
            end
            begin
              mem_check[21][5].run()  ;
            end
            begin
              rf_driver[21][5].run()  ;
            end

            begin
              gen[21][6].run()  ;
            end
            begin
              drv[21][6].run()  ;
            end
            begin
              mem_check[21][6].run()  ;
            end
            begin
              rf_driver[21][6].run()  ;
            end

            begin
              gen[21][7].run()  ;
            end
            begin
              drv[21][7].run()  ;
            end
            begin
              mem_check[21][7].run()  ;
            end
            begin
              rf_driver[21][7].run()  ;
            end

            begin
              gen[21][8].run()  ;
            end
            begin
              drv[21][8].run()  ;
            end
            begin
              mem_check[21][8].run()  ;
            end
            begin
              rf_driver[21][8].run()  ;
            end

            begin
              gen[21][9].run()  ;
            end
            begin
              drv[21][9].run()  ;
            end
            begin
              mem_check[21][9].run()  ;
            end
            begin
              rf_driver[21][9].run()  ;
            end

            begin
              gen[21][10].run()  ;
            end
            begin
              drv[21][10].run()  ;
            end
            begin
              mem_check[21][10].run()  ;
            end
            begin
              rf_driver[21][10].run()  ;
            end

            begin
              gen[21][11].run()  ;
            end
            begin
              drv[21][11].run()  ;
            end
            begin
              mem_check[21][11].run()  ;
            end
            begin
              rf_driver[21][11].run()  ;
            end

            begin
              gen[21][12].run()  ;
            end
            begin
              drv[21][12].run()  ;
            end
            begin
              mem_check[21][12].run()  ;
            end
            begin
              rf_driver[21][12].run()  ;
            end

            begin
              gen[21][13].run()  ;
            end
            begin
              drv[21][13].run()  ;
            end
            begin
              mem_check[21][13].run()  ;
            end
            begin
              rf_driver[21][13].run()  ;
            end

            begin
              gen[21][14].run()  ;
            end
            begin
              drv[21][14].run()  ;
            end
            begin
              mem_check[21][14].run()  ;
            end
            begin
              rf_driver[21][14].run()  ;
            end

            begin
              gen[21][15].run()  ;
            end
            begin
              drv[21][15].run()  ;
            end
            begin
              mem_check[21][15].run()  ;
            end
            begin
              rf_driver[21][15].run()  ;
            end

            begin
              gen[21][16].run()  ;
            end
            begin
              drv[21][16].run()  ;
            end
            begin
              mem_check[21][16].run()  ;
            end
            begin
              rf_driver[21][16].run()  ;
            end

            begin
              gen[21][17].run()  ;
            end
            begin
              drv[21][17].run()  ;
            end
            begin
              mem_check[21][17].run()  ;
            end
            begin
              rf_driver[21][17].run()  ;
            end

            begin
              gen[21][18].run()  ;
            end
            begin
              drv[21][18].run()  ;
            end
            begin
              mem_check[21][18].run()  ;
            end
            begin
              rf_driver[21][18].run()  ;
            end

            begin
              gen[21][19].run()  ;
            end
            begin
              drv[21][19].run()  ;
            end
            begin
              mem_check[21][19].run()  ;
            end
            begin
              rf_driver[21][19].run()  ;
            end

            begin
              gen[21][20].run()  ;
            end
            begin
              drv[21][20].run()  ;
            end
            begin
              mem_check[21][20].run()  ;
            end
            begin
              rf_driver[21][20].run()  ;
            end

            begin
              gen[21][21].run()  ;
            end
            begin
              drv[21][21].run()  ;
            end
            begin
              mem_check[21][21].run()  ;
            end
            begin
              rf_driver[21][21].run()  ;
            end

            begin
              gen[21][22].run()  ;
            end
            begin
              drv[21][22].run()  ;
            end
            begin
              mem_check[21][22].run()  ;
            end
            begin
              rf_driver[21][22].run()  ;
            end

            begin
              gen[21][23].run()  ;
            end
            begin
              drv[21][23].run()  ;
            end
            begin
              mem_check[21][23].run()  ;
            end
            begin
              rf_driver[21][23].run()  ;
            end

            begin
              gen[21][24].run()  ;
            end
            begin
              drv[21][24].run()  ;
            end
            begin
              mem_check[21][24].run()  ;
            end
            begin
              rf_driver[21][24].run()  ;
            end

            begin
              gen[21][25].run()  ;
            end
            begin
              drv[21][25].run()  ;
            end
            begin
              mem_check[21][25].run()  ;
            end
            begin
              rf_driver[21][25].run()  ;
            end

            begin
              gen[21][26].run()  ;
            end
            begin
              drv[21][26].run()  ;
            end
            begin
              mem_check[21][26].run()  ;
            end
            begin
              rf_driver[21][26].run()  ;
            end

            begin
              gen[21][27].run()  ;
            end
            begin
              drv[21][27].run()  ;
            end
            begin
              mem_check[21][27].run()  ;
            end
            begin
              rf_driver[21][27].run()  ;
            end

            begin
              gen[21][28].run()  ;
            end
            begin
              drv[21][28].run()  ;
            end
            begin
              mem_check[21][28].run()  ;
            end
            begin
              rf_driver[21][28].run()  ;
            end

            begin
              gen[21][29].run()  ;
            end
            begin
              drv[21][29].run()  ;
            end
            begin
              mem_check[21][29].run()  ;
            end
            begin
              rf_driver[21][29].run()  ;
            end

            begin
              gen[21][30].run()  ;
            end
            begin
              drv[21][30].run()  ;
            end
            begin
              mem_check[21][30].run()  ;
            end
            begin
              rf_driver[21][30].run()  ;
            end

            begin
              gen[21][31].run()  ;
            end
            begin
              drv[21][31].run()  ;
            end
            begin
              mem_check[21][31].run()  ;
            end
            begin
              rf_driver[21][31].run()  ;
            end

            begin
              ldst_driver[22].run()  ;
            end
            begin
              mgr[22].run()  ;
            end
            begin
              oob_drv[22].run()  ;
            end
            begin
              up_check[22].run()  ;
            end
            begin
              gen[22][0].run()  ;
            end
            begin
              drv[22][0].run()  ;
            end
            begin
              mem_check[22][0].run()  ;
            end
            begin
              rf_driver[22][0].run()  ;
            end

            begin
              gen[22][1].run()  ;
            end
            begin
              drv[22][1].run()  ;
            end
            begin
              mem_check[22][1].run()  ;
            end
            begin
              rf_driver[22][1].run()  ;
            end

            begin
              gen[22][2].run()  ;
            end
            begin
              drv[22][2].run()  ;
            end
            begin
              mem_check[22][2].run()  ;
            end
            begin
              rf_driver[22][2].run()  ;
            end

            begin
              gen[22][3].run()  ;
            end
            begin
              drv[22][3].run()  ;
            end
            begin
              mem_check[22][3].run()  ;
            end
            begin
              rf_driver[22][3].run()  ;
            end

            begin
              gen[22][4].run()  ;
            end
            begin
              drv[22][4].run()  ;
            end
            begin
              mem_check[22][4].run()  ;
            end
            begin
              rf_driver[22][4].run()  ;
            end

            begin
              gen[22][5].run()  ;
            end
            begin
              drv[22][5].run()  ;
            end
            begin
              mem_check[22][5].run()  ;
            end
            begin
              rf_driver[22][5].run()  ;
            end

            begin
              gen[22][6].run()  ;
            end
            begin
              drv[22][6].run()  ;
            end
            begin
              mem_check[22][6].run()  ;
            end
            begin
              rf_driver[22][6].run()  ;
            end

            begin
              gen[22][7].run()  ;
            end
            begin
              drv[22][7].run()  ;
            end
            begin
              mem_check[22][7].run()  ;
            end
            begin
              rf_driver[22][7].run()  ;
            end

            begin
              gen[22][8].run()  ;
            end
            begin
              drv[22][8].run()  ;
            end
            begin
              mem_check[22][8].run()  ;
            end
            begin
              rf_driver[22][8].run()  ;
            end

            begin
              gen[22][9].run()  ;
            end
            begin
              drv[22][9].run()  ;
            end
            begin
              mem_check[22][9].run()  ;
            end
            begin
              rf_driver[22][9].run()  ;
            end

            begin
              gen[22][10].run()  ;
            end
            begin
              drv[22][10].run()  ;
            end
            begin
              mem_check[22][10].run()  ;
            end
            begin
              rf_driver[22][10].run()  ;
            end

            begin
              gen[22][11].run()  ;
            end
            begin
              drv[22][11].run()  ;
            end
            begin
              mem_check[22][11].run()  ;
            end
            begin
              rf_driver[22][11].run()  ;
            end

            begin
              gen[22][12].run()  ;
            end
            begin
              drv[22][12].run()  ;
            end
            begin
              mem_check[22][12].run()  ;
            end
            begin
              rf_driver[22][12].run()  ;
            end

            begin
              gen[22][13].run()  ;
            end
            begin
              drv[22][13].run()  ;
            end
            begin
              mem_check[22][13].run()  ;
            end
            begin
              rf_driver[22][13].run()  ;
            end

            begin
              gen[22][14].run()  ;
            end
            begin
              drv[22][14].run()  ;
            end
            begin
              mem_check[22][14].run()  ;
            end
            begin
              rf_driver[22][14].run()  ;
            end

            begin
              gen[22][15].run()  ;
            end
            begin
              drv[22][15].run()  ;
            end
            begin
              mem_check[22][15].run()  ;
            end
            begin
              rf_driver[22][15].run()  ;
            end

            begin
              gen[22][16].run()  ;
            end
            begin
              drv[22][16].run()  ;
            end
            begin
              mem_check[22][16].run()  ;
            end
            begin
              rf_driver[22][16].run()  ;
            end

            begin
              gen[22][17].run()  ;
            end
            begin
              drv[22][17].run()  ;
            end
            begin
              mem_check[22][17].run()  ;
            end
            begin
              rf_driver[22][17].run()  ;
            end

            begin
              gen[22][18].run()  ;
            end
            begin
              drv[22][18].run()  ;
            end
            begin
              mem_check[22][18].run()  ;
            end
            begin
              rf_driver[22][18].run()  ;
            end

            begin
              gen[22][19].run()  ;
            end
            begin
              drv[22][19].run()  ;
            end
            begin
              mem_check[22][19].run()  ;
            end
            begin
              rf_driver[22][19].run()  ;
            end

            begin
              gen[22][20].run()  ;
            end
            begin
              drv[22][20].run()  ;
            end
            begin
              mem_check[22][20].run()  ;
            end
            begin
              rf_driver[22][20].run()  ;
            end

            begin
              gen[22][21].run()  ;
            end
            begin
              drv[22][21].run()  ;
            end
            begin
              mem_check[22][21].run()  ;
            end
            begin
              rf_driver[22][21].run()  ;
            end

            begin
              gen[22][22].run()  ;
            end
            begin
              drv[22][22].run()  ;
            end
            begin
              mem_check[22][22].run()  ;
            end
            begin
              rf_driver[22][22].run()  ;
            end

            begin
              gen[22][23].run()  ;
            end
            begin
              drv[22][23].run()  ;
            end
            begin
              mem_check[22][23].run()  ;
            end
            begin
              rf_driver[22][23].run()  ;
            end

            begin
              gen[22][24].run()  ;
            end
            begin
              drv[22][24].run()  ;
            end
            begin
              mem_check[22][24].run()  ;
            end
            begin
              rf_driver[22][24].run()  ;
            end

            begin
              gen[22][25].run()  ;
            end
            begin
              drv[22][25].run()  ;
            end
            begin
              mem_check[22][25].run()  ;
            end
            begin
              rf_driver[22][25].run()  ;
            end

            begin
              gen[22][26].run()  ;
            end
            begin
              drv[22][26].run()  ;
            end
            begin
              mem_check[22][26].run()  ;
            end
            begin
              rf_driver[22][26].run()  ;
            end

            begin
              gen[22][27].run()  ;
            end
            begin
              drv[22][27].run()  ;
            end
            begin
              mem_check[22][27].run()  ;
            end
            begin
              rf_driver[22][27].run()  ;
            end

            begin
              gen[22][28].run()  ;
            end
            begin
              drv[22][28].run()  ;
            end
            begin
              mem_check[22][28].run()  ;
            end
            begin
              rf_driver[22][28].run()  ;
            end

            begin
              gen[22][29].run()  ;
            end
            begin
              drv[22][29].run()  ;
            end
            begin
              mem_check[22][29].run()  ;
            end
            begin
              rf_driver[22][29].run()  ;
            end

            begin
              gen[22][30].run()  ;
            end
            begin
              drv[22][30].run()  ;
            end
            begin
              mem_check[22][30].run()  ;
            end
            begin
              rf_driver[22][30].run()  ;
            end

            begin
              gen[22][31].run()  ;
            end
            begin
              drv[22][31].run()  ;
            end
            begin
              mem_check[22][31].run()  ;
            end
            begin
              rf_driver[22][31].run()  ;
            end

            begin
              ldst_driver[23].run()  ;
            end
            begin
              mgr[23].run()  ;
            end
            begin
              oob_drv[23].run()  ;
            end
            begin
              up_check[23].run()  ;
            end
            begin
              gen[23][0].run()  ;
            end
            begin
              drv[23][0].run()  ;
            end
            begin
              mem_check[23][0].run()  ;
            end
            begin
              rf_driver[23][0].run()  ;
            end

            begin
              gen[23][1].run()  ;
            end
            begin
              drv[23][1].run()  ;
            end
            begin
              mem_check[23][1].run()  ;
            end
            begin
              rf_driver[23][1].run()  ;
            end

            begin
              gen[23][2].run()  ;
            end
            begin
              drv[23][2].run()  ;
            end
            begin
              mem_check[23][2].run()  ;
            end
            begin
              rf_driver[23][2].run()  ;
            end

            begin
              gen[23][3].run()  ;
            end
            begin
              drv[23][3].run()  ;
            end
            begin
              mem_check[23][3].run()  ;
            end
            begin
              rf_driver[23][3].run()  ;
            end

            begin
              gen[23][4].run()  ;
            end
            begin
              drv[23][4].run()  ;
            end
            begin
              mem_check[23][4].run()  ;
            end
            begin
              rf_driver[23][4].run()  ;
            end

            begin
              gen[23][5].run()  ;
            end
            begin
              drv[23][5].run()  ;
            end
            begin
              mem_check[23][5].run()  ;
            end
            begin
              rf_driver[23][5].run()  ;
            end

            begin
              gen[23][6].run()  ;
            end
            begin
              drv[23][6].run()  ;
            end
            begin
              mem_check[23][6].run()  ;
            end
            begin
              rf_driver[23][6].run()  ;
            end

            begin
              gen[23][7].run()  ;
            end
            begin
              drv[23][7].run()  ;
            end
            begin
              mem_check[23][7].run()  ;
            end
            begin
              rf_driver[23][7].run()  ;
            end

            begin
              gen[23][8].run()  ;
            end
            begin
              drv[23][8].run()  ;
            end
            begin
              mem_check[23][8].run()  ;
            end
            begin
              rf_driver[23][8].run()  ;
            end

            begin
              gen[23][9].run()  ;
            end
            begin
              drv[23][9].run()  ;
            end
            begin
              mem_check[23][9].run()  ;
            end
            begin
              rf_driver[23][9].run()  ;
            end

            begin
              gen[23][10].run()  ;
            end
            begin
              drv[23][10].run()  ;
            end
            begin
              mem_check[23][10].run()  ;
            end
            begin
              rf_driver[23][10].run()  ;
            end

            begin
              gen[23][11].run()  ;
            end
            begin
              drv[23][11].run()  ;
            end
            begin
              mem_check[23][11].run()  ;
            end
            begin
              rf_driver[23][11].run()  ;
            end

            begin
              gen[23][12].run()  ;
            end
            begin
              drv[23][12].run()  ;
            end
            begin
              mem_check[23][12].run()  ;
            end
            begin
              rf_driver[23][12].run()  ;
            end

            begin
              gen[23][13].run()  ;
            end
            begin
              drv[23][13].run()  ;
            end
            begin
              mem_check[23][13].run()  ;
            end
            begin
              rf_driver[23][13].run()  ;
            end

            begin
              gen[23][14].run()  ;
            end
            begin
              drv[23][14].run()  ;
            end
            begin
              mem_check[23][14].run()  ;
            end
            begin
              rf_driver[23][14].run()  ;
            end

            begin
              gen[23][15].run()  ;
            end
            begin
              drv[23][15].run()  ;
            end
            begin
              mem_check[23][15].run()  ;
            end
            begin
              rf_driver[23][15].run()  ;
            end

            begin
              gen[23][16].run()  ;
            end
            begin
              drv[23][16].run()  ;
            end
            begin
              mem_check[23][16].run()  ;
            end
            begin
              rf_driver[23][16].run()  ;
            end

            begin
              gen[23][17].run()  ;
            end
            begin
              drv[23][17].run()  ;
            end
            begin
              mem_check[23][17].run()  ;
            end
            begin
              rf_driver[23][17].run()  ;
            end

            begin
              gen[23][18].run()  ;
            end
            begin
              drv[23][18].run()  ;
            end
            begin
              mem_check[23][18].run()  ;
            end
            begin
              rf_driver[23][18].run()  ;
            end

            begin
              gen[23][19].run()  ;
            end
            begin
              drv[23][19].run()  ;
            end
            begin
              mem_check[23][19].run()  ;
            end
            begin
              rf_driver[23][19].run()  ;
            end

            begin
              gen[23][20].run()  ;
            end
            begin
              drv[23][20].run()  ;
            end
            begin
              mem_check[23][20].run()  ;
            end
            begin
              rf_driver[23][20].run()  ;
            end

            begin
              gen[23][21].run()  ;
            end
            begin
              drv[23][21].run()  ;
            end
            begin
              mem_check[23][21].run()  ;
            end
            begin
              rf_driver[23][21].run()  ;
            end

            begin
              gen[23][22].run()  ;
            end
            begin
              drv[23][22].run()  ;
            end
            begin
              mem_check[23][22].run()  ;
            end
            begin
              rf_driver[23][22].run()  ;
            end

            begin
              gen[23][23].run()  ;
            end
            begin
              drv[23][23].run()  ;
            end
            begin
              mem_check[23][23].run()  ;
            end
            begin
              rf_driver[23][23].run()  ;
            end

            begin
              gen[23][24].run()  ;
            end
            begin
              drv[23][24].run()  ;
            end
            begin
              mem_check[23][24].run()  ;
            end
            begin
              rf_driver[23][24].run()  ;
            end

            begin
              gen[23][25].run()  ;
            end
            begin
              drv[23][25].run()  ;
            end
            begin
              mem_check[23][25].run()  ;
            end
            begin
              rf_driver[23][25].run()  ;
            end

            begin
              gen[23][26].run()  ;
            end
            begin
              drv[23][26].run()  ;
            end
            begin
              mem_check[23][26].run()  ;
            end
            begin
              rf_driver[23][26].run()  ;
            end

            begin
              gen[23][27].run()  ;
            end
            begin
              drv[23][27].run()  ;
            end
            begin
              mem_check[23][27].run()  ;
            end
            begin
              rf_driver[23][27].run()  ;
            end

            begin
              gen[23][28].run()  ;
            end
            begin
              drv[23][28].run()  ;
            end
            begin
              mem_check[23][28].run()  ;
            end
            begin
              rf_driver[23][28].run()  ;
            end

            begin
              gen[23][29].run()  ;
            end
            begin
              drv[23][29].run()  ;
            end
            begin
              mem_check[23][29].run()  ;
            end
            begin
              rf_driver[23][29].run()  ;
            end

            begin
              gen[23][30].run()  ;
            end
            begin
              drv[23][30].run()  ;
            end
            begin
              mem_check[23][30].run()  ;
            end
            begin
              rf_driver[23][30].run()  ;
            end

            begin
              gen[23][31].run()  ;
            end
            begin
              drv[23][31].run()  ;
            end
            begin
              mem_check[23][31].run()  ;
            end
            begin
              rf_driver[23][31].run()  ;
            end

            begin
              ldst_driver[24].run()  ;
            end
            begin
              mgr[24].run()  ;
            end
            begin
              oob_drv[24].run()  ;
            end
            begin
              up_check[24].run()  ;
            end
            begin
              gen[24][0].run()  ;
            end
            begin
              drv[24][0].run()  ;
            end
            begin
              mem_check[24][0].run()  ;
            end
            begin
              rf_driver[24][0].run()  ;
            end

            begin
              gen[24][1].run()  ;
            end
            begin
              drv[24][1].run()  ;
            end
            begin
              mem_check[24][1].run()  ;
            end
            begin
              rf_driver[24][1].run()  ;
            end

            begin
              gen[24][2].run()  ;
            end
            begin
              drv[24][2].run()  ;
            end
            begin
              mem_check[24][2].run()  ;
            end
            begin
              rf_driver[24][2].run()  ;
            end

            begin
              gen[24][3].run()  ;
            end
            begin
              drv[24][3].run()  ;
            end
            begin
              mem_check[24][3].run()  ;
            end
            begin
              rf_driver[24][3].run()  ;
            end

            begin
              gen[24][4].run()  ;
            end
            begin
              drv[24][4].run()  ;
            end
            begin
              mem_check[24][4].run()  ;
            end
            begin
              rf_driver[24][4].run()  ;
            end

            begin
              gen[24][5].run()  ;
            end
            begin
              drv[24][5].run()  ;
            end
            begin
              mem_check[24][5].run()  ;
            end
            begin
              rf_driver[24][5].run()  ;
            end

            begin
              gen[24][6].run()  ;
            end
            begin
              drv[24][6].run()  ;
            end
            begin
              mem_check[24][6].run()  ;
            end
            begin
              rf_driver[24][6].run()  ;
            end

            begin
              gen[24][7].run()  ;
            end
            begin
              drv[24][7].run()  ;
            end
            begin
              mem_check[24][7].run()  ;
            end
            begin
              rf_driver[24][7].run()  ;
            end

            begin
              gen[24][8].run()  ;
            end
            begin
              drv[24][8].run()  ;
            end
            begin
              mem_check[24][8].run()  ;
            end
            begin
              rf_driver[24][8].run()  ;
            end

            begin
              gen[24][9].run()  ;
            end
            begin
              drv[24][9].run()  ;
            end
            begin
              mem_check[24][9].run()  ;
            end
            begin
              rf_driver[24][9].run()  ;
            end

            begin
              gen[24][10].run()  ;
            end
            begin
              drv[24][10].run()  ;
            end
            begin
              mem_check[24][10].run()  ;
            end
            begin
              rf_driver[24][10].run()  ;
            end

            begin
              gen[24][11].run()  ;
            end
            begin
              drv[24][11].run()  ;
            end
            begin
              mem_check[24][11].run()  ;
            end
            begin
              rf_driver[24][11].run()  ;
            end

            begin
              gen[24][12].run()  ;
            end
            begin
              drv[24][12].run()  ;
            end
            begin
              mem_check[24][12].run()  ;
            end
            begin
              rf_driver[24][12].run()  ;
            end

            begin
              gen[24][13].run()  ;
            end
            begin
              drv[24][13].run()  ;
            end
            begin
              mem_check[24][13].run()  ;
            end
            begin
              rf_driver[24][13].run()  ;
            end

            begin
              gen[24][14].run()  ;
            end
            begin
              drv[24][14].run()  ;
            end
            begin
              mem_check[24][14].run()  ;
            end
            begin
              rf_driver[24][14].run()  ;
            end

            begin
              gen[24][15].run()  ;
            end
            begin
              drv[24][15].run()  ;
            end
            begin
              mem_check[24][15].run()  ;
            end
            begin
              rf_driver[24][15].run()  ;
            end

            begin
              gen[24][16].run()  ;
            end
            begin
              drv[24][16].run()  ;
            end
            begin
              mem_check[24][16].run()  ;
            end
            begin
              rf_driver[24][16].run()  ;
            end

            begin
              gen[24][17].run()  ;
            end
            begin
              drv[24][17].run()  ;
            end
            begin
              mem_check[24][17].run()  ;
            end
            begin
              rf_driver[24][17].run()  ;
            end

            begin
              gen[24][18].run()  ;
            end
            begin
              drv[24][18].run()  ;
            end
            begin
              mem_check[24][18].run()  ;
            end
            begin
              rf_driver[24][18].run()  ;
            end

            begin
              gen[24][19].run()  ;
            end
            begin
              drv[24][19].run()  ;
            end
            begin
              mem_check[24][19].run()  ;
            end
            begin
              rf_driver[24][19].run()  ;
            end

            begin
              gen[24][20].run()  ;
            end
            begin
              drv[24][20].run()  ;
            end
            begin
              mem_check[24][20].run()  ;
            end
            begin
              rf_driver[24][20].run()  ;
            end

            begin
              gen[24][21].run()  ;
            end
            begin
              drv[24][21].run()  ;
            end
            begin
              mem_check[24][21].run()  ;
            end
            begin
              rf_driver[24][21].run()  ;
            end

            begin
              gen[24][22].run()  ;
            end
            begin
              drv[24][22].run()  ;
            end
            begin
              mem_check[24][22].run()  ;
            end
            begin
              rf_driver[24][22].run()  ;
            end

            begin
              gen[24][23].run()  ;
            end
            begin
              drv[24][23].run()  ;
            end
            begin
              mem_check[24][23].run()  ;
            end
            begin
              rf_driver[24][23].run()  ;
            end

            begin
              gen[24][24].run()  ;
            end
            begin
              drv[24][24].run()  ;
            end
            begin
              mem_check[24][24].run()  ;
            end
            begin
              rf_driver[24][24].run()  ;
            end

            begin
              gen[24][25].run()  ;
            end
            begin
              drv[24][25].run()  ;
            end
            begin
              mem_check[24][25].run()  ;
            end
            begin
              rf_driver[24][25].run()  ;
            end

            begin
              gen[24][26].run()  ;
            end
            begin
              drv[24][26].run()  ;
            end
            begin
              mem_check[24][26].run()  ;
            end
            begin
              rf_driver[24][26].run()  ;
            end

            begin
              gen[24][27].run()  ;
            end
            begin
              drv[24][27].run()  ;
            end
            begin
              mem_check[24][27].run()  ;
            end
            begin
              rf_driver[24][27].run()  ;
            end

            begin
              gen[24][28].run()  ;
            end
            begin
              drv[24][28].run()  ;
            end
            begin
              mem_check[24][28].run()  ;
            end
            begin
              rf_driver[24][28].run()  ;
            end

            begin
              gen[24][29].run()  ;
            end
            begin
              drv[24][29].run()  ;
            end
            begin
              mem_check[24][29].run()  ;
            end
            begin
              rf_driver[24][29].run()  ;
            end

            begin
              gen[24][30].run()  ;
            end
            begin
              drv[24][30].run()  ;
            end
            begin
              mem_check[24][30].run()  ;
            end
            begin
              rf_driver[24][30].run()  ;
            end

            begin
              gen[24][31].run()  ;
            end
            begin
              drv[24][31].run()  ;
            end
            begin
              mem_check[24][31].run()  ;
            end
            begin
              rf_driver[24][31].run()  ;
            end

            begin
              ldst_driver[25].run()  ;
            end
            begin
              mgr[25].run()  ;
            end
            begin
              oob_drv[25].run()  ;
            end
            begin
              up_check[25].run()  ;
            end
            begin
              gen[25][0].run()  ;
            end
            begin
              drv[25][0].run()  ;
            end
            begin
              mem_check[25][0].run()  ;
            end
            begin
              rf_driver[25][0].run()  ;
            end

            begin
              gen[25][1].run()  ;
            end
            begin
              drv[25][1].run()  ;
            end
            begin
              mem_check[25][1].run()  ;
            end
            begin
              rf_driver[25][1].run()  ;
            end

            begin
              gen[25][2].run()  ;
            end
            begin
              drv[25][2].run()  ;
            end
            begin
              mem_check[25][2].run()  ;
            end
            begin
              rf_driver[25][2].run()  ;
            end

            begin
              gen[25][3].run()  ;
            end
            begin
              drv[25][3].run()  ;
            end
            begin
              mem_check[25][3].run()  ;
            end
            begin
              rf_driver[25][3].run()  ;
            end

            begin
              gen[25][4].run()  ;
            end
            begin
              drv[25][4].run()  ;
            end
            begin
              mem_check[25][4].run()  ;
            end
            begin
              rf_driver[25][4].run()  ;
            end

            begin
              gen[25][5].run()  ;
            end
            begin
              drv[25][5].run()  ;
            end
            begin
              mem_check[25][5].run()  ;
            end
            begin
              rf_driver[25][5].run()  ;
            end

            begin
              gen[25][6].run()  ;
            end
            begin
              drv[25][6].run()  ;
            end
            begin
              mem_check[25][6].run()  ;
            end
            begin
              rf_driver[25][6].run()  ;
            end

            begin
              gen[25][7].run()  ;
            end
            begin
              drv[25][7].run()  ;
            end
            begin
              mem_check[25][7].run()  ;
            end
            begin
              rf_driver[25][7].run()  ;
            end

            begin
              gen[25][8].run()  ;
            end
            begin
              drv[25][8].run()  ;
            end
            begin
              mem_check[25][8].run()  ;
            end
            begin
              rf_driver[25][8].run()  ;
            end

            begin
              gen[25][9].run()  ;
            end
            begin
              drv[25][9].run()  ;
            end
            begin
              mem_check[25][9].run()  ;
            end
            begin
              rf_driver[25][9].run()  ;
            end

            begin
              gen[25][10].run()  ;
            end
            begin
              drv[25][10].run()  ;
            end
            begin
              mem_check[25][10].run()  ;
            end
            begin
              rf_driver[25][10].run()  ;
            end

            begin
              gen[25][11].run()  ;
            end
            begin
              drv[25][11].run()  ;
            end
            begin
              mem_check[25][11].run()  ;
            end
            begin
              rf_driver[25][11].run()  ;
            end

            begin
              gen[25][12].run()  ;
            end
            begin
              drv[25][12].run()  ;
            end
            begin
              mem_check[25][12].run()  ;
            end
            begin
              rf_driver[25][12].run()  ;
            end

            begin
              gen[25][13].run()  ;
            end
            begin
              drv[25][13].run()  ;
            end
            begin
              mem_check[25][13].run()  ;
            end
            begin
              rf_driver[25][13].run()  ;
            end

            begin
              gen[25][14].run()  ;
            end
            begin
              drv[25][14].run()  ;
            end
            begin
              mem_check[25][14].run()  ;
            end
            begin
              rf_driver[25][14].run()  ;
            end

            begin
              gen[25][15].run()  ;
            end
            begin
              drv[25][15].run()  ;
            end
            begin
              mem_check[25][15].run()  ;
            end
            begin
              rf_driver[25][15].run()  ;
            end

            begin
              gen[25][16].run()  ;
            end
            begin
              drv[25][16].run()  ;
            end
            begin
              mem_check[25][16].run()  ;
            end
            begin
              rf_driver[25][16].run()  ;
            end

            begin
              gen[25][17].run()  ;
            end
            begin
              drv[25][17].run()  ;
            end
            begin
              mem_check[25][17].run()  ;
            end
            begin
              rf_driver[25][17].run()  ;
            end

            begin
              gen[25][18].run()  ;
            end
            begin
              drv[25][18].run()  ;
            end
            begin
              mem_check[25][18].run()  ;
            end
            begin
              rf_driver[25][18].run()  ;
            end

            begin
              gen[25][19].run()  ;
            end
            begin
              drv[25][19].run()  ;
            end
            begin
              mem_check[25][19].run()  ;
            end
            begin
              rf_driver[25][19].run()  ;
            end

            begin
              gen[25][20].run()  ;
            end
            begin
              drv[25][20].run()  ;
            end
            begin
              mem_check[25][20].run()  ;
            end
            begin
              rf_driver[25][20].run()  ;
            end

            begin
              gen[25][21].run()  ;
            end
            begin
              drv[25][21].run()  ;
            end
            begin
              mem_check[25][21].run()  ;
            end
            begin
              rf_driver[25][21].run()  ;
            end

            begin
              gen[25][22].run()  ;
            end
            begin
              drv[25][22].run()  ;
            end
            begin
              mem_check[25][22].run()  ;
            end
            begin
              rf_driver[25][22].run()  ;
            end

            begin
              gen[25][23].run()  ;
            end
            begin
              drv[25][23].run()  ;
            end
            begin
              mem_check[25][23].run()  ;
            end
            begin
              rf_driver[25][23].run()  ;
            end

            begin
              gen[25][24].run()  ;
            end
            begin
              drv[25][24].run()  ;
            end
            begin
              mem_check[25][24].run()  ;
            end
            begin
              rf_driver[25][24].run()  ;
            end

            begin
              gen[25][25].run()  ;
            end
            begin
              drv[25][25].run()  ;
            end
            begin
              mem_check[25][25].run()  ;
            end
            begin
              rf_driver[25][25].run()  ;
            end

            begin
              gen[25][26].run()  ;
            end
            begin
              drv[25][26].run()  ;
            end
            begin
              mem_check[25][26].run()  ;
            end
            begin
              rf_driver[25][26].run()  ;
            end

            begin
              gen[25][27].run()  ;
            end
            begin
              drv[25][27].run()  ;
            end
            begin
              mem_check[25][27].run()  ;
            end
            begin
              rf_driver[25][27].run()  ;
            end

            begin
              gen[25][28].run()  ;
            end
            begin
              drv[25][28].run()  ;
            end
            begin
              mem_check[25][28].run()  ;
            end
            begin
              rf_driver[25][28].run()  ;
            end

            begin
              gen[25][29].run()  ;
            end
            begin
              drv[25][29].run()  ;
            end
            begin
              mem_check[25][29].run()  ;
            end
            begin
              rf_driver[25][29].run()  ;
            end

            begin
              gen[25][30].run()  ;
            end
            begin
              drv[25][30].run()  ;
            end
            begin
              mem_check[25][30].run()  ;
            end
            begin
              rf_driver[25][30].run()  ;
            end

            begin
              gen[25][31].run()  ;
            end
            begin
              drv[25][31].run()  ;
            end
            begin
              mem_check[25][31].run()  ;
            end
            begin
              rf_driver[25][31].run()  ;
            end

            begin
              ldst_driver[26].run()  ;
            end
            begin
              mgr[26].run()  ;
            end
            begin
              oob_drv[26].run()  ;
            end
            begin
              up_check[26].run()  ;
            end
            begin
              gen[26][0].run()  ;
            end
            begin
              drv[26][0].run()  ;
            end
            begin
              mem_check[26][0].run()  ;
            end
            begin
              rf_driver[26][0].run()  ;
            end

            begin
              gen[26][1].run()  ;
            end
            begin
              drv[26][1].run()  ;
            end
            begin
              mem_check[26][1].run()  ;
            end
            begin
              rf_driver[26][1].run()  ;
            end

            begin
              gen[26][2].run()  ;
            end
            begin
              drv[26][2].run()  ;
            end
            begin
              mem_check[26][2].run()  ;
            end
            begin
              rf_driver[26][2].run()  ;
            end

            begin
              gen[26][3].run()  ;
            end
            begin
              drv[26][3].run()  ;
            end
            begin
              mem_check[26][3].run()  ;
            end
            begin
              rf_driver[26][3].run()  ;
            end

            begin
              gen[26][4].run()  ;
            end
            begin
              drv[26][4].run()  ;
            end
            begin
              mem_check[26][4].run()  ;
            end
            begin
              rf_driver[26][4].run()  ;
            end

            begin
              gen[26][5].run()  ;
            end
            begin
              drv[26][5].run()  ;
            end
            begin
              mem_check[26][5].run()  ;
            end
            begin
              rf_driver[26][5].run()  ;
            end

            begin
              gen[26][6].run()  ;
            end
            begin
              drv[26][6].run()  ;
            end
            begin
              mem_check[26][6].run()  ;
            end
            begin
              rf_driver[26][6].run()  ;
            end

            begin
              gen[26][7].run()  ;
            end
            begin
              drv[26][7].run()  ;
            end
            begin
              mem_check[26][7].run()  ;
            end
            begin
              rf_driver[26][7].run()  ;
            end

            begin
              gen[26][8].run()  ;
            end
            begin
              drv[26][8].run()  ;
            end
            begin
              mem_check[26][8].run()  ;
            end
            begin
              rf_driver[26][8].run()  ;
            end

            begin
              gen[26][9].run()  ;
            end
            begin
              drv[26][9].run()  ;
            end
            begin
              mem_check[26][9].run()  ;
            end
            begin
              rf_driver[26][9].run()  ;
            end

            begin
              gen[26][10].run()  ;
            end
            begin
              drv[26][10].run()  ;
            end
            begin
              mem_check[26][10].run()  ;
            end
            begin
              rf_driver[26][10].run()  ;
            end

            begin
              gen[26][11].run()  ;
            end
            begin
              drv[26][11].run()  ;
            end
            begin
              mem_check[26][11].run()  ;
            end
            begin
              rf_driver[26][11].run()  ;
            end

            begin
              gen[26][12].run()  ;
            end
            begin
              drv[26][12].run()  ;
            end
            begin
              mem_check[26][12].run()  ;
            end
            begin
              rf_driver[26][12].run()  ;
            end

            begin
              gen[26][13].run()  ;
            end
            begin
              drv[26][13].run()  ;
            end
            begin
              mem_check[26][13].run()  ;
            end
            begin
              rf_driver[26][13].run()  ;
            end

            begin
              gen[26][14].run()  ;
            end
            begin
              drv[26][14].run()  ;
            end
            begin
              mem_check[26][14].run()  ;
            end
            begin
              rf_driver[26][14].run()  ;
            end

            begin
              gen[26][15].run()  ;
            end
            begin
              drv[26][15].run()  ;
            end
            begin
              mem_check[26][15].run()  ;
            end
            begin
              rf_driver[26][15].run()  ;
            end

            begin
              gen[26][16].run()  ;
            end
            begin
              drv[26][16].run()  ;
            end
            begin
              mem_check[26][16].run()  ;
            end
            begin
              rf_driver[26][16].run()  ;
            end

            begin
              gen[26][17].run()  ;
            end
            begin
              drv[26][17].run()  ;
            end
            begin
              mem_check[26][17].run()  ;
            end
            begin
              rf_driver[26][17].run()  ;
            end

            begin
              gen[26][18].run()  ;
            end
            begin
              drv[26][18].run()  ;
            end
            begin
              mem_check[26][18].run()  ;
            end
            begin
              rf_driver[26][18].run()  ;
            end

            begin
              gen[26][19].run()  ;
            end
            begin
              drv[26][19].run()  ;
            end
            begin
              mem_check[26][19].run()  ;
            end
            begin
              rf_driver[26][19].run()  ;
            end

            begin
              gen[26][20].run()  ;
            end
            begin
              drv[26][20].run()  ;
            end
            begin
              mem_check[26][20].run()  ;
            end
            begin
              rf_driver[26][20].run()  ;
            end

            begin
              gen[26][21].run()  ;
            end
            begin
              drv[26][21].run()  ;
            end
            begin
              mem_check[26][21].run()  ;
            end
            begin
              rf_driver[26][21].run()  ;
            end

            begin
              gen[26][22].run()  ;
            end
            begin
              drv[26][22].run()  ;
            end
            begin
              mem_check[26][22].run()  ;
            end
            begin
              rf_driver[26][22].run()  ;
            end

            begin
              gen[26][23].run()  ;
            end
            begin
              drv[26][23].run()  ;
            end
            begin
              mem_check[26][23].run()  ;
            end
            begin
              rf_driver[26][23].run()  ;
            end

            begin
              gen[26][24].run()  ;
            end
            begin
              drv[26][24].run()  ;
            end
            begin
              mem_check[26][24].run()  ;
            end
            begin
              rf_driver[26][24].run()  ;
            end

            begin
              gen[26][25].run()  ;
            end
            begin
              drv[26][25].run()  ;
            end
            begin
              mem_check[26][25].run()  ;
            end
            begin
              rf_driver[26][25].run()  ;
            end

            begin
              gen[26][26].run()  ;
            end
            begin
              drv[26][26].run()  ;
            end
            begin
              mem_check[26][26].run()  ;
            end
            begin
              rf_driver[26][26].run()  ;
            end

            begin
              gen[26][27].run()  ;
            end
            begin
              drv[26][27].run()  ;
            end
            begin
              mem_check[26][27].run()  ;
            end
            begin
              rf_driver[26][27].run()  ;
            end

            begin
              gen[26][28].run()  ;
            end
            begin
              drv[26][28].run()  ;
            end
            begin
              mem_check[26][28].run()  ;
            end
            begin
              rf_driver[26][28].run()  ;
            end

            begin
              gen[26][29].run()  ;
            end
            begin
              drv[26][29].run()  ;
            end
            begin
              mem_check[26][29].run()  ;
            end
            begin
              rf_driver[26][29].run()  ;
            end

            begin
              gen[26][30].run()  ;
            end
            begin
              drv[26][30].run()  ;
            end
            begin
              mem_check[26][30].run()  ;
            end
            begin
              rf_driver[26][30].run()  ;
            end

            begin
              gen[26][31].run()  ;
            end
            begin
              drv[26][31].run()  ;
            end
            begin
              mem_check[26][31].run()  ;
            end
            begin
              rf_driver[26][31].run()  ;
            end

            begin
              ldst_driver[27].run()  ;
            end
            begin
              mgr[27].run()  ;
            end
            begin
              oob_drv[27].run()  ;
            end
            begin
              up_check[27].run()  ;
            end
            begin
              gen[27][0].run()  ;
            end
            begin
              drv[27][0].run()  ;
            end
            begin
              mem_check[27][0].run()  ;
            end
            begin
              rf_driver[27][0].run()  ;
            end

            begin
              gen[27][1].run()  ;
            end
            begin
              drv[27][1].run()  ;
            end
            begin
              mem_check[27][1].run()  ;
            end
            begin
              rf_driver[27][1].run()  ;
            end

            begin
              gen[27][2].run()  ;
            end
            begin
              drv[27][2].run()  ;
            end
            begin
              mem_check[27][2].run()  ;
            end
            begin
              rf_driver[27][2].run()  ;
            end

            begin
              gen[27][3].run()  ;
            end
            begin
              drv[27][3].run()  ;
            end
            begin
              mem_check[27][3].run()  ;
            end
            begin
              rf_driver[27][3].run()  ;
            end

            begin
              gen[27][4].run()  ;
            end
            begin
              drv[27][4].run()  ;
            end
            begin
              mem_check[27][4].run()  ;
            end
            begin
              rf_driver[27][4].run()  ;
            end

            begin
              gen[27][5].run()  ;
            end
            begin
              drv[27][5].run()  ;
            end
            begin
              mem_check[27][5].run()  ;
            end
            begin
              rf_driver[27][5].run()  ;
            end

            begin
              gen[27][6].run()  ;
            end
            begin
              drv[27][6].run()  ;
            end
            begin
              mem_check[27][6].run()  ;
            end
            begin
              rf_driver[27][6].run()  ;
            end

            begin
              gen[27][7].run()  ;
            end
            begin
              drv[27][7].run()  ;
            end
            begin
              mem_check[27][7].run()  ;
            end
            begin
              rf_driver[27][7].run()  ;
            end

            begin
              gen[27][8].run()  ;
            end
            begin
              drv[27][8].run()  ;
            end
            begin
              mem_check[27][8].run()  ;
            end
            begin
              rf_driver[27][8].run()  ;
            end

            begin
              gen[27][9].run()  ;
            end
            begin
              drv[27][9].run()  ;
            end
            begin
              mem_check[27][9].run()  ;
            end
            begin
              rf_driver[27][9].run()  ;
            end

            begin
              gen[27][10].run()  ;
            end
            begin
              drv[27][10].run()  ;
            end
            begin
              mem_check[27][10].run()  ;
            end
            begin
              rf_driver[27][10].run()  ;
            end

            begin
              gen[27][11].run()  ;
            end
            begin
              drv[27][11].run()  ;
            end
            begin
              mem_check[27][11].run()  ;
            end
            begin
              rf_driver[27][11].run()  ;
            end

            begin
              gen[27][12].run()  ;
            end
            begin
              drv[27][12].run()  ;
            end
            begin
              mem_check[27][12].run()  ;
            end
            begin
              rf_driver[27][12].run()  ;
            end

            begin
              gen[27][13].run()  ;
            end
            begin
              drv[27][13].run()  ;
            end
            begin
              mem_check[27][13].run()  ;
            end
            begin
              rf_driver[27][13].run()  ;
            end

            begin
              gen[27][14].run()  ;
            end
            begin
              drv[27][14].run()  ;
            end
            begin
              mem_check[27][14].run()  ;
            end
            begin
              rf_driver[27][14].run()  ;
            end

            begin
              gen[27][15].run()  ;
            end
            begin
              drv[27][15].run()  ;
            end
            begin
              mem_check[27][15].run()  ;
            end
            begin
              rf_driver[27][15].run()  ;
            end

            begin
              gen[27][16].run()  ;
            end
            begin
              drv[27][16].run()  ;
            end
            begin
              mem_check[27][16].run()  ;
            end
            begin
              rf_driver[27][16].run()  ;
            end

            begin
              gen[27][17].run()  ;
            end
            begin
              drv[27][17].run()  ;
            end
            begin
              mem_check[27][17].run()  ;
            end
            begin
              rf_driver[27][17].run()  ;
            end

            begin
              gen[27][18].run()  ;
            end
            begin
              drv[27][18].run()  ;
            end
            begin
              mem_check[27][18].run()  ;
            end
            begin
              rf_driver[27][18].run()  ;
            end

            begin
              gen[27][19].run()  ;
            end
            begin
              drv[27][19].run()  ;
            end
            begin
              mem_check[27][19].run()  ;
            end
            begin
              rf_driver[27][19].run()  ;
            end

            begin
              gen[27][20].run()  ;
            end
            begin
              drv[27][20].run()  ;
            end
            begin
              mem_check[27][20].run()  ;
            end
            begin
              rf_driver[27][20].run()  ;
            end

            begin
              gen[27][21].run()  ;
            end
            begin
              drv[27][21].run()  ;
            end
            begin
              mem_check[27][21].run()  ;
            end
            begin
              rf_driver[27][21].run()  ;
            end

            begin
              gen[27][22].run()  ;
            end
            begin
              drv[27][22].run()  ;
            end
            begin
              mem_check[27][22].run()  ;
            end
            begin
              rf_driver[27][22].run()  ;
            end

            begin
              gen[27][23].run()  ;
            end
            begin
              drv[27][23].run()  ;
            end
            begin
              mem_check[27][23].run()  ;
            end
            begin
              rf_driver[27][23].run()  ;
            end

            begin
              gen[27][24].run()  ;
            end
            begin
              drv[27][24].run()  ;
            end
            begin
              mem_check[27][24].run()  ;
            end
            begin
              rf_driver[27][24].run()  ;
            end

            begin
              gen[27][25].run()  ;
            end
            begin
              drv[27][25].run()  ;
            end
            begin
              mem_check[27][25].run()  ;
            end
            begin
              rf_driver[27][25].run()  ;
            end

            begin
              gen[27][26].run()  ;
            end
            begin
              drv[27][26].run()  ;
            end
            begin
              mem_check[27][26].run()  ;
            end
            begin
              rf_driver[27][26].run()  ;
            end

            begin
              gen[27][27].run()  ;
            end
            begin
              drv[27][27].run()  ;
            end
            begin
              mem_check[27][27].run()  ;
            end
            begin
              rf_driver[27][27].run()  ;
            end

            begin
              gen[27][28].run()  ;
            end
            begin
              drv[27][28].run()  ;
            end
            begin
              mem_check[27][28].run()  ;
            end
            begin
              rf_driver[27][28].run()  ;
            end

            begin
              gen[27][29].run()  ;
            end
            begin
              drv[27][29].run()  ;
            end
            begin
              mem_check[27][29].run()  ;
            end
            begin
              rf_driver[27][29].run()  ;
            end

            begin
              gen[27][30].run()  ;
            end
            begin
              drv[27][30].run()  ;
            end
            begin
              mem_check[27][30].run()  ;
            end
            begin
              rf_driver[27][30].run()  ;
            end

            begin
              gen[27][31].run()  ;
            end
            begin
              drv[27][31].run()  ;
            end
            begin
              mem_check[27][31].run()  ;
            end
            begin
              rf_driver[27][31].run()  ;
            end

            begin
              ldst_driver[28].run()  ;
            end
            begin
              mgr[28].run()  ;
            end
            begin
              oob_drv[28].run()  ;
            end
            begin
              up_check[28].run()  ;
            end
            begin
              gen[28][0].run()  ;
            end
            begin
              drv[28][0].run()  ;
            end
            begin
              mem_check[28][0].run()  ;
            end
            begin
              rf_driver[28][0].run()  ;
            end

            begin
              gen[28][1].run()  ;
            end
            begin
              drv[28][1].run()  ;
            end
            begin
              mem_check[28][1].run()  ;
            end
            begin
              rf_driver[28][1].run()  ;
            end

            begin
              gen[28][2].run()  ;
            end
            begin
              drv[28][2].run()  ;
            end
            begin
              mem_check[28][2].run()  ;
            end
            begin
              rf_driver[28][2].run()  ;
            end

            begin
              gen[28][3].run()  ;
            end
            begin
              drv[28][3].run()  ;
            end
            begin
              mem_check[28][3].run()  ;
            end
            begin
              rf_driver[28][3].run()  ;
            end

            begin
              gen[28][4].run()  ;
            end
            begin
              drv[28][4].run()  ;
            end
            begin
              mem_check[28][4].run()  ;
            end
            begin
              rf_driver[28][4].run()  ;
            end

            begin
              gen[28][5].run()  ;
            end
            begin
              drv[28][5].run()  ;
            end
            begin
              mem_check[28][5].run()  ;
            end
            begin
              rf_driver[28][5].run()  ;
            end

            begin
              gen[28][6].run()  ;
            end
            begin
              drv[28][6].run()  ;
            end
            begin
              mem_check[28][6].run()  ;
            end
            begin
              rf_driver[28][6].run()  ;
            end

            begin
              gen[28][7].run()  ;
            end
            begin
              drv[28][7].run()  ;
            end
            begin
              mem_check[28][7].run()  ;
            end
            begin
              rf_driver[28][7].run()  ;
            end

            begin
              gen[28][8].run()  ;
            end
            begin
              drv[28][8].run()  ;
            end
            begin
              mem_check[28][8].run()  ;
            end
            begin
              rf_driver[28][8].run()  ;
            end

            begin
              gen[28][9].run()  ;
            end
            begin
              drv[28][9].run()  ;
            end
            begin
              mem_check[28][9].run()  ;
            end
            begin
              rf_driver[28][9].run()  ;
            end

            begin
              gen[28][10].run()  ;
            end
            begin
              drv[28][10].run()  ;
            end
            begin
              mem_check[28][10].run()  ;
            end
            begin
              rf_driver[28][10].run()  ;
            end

            begin
              gen[28][11].run()  ;
            end
            begin
              drv[28][11].run()  ;
            end
            begin
              mem_check[28][11].run()  ;
            end
            begin
              rf_driver[28][11].run()  ;
            end

            begin
              gen[28][12].run()  ;
            end
            begin
              drv[28][12].run()  ;
            end
            begin
              mem_check[28][12].run()  ;
            end
            begin
              rf_driver[28][12].run()  ;
            end

            begin
              gen[28][13].run()  ;
            end
            begin
              drv[28][13].run()  ;
            end
            begin
              mem_check[28][13].run()  ;
            end
            begin
              rf_driver[28][13].run()  ;
            end

            begin
              gen[28][14].run()  ;
            end
            begin
              drv[28][14].run()  ;
            end
            begin
              mem_check[28][14].run()  ;
            end
            begin
              rf_driver[28][14].run()  ;
            end

            begin
              gen[28][15].run()  ;
            end
            begin
              drv[28][15].run()  ;
            end
            begin
              mem_check[28][15].run()  ;
            end
            begin
              rf_driver[28][15].run()  ;
            end

            begin
              gen[28][16].run()  ;
            end
            begin
              drv[28][16].run()  ;
            end
            begin
              mem_check[28][16].run()  ;
            end
            begin
              rf_driver[28][16].run()  ;
            end

            begin
              gen[28][17].run()  ;
            end
            begin
              drv[28][17].run()  ;
            end
            begin
              mem_check[28][17].run()  ;
            end
            begin
              rf_driver[28][17].run()  ;
            end

            begin
              gen[28][18].run()  ;
            end
            begin
              drv[28][18].run()  ;
            end
            begin
              mem_check[28][18].run()  ;
            end
            begin
              rf_driver[28][18].run()  ;
            end

            begin
              gen[28][19].run()  ;
            end
            begin
              drv[28][19].run()  ;
            end
            begin
              mem_check[28][19].run()  ;
            end
            begin
              rf_driver[28][19].run()  ;
            end

            begin
              gen[28][20].run()  ;
            end
            begin
              drv[28][20].run()  ;
            end
            begin
              mem_check[28][20].run()  ;
            end
            begin
              rf_driver[28][20].run()  ;
            end

            begin
              gen[28][21].run()  ;
            end
            begin
              drv[28][21].run()  ;
            end
            begin
              mem_check[28][21].run()  ;
            end
            begin
              rf_driver[28][21].run()  ;
            end

            begin
              gen[28][22].run()  ;
            end
            begin
              drv[28][22].run()  ;
            end
            begin
              mem_check[28][22].run()  ;
            end
            begin
              rf_driver[28][22].run()  ;
            end

            begin
              gen[28][23].run()  ;
            end
            begin
              drv[28][23].run()  ;
            end
            begin
              mem_check[28][23].run()  ;
            end
            begin
              rf_driver[28][23].run()  ;
            end

            begin
              gen[28][24].run()  ;
            end
            begin
              drv[28][24].run()  ;
            end
            begin
              mem_check[28][24].run()  ;
            end
            begin
              rf_driver[28][24].run()  ;
            end

            begin
              gen[28][25].run()  ;
            end
            begin
              drv[28][25].run()  ;
            end
            begin
              mem_check[28][25].run()  ;
            end
            begin
              rf_driver[28][25].run()  ;
            end

            begin
              gen[28][26].run()  ;
            end
            begin
              drv[28][26].run()  ;
            end
            begin
              mem_check[28][26].run()  ;
            end
            begin
              rf_driver[28][26].run()  ;
            end

            begin
              gen[28][27].run()  ;
            end
            begin
              drv[28][27].run()  ;
            end
            begin
              mem_check[28][27].run()  ;
            end
            begin
              rf_driver[28][27].run()  ;
            end

            begin
              gen[28][28].run()  ;
            end
            begin
              drv[28][28].run()  ;
            end
            begin
              mem_check[28][28].run()  ;
            end
            begin
              rf_driver[28][28].run()  ;
            end

            begin
              gen[28][29].run()  ;
            end
            begin
              drv[28][29].run()  ;
            end
            begin
              mem_check[28][29].run()  ;
            end
            begin
              rf_driver[28][29].run()  ;
            end

            begin
              gen[28][30].run()  ;
            end
            begin
              drv[28][30].run()  ;
            end
            begin
              mem_check[28][30].run()  ;
            end
            begin
              rf_driver[28][30].run()  ;
            end

            begin
              gen[28][31].run()  ;
            end
            begin
              drv[28][31].run()  ;
            end
            begin
              mem_check[28][31].run()  ;
            end
            begin
              rf_driver[28][31].run()  ;
            end

            begin
              ldst_driver[29].run()  ;
            end
            begin
              mgr[29].run()  ;
            end
            begin
              oob_drv[29].run()  ;
            end
            begin
              up_check[29].run()  ;
            end
            begin
              gen[29][0].run()  ;
            end
            begin
              drv[29][0].run()  ;
            end
            begin
              mem_check[29][0].run()  ;
            end
            begin
              rf_driver[29][0].run()  ;
            end

            begin
              gen[29][1].run()  ;
            end
            begin
              drv[29][1].run()  ;
            end
            begin
              mem_check[29][1].run()  ;
            end
            begin
              rf_driver[29][1].run()  ;
            end

            begin
              gen[29][2].run()  ;
            end
            begin
              drv[29][2].run()  ;
            end
            begin
              mem_check[29][2].run()  ;
            end
            begin
              rf_driver[29][2].run()  ;
            end

            begin
              gen[29][3].run()  ;
            end
            begin
              drv[29][3].run()  ;
            end
            begin
              mem_check[29][3].run()  ;
            end
            begin
              rf_driver[29][3].run()  ;
            end

            begin
              gen[29][4].run()  ;
            end
            begin
              drv[29][4].run()  ;
            end
            begin
              mem_check[29][4].run()  ;
            end
            begin
              rf_driver[29][4].run()  ;
            end

            begin
              gen[29][5].run()  ;
            end
            begin
              drv[29][5].run()  ;
            end
            begin
              mem_check[29][5].run()  ;
            end
            begin
              rf_driver[29][5].run()  ;
            end

            begin
              gen[29][6].run()  ;
            end
            begin
              drv[29][6].run()  ;
            end
            begin
              mem_check[29][6].run()  ;
            end
            begin
              rf_driver[29][6].run()  ;
            end

            begin
              gen[29][7].run()  ;
            end
            begin
              drv[29][7].run()  ;
            end
            begin
              mem_check[29][7].run()  ;
            end
            begin
              rf_driver[29][7].run()  ;
            end

            begin
              gen[29][8].run()  ;
            end
            begin
              drv[29][8].run()  ;
            end
            begin
              mem_check[29][8].run()  ;
            end
            begin
              rf_driver[29][8].run()  ;
            end

            begin
              gen[29][9].run()  ;
            end
            begin
              drv[29][9].run()  ;
            end
            begin
              mem_check[29][9].run()  ;
            end
            begin
              rf_driver[29][9].run()  ;
            end

            begin
              gen[29][10].run()  ;
            end
            begin
              drv[29][10].run()  ;
            end
            begin
              mem_check[29][10].run()  ;
            end
            begin
              rf_driver[29][10].run()  ;
            end

            begin
              gen[29][11].run()  ;
            end
            begin
              drv[29][11].run()  ;
            end
            begin
              mem_check[29][11].run()  ;
            end
            begin
              rf_driver[29][11].run()  ;
            end

            begin
              gen[29][12].run()  ;
            end
            begin
              drv[29][12].run()  ;
            end
            begin
              mem_check[29][12].run()  ;
            end
            begin
              rf_driver[29][12].run()  ;
            end

            begin
              gen[29][13].run()  ;
            end
            begin
              drv[29][13].run()  ;
            end
            begin
              mem_check[29][13].run()  ;
            end
            begin
              rf_driver[29][13].run()  ;
            end

            begin
              gen[29][14].run()  ;
            end
            begin
              drv[29][14].run()  ;
            end
            begin
              mem_check[29][14].run()  ;
            end
            begin
              rf_driver[29][14].run()  ;
            end

            begin
              gen[29][15].run()  ;
            end
            begin
              drv[29][15].run()  ;
            end
            begin
              mem_check[29][15].run()  ;
            end
            begin
              rf_driver[29][15].run()  ;
            end

            begin
              gen[29][16].run()  ;
            end
            begin
              drv[29][16].run()  ;
            end
            begin
              mem_check[29][16].run()  ;
            end
            begin
              rf_driver[29][16].run()  ;
            end

            begin
              gen[29][17].run()  ;
            end
            begin
              drv[29][17].run()  ;
            end
            begin
              mem_check[29][17].run()  ;
            end
            begin
              rf_driver[29][17].run()  ;
            end

            begin
              gen[29][18].run()  ;
            end
            begin
              drv[29][18].run()  ;
            end
            begin
              mem_check[29][18].run()  ;
            end
            begin
              rf_driver[29][18].run()  ;
            end

            begin
              gen[29][19].run()  ;
            end
            begin
              drv[29][19].run()  ;
            end
            begin
              mem_check[29][19].run()  ;
            end
            begin
              rf_driver[29][19].run()  ;
            end

            begin
              gen[29][20].run()  ;
            end
            begin
              drv[29][20].run()  ;
            end
            begin
              mem_check[29][20].run()  ;
            end
            begin
              rf_driver[29][20].run()  ;
            end

            begin
              gen[29][21].run()  ;
            end
            begin
              drv[29][21].run()  ;
            end
            begin
              mem_check[29][21].run()  ;
            end
            begin
              rf_driver[29][21].run()  ;
            end

            begin
              gen[29][22].run()  ;
            end
            begin
              drv[29][22].run()  ;
            end
            begin
              mem_check[29][22].run()  ;
            end
            begin
              rf_driver[29][22].run()  ;
            end

            begin
              gen[29][23].run()  ;
            end
            begin
              drv[29][23].run()  ;
            end
            begin
              mem_check[29][23].run()  ;
            end
            begin
              rf_driver[29][23].run()  ;
            end

            begin
              gen[29][24].run()  ;
            end
            begin
              drv[29][24].run()  ;
            end
            begin
              mem_check[29][24].run()  ;
            end
            begin
              rf_driver[29][24].run()  ;
            end

            begin
              gen[29][25].run()  ;
            end
            begin
              drv[29][25].run()  ;
            end
            begin
              mem_check[29][25].run()  ;
            end
            begin
              rf_driver[29][25].run()  ;
            end

            begin
              gen[29][26].run()  ;
            end
            begin
              drv[29][26].run()  ;
            end
            begin
              mem_check[29][26].run()  ;
            end
            begin
              rf_driver[29][26].run()  ;
            end

            begin
              gen[29][27].run()  ;
            end
            begin
              drv[29][27].run()  ;
            end
            begin
              mem_check[29][27].run()  ;
            end
            begin
              rf_driver[29][27].run()  ;
            end

            begin
              gen[29][28].run()  ;
            end
            begin
              drv[29][28].run()  ;
            end
            begin
              mem_check[29][28].run()  ;
            end
            begin
              rf_driver[29][28].run()  ;
            end

            begin
              gen[29][29].run()  ;
            end
            begin
              drv[29][29].run()  ;
            end
            begin
              mem_check[29][29].run()  ;
            end
            begin
              rf_driver[29][29].run()  ;
            end

            begin
              gen[29][30].run()  ;
            end
            begin
              drv[29][30].run()  ;
            end
            begin
              mem_check[29][30].run()  ;
            end
            begin
              rf_driver[29][30].run()  ;
            end

            begin
              gen[29][31].run()  ;
            end
            begin
              drv[29][31].run()  ;
            end
            begin
              mem_check[29][31].run()  ;
            end
            begin
              rf_driver[29][31].run()  ;
            end

            begin
              ldst_driver[30].run()  ;
            end
            begin
              mgr[30].run()  ;
            end
            begin
              oob_drv[30].run()  ;
            end
            begin
              up_check[30].run()  ;
            end
            begin
              gen[30][0].run()  ;
            end
            begin
              drv[30][0].run()  ;
            end
            begin
              mem_check[30][0].run()  ;
            end
            begin
              rf_driver[30][0].run()  ;
            end

            begin
              gen[30][1].run()  ;
            end
            begin
              drv[30][1].run()  ;
            end
            begin
              mem_check[30][1].run()  ;
            end
            begin
              rf_driver[30][1].run()  ;
            end

            begin
              gen[30][2].run()  ;
            end
            begin
              drv[30][2].run()  ;
            end
            begin
              mem_check[30][2].run()  ;
            end
            begin
              rf_driver[30][2].run()  ;
            end

            begin
              gen[30][3].run()  ;
            end
            begin
              drv[30][3].run()  ;
            end
            begin
              mem_check[30][3].run()  ;
            end
            begin
              rf_driver[30][3].run()  ;
            end

            begin
              gen[30][4].run()  ;
            end
            begin
              drv[30][4].run()  ;
            end
            begin
              mem_check[30][4].run()  ;
            end
            begin
              rf_driver[30][4].run()  ;
            end

            begin
              gen[30][5].run()  ;
            end
            begin
              drv[30][5].run()  ;
            end
            begin
              mem_check[30][5].run()  ;
            end
            begin
              rf_driver[30][5].run()  ;
            end

            begin
              gen[30][6].run()  ;
            end
            begin
              drv[30][6].run()  ;
            end
            begin
              mem_check[30][6].run()  ;
            end
            begin
              rf_driver[30][6].run()  ;
            end

            begin
              gen[30][7].run()  ;
            end
            begin
              drv[30][7].run()  ;
            end
            begin
              mem_check[30][7].run()  ;
            end
            begin
              rf_driver[30][7].run()  ;
            end

            begin
              gen[30][8].run()  ;
            end
            begin
              drv[30][8].run()  ;
            end
            begin
              mem_check[30][8].run()  ;
            end
            begin
              rf_driver[30][8].run()  ;
            end

            begin
              gen[30][9].run()  ;
            end
            begin
              drv[30][9].run()  ;
            end
            begin
              mem_check[30][9].run()  ;
            end
            begin
              rf_driver[30][9].run()  ;
            end

            begin
              gen[30][10].run()  ;
            end
            begin
              drv[30][10].run()  ;
            end
            begin
              mem_check[30][10].run()  ;
            end
            begin
              rf_driver[30][10].run()  ;
            end

            begin
              gen[30][11].run()  ;
            end
            begin
              drv[30][11].run()  ;
            end
            begin
              mem_check[30][11].run()  ;
            end
            begin
              rf_driver[30][11].run()  ;
            end

            begin
              gen[30][12].run()  ;
            end
            begin
              drv[30][12].run()  ;
            end
            begin
              mem_check[30][12].run()  ;
            end
            begin
              rf_driver[30][12].run()  ;
            end

            begin
              gen[30][13].run()  ;
            end
            begin
              drv[30][13].run()  ;
            end
            begin
              mem_check[30][13].run()  ;
            end
            begin
              rf_driver[30][13].run()  ;
            end

            begin
              gen[30][14].run()  ;
            end
            begin
              drv[30][14].run()  ;
            end
            begin
              mem_check[30][14].run()  ;
            end
            begin
              rf_driver[30][14].run()  ;
            end

            begin
              gen[30][15].run()  ;
            end
            begin
              drv[30][15].run()  ;
            end
            begin
              mem_check[30][15].run()  ;
            end
            begin
              rf_driver[30][15].run()  ;
            end

            begin
              gen[30][16].run()  ;
            end
            begin
              drv[30][16].run()  ;
            end
            begin
              mem_check[30][16].run()  ;
            end
            begin
              rf_driver[30][16].run()  ;
            end

            begin
              gen[30][17].run()  ;
            end
            begin
              drv[30][17].run()  ;
            end
            begin
              mem_check[30][17].run()  ;
            end
            begin
              rf_driver[30][17].run()  ;
            end

            begin
              gen[30][18].run()  ;
            end
            begin
              drv[30][18].run()  ;
            end
            begin
              mem_check[30][18].run()  ;
            end
            begin
              rf_driver[30][18].run()  ;
            end

            begin
              gen[30][19].run()  ;
            end
            begin
              drv[30][19].run()  ;
            end
            begin
              mem_check[30][19].run()  ;
            end
            begin
              rf_driver[30][19].run()  ;
            end

            begin
              gen[30][20].run()  ;
            end
            begin
              drv[30][20].run()  ;
            end
            begin
              mem_check[30][20].run()  ;
            end
            begin
              rf_driver[30][20].run()  ;
            end

            begin
              gen[30][21].run()  ;
            end
            begin
              drv[30][21].run()  ;
            end
            begin
              mem_check[30][21].run()  ;
            end
            begin
              rf_driver[30][21].run()  ;
            end

            begin
              gen[30][22].run()  ;
            end
            begin
              drv[30][22].run()  ;
            end
            begin
              mem_check[30][22].run()  ;
            end
            begin
              rf_driver[30][22].run()  ;
            end

            begin
              gen[30][23].run()  ;
            end
            begin
              drv[30][23].run()  ;
            end
            begin
              mem_check[30][23].run()  ;
            end
            begin
              rf_driver[30][23].run()  ;
            end

            begin
              gen[30][24].run()  ;
            end
            begin
              drv[30][24].run()  ;
            end
            begin
              mem_check[30][24].run()  ;
            end
            begin
              rf_driver[30][24].run()  ;
            end

            begin
              gen[30][25].run()  ;
            end
            begin
              drv[30][25].run()  ;
            end
            begin
              mem_check[30][25].run()  ;
            end
            begin
              rf_driver[30][25].run()  ;
            end

            begin
              gen[30][26].run()  ;
            end
            begin
              drv[30][26].run()  ;
            end
            begin
              mem_check[30][26].run()  ;
            end
            begin
              rf_driver[30][26].run()  ;
            end

            begin
              gen[30][27].run()  ;
            end
            begin
              drv[30][27].run()  ;
            end
            begin
              mem_check[30][27].run()  ;
            end
            begin
              rf_driver[30][27].run()  ;
            end

            begin
              gen[30][28].run()  ;
            end
            begin
              drv[30][28].run()  ;
            end
            begin
              mem_check[30][28].run()  ;
            end
            begin
              rf_driver[30][28].run()  ;
            end

            begin
              gen[30][29].run()  ;
            end
            begin
              drv[30][29].run()  ;
            end
            begin
              mem_check[30][29].run()  ;
            end
            begin
              rf_driver[30][29].run()  ;
            end

            begin
              gen[30][30].run()  ;
            end
            begin
              drv[30][30].run()  ;
            end
            begin
              mem_check[30][30].run()  ;
            end
            begin
              rf_driver[30][30].run()  ;
            end

            begin
              gen[30][31].run()  ;
            end
            begin
              drv[30][31].run()  ;
            end
            begin
              mem_check[30][31].run()  ;
            end
            begin
              rf_driver[30][31].run()  ;
            end

            begin
              ldst_driver[31].run()  ;
            end
            begin
              mgr[31].run()  ;
            end
            begin
              oob_drv[31].run()  ;
            end
            begin
              up_check[31].run()  ;
            end
            begin
              gen[31][0].run()  ;
            end
            begin
              drv[31][0].run()  ;
            end
            begin
              mem_check[31][0].run()  ;
            end
            begin
              rf_driver[31][0].run()  ;
            end

            begin
              gen[31][1].run()  ;
            end
            begin
              drv[31][1].run()  ;
            end
            begin
              mem_check[31][1].run()  ;
            end
            begin
              rf_driver[31][1].run()  ;
            end

            begin
              gen[31][2].run()  ;
            end
            begin
              drv[31][2].run()  ;
            end
            begin
              mem_check[31][2].run()  ;
            end
            begin
              rf_driver[31][2].run()  ;
            end

            begin
              gen[31][3].run()  ;
            end
            begin
              drv[31][3].run()  ;
            end
            begin
              mem_check[31][3].run()  ;
            end
            begin
              rf_driver[31][3].run()  ;
            end

            begin
              gen[31][4].run()  ;
            end
            begin
              drv[31][4].run()  ;
            end
            begin
              mem_check[31][4].run()  ;
            end
            begin
              rf_driver[31][4].run()  ;
            end

            begin
              gen[31][5].run()  ;
            end
            begin
              drv[31][5].run()  ;
            end
            begin
              mem_check[31][5].run()  ;
            end
            begin
              rf_driver[31][5].run()  ;
            end

            begin
              gen[31][6].run()  ;
            end
            begin
              drv[31][6].run()  ;
            end
            begin
              mem_check[31][6].run()  ;
            end
            begin
              rf_driver[31][6].run()  ;
            end

            begin
              gen[31][7].run()  ;
            end
            begin
              drv[31][7].run()  ;
            end
            begin
              mem_check[31][7].run()  ;
            end
            begin
              rf_driver[31][7].run()  ;
            end

            begin
              gen[31][8].run()  ;
            end
            begin
              drv[31][8].run()  ;
            end
            begin
              mem_check[31][8].run()  ;
            end
            begin
              rf_driver[31][8].run()  ;
            end

            begin
              gen[31][9].run()  ;
            end
            begin
              drv[31][9].run()  ;
            end
            begin
              mem_check[31][9].run()  ;
            end
            begin
              rf_driver[31][9].run()  ;
            end

            begin
              gen[31][10].run()  ;
            end
            begin
              drv[31][10].run()  ;
            end
            begin
              mem_check[31][10].run()  ;
            end
            begin
              rf_driver[31][10].run()  ;
            end

            begin
              gen[31][11].run()  ;
            end
            begin
              drv[31][11].run()  ;
            end
            begin
              mem_check[31][11].run()  ;
            end
            begin
              rf_driver[31][11].run()  ;
            end

            begin
              gen[31][12].run()  ;
            end
            begin
              drv[31][12].run()  ;
            end
            begin
              mem_check[31][12].run()  ;
            end
            begin
              rf_driver[31][12].run()  ;
            end

            begin
              gen[31][13].run()  ;
            end
            begin
              drv[31][13].run()  ;
            end
            begin
              mem_check[31][13].run()  ;
            end
            begin
              rf_driver[31][13].run()  ;
            end

            begin
              gen[31][14].run()  ;
            end
            begin
              drv[31][14].run()  ;
            end
            begin
              mem_check[31][14].run()  ;
            end
            begin
              rf_driver[31][14].run()  ;
            end

            begin
              gen[31][15].run()  ;
            end
            begin
              drv[31][15].run()  ;
            end
            begin
              mem_check[31][15].run()  ;
            end
            begin
              rf_driver[31][15].run()  ;
            end

            begin
              gen[31][16].run()  ;
            end
            begin
              drv[31][16].run()  ;
            end
            begin
              mem_check[31][16].run()  ;
            end
            begin
              rf_driver[31][16].run()  ;
            end

            begin
              gen[31][17].run()  ;
            end
            begin
              drv[31][17].run()  ;
            end
            begin
              mem_check[31][17].run()  ;
            end
            begin
              rf_driver[31][17].run()  ;
            end

            begin
              gen[31][18].run()  ;
            end
            begin
              drv[31][18].run()  ;
            end
            begin
              mem_check[31][18].run()  ;
            end
            begin
              rf_driver[31][18].run()  ;
            end

            begin
              gen[31][19].run()  ;
            end
            begin
              drv[31][19].run()  ;
            end
            begin
              mem_check[31][19].run()  ;
            end
            begin
              rf_driver[31][19].run()  ;
            end

            begin
              gen[31][20].run()  ;
            end
            begin
              drv[31][20].run()  ;
            end
            begin
              mem_check[31][20].run()  ;
            end
            begin
              rf_driver[31][20].run()  ;
            end

            begin
              gen[31][21].run()  ;
            end
            begin
              drv[31][21].run()  ;
            end
            begin
              mem_check[31][21].run()  ;
            end
            begin
              rf_driver[31][21].run()  ;
            end

            begin
              gen[31][22].run()  ;
            end
            begin
              drv[31][22].run()  ;
            end
            begin
              mem_check[31][22].run()  ;
            end
            begin
              rf_driver[31][22].run()  ;
            end

            begin
              gen[31][23].run()  ;
            end
            begin
              drv[31][23].run()  ;
            end
            begin
              mem_check[31][23].run()  ;
            end
            begin
              rf_driver[31][23].run()  ;
            end

            begin
              gen[31][24].run()  ;
            end
            begin
              drv[31][24].run()  ;
            end
            begin
              mem_check[31][24].run()  ;
            end
            begin
              rf_driver[31][24].run()  ;
            end

            begin
              gen[31][25].run()  ;
            end
            begin
              drv[31][25].run()  ;
            end
            begin
              mem_check[31][25].run()  ;
            end
            begin
              rf_driver[31][25].run()  ;
            end

            begin
              gen[31][26].run()  ;
            end
            begin
              drv[31][26].run()  ;
            end
            begin
              mem_check[31][26].run()  ;
            end
            begin
              rf_driver[31][26].run()  ;
            end

            begin
              gen[31][27].run()  ;
            end
            begin
              drv[31][27].run()  ;
            end
            begin
              mem_check[31][27].run()  ;
            end
            begin
              rf_driver[31][27].run()  ;
            end

            begin
              gen[31][28].run()  ;
            end
            begin
              drv[31][28].run()  ;
            end
            begin
              mem_check[31][28].run()  ;
            end
            begin
              rf_driver[31][28].run()  ;
            end

            begin
              gen[31][29].run()  ;
            end
            begin
              drv[31][29].run()  ;
            end
            begin
              mem_check[31][29].run()  ;
            end
            begin
              rf_driver[31][29].run()  ;
            end

            begin
              gen[31][30].run()  ;
            end
            begin
              drv[31][30].run()  ;
            end
            begin
              mem_check[31][30].run()  ;
            end
            begin
              rf_driver[31][30].run()  ;
            end

            begin
              gen[31][31].run()  ;
            end
            begin
              drv[31][31].run()  ;
            end
            begin
              mem_check[31][31].run()  ;
            end
            begin
              rf_driver[31][31].run()  ;
            end

            begin
              ldst_driver[32].run()  ;
            end
            begin
              mgr[32].run()  ;
            end
            begin
              oob_drv[32].run()  ;
            end
            begin
              up_check[32].run()  ;
            end
            begin
              gen[32][0].run()  ;
            end
            begin
              drv[32][0].run()  ;
            end
            begin
              mem_check[32][0].run()  ;
            end
            begin
              rf_driver[32][0].run()  ;
            end

            begin
              gen[32][1].run()  ;
            end
            begin
              drv[32][1].run()  ;
            end
            begin
              mem_check[32][1].run()  ;
            end
            begin
              rf_driver[32][1].run()  ;
            end

            begin
              gen[32][2].run()  ;
            end
            begin
              drv[32][2].run()  ;
            end
            begin
              mem_check[32][2].run()  ;
            end
            begin
              rf_driver[32][2].run()  ;
            end

            begin
              gen[32][3].run()  ;
            end
            begin
              drv[32][3].run()  ;
            end
            begin
              mem_check[32][3].run()  ;
            end
            begin
              rf_driver[32][3].run()  ;
            end

            begin
              gen[32][4].run()  ;
            end
            begin
              drv[32][4].run()  ;
            end
            begin
              mem_check[32][4].run()  ;
            end
            begin
              rf_driver[32][4].run()  ;
            end

            begin
              gen[32][5].run()  ;
            end
            begin
              drv[32][5].run()  ;
            end
            begin
              mem_check[32][5].run()  ;
            end
            begin
              rf_driver[32][5].run()  ;
            end

            begin
              gen[32][6].run()  ;
            end
            begin
              drv[32][6].run()  ;
            end
            begin
              mem_check[32][6].run()  ;
            end
            begin
              rf_driver[32][6].run()  ;
            end

            begin
              gen[32][7].run()  ;
            end
            begin
              drv[32][7].run()  ;
            end
            begin
              mem_check[32][7].run()  ;
            end
            begin
              rf_driver[32][7].run()  ;
            end

            begin
              gen[32][8].run()  ;
            end
            begin
              drv[32][8].run()  ;
            end
            begin
              mem_check[32][8].run()  ;
            end
            begin
              rf_driver[32][8].run()  ;
            end

            begin
              gen[32][9].run()  ;
            end
            begin
              drv[32][9].run()  ;
            end
            begin
              mem_check[32][9].run()  ;
            end
            begin
              rf_driver[32][9].run()  ;
            end

            begin
              gen[32][10].run()  ;
            end
            begin
              drv[32][10].run()  ;
            end
            begin
              mem_check[32][10].run()  ;
            end
            begin
              rf_driver[32][10].run()  ;
            end

            begin
              gen[32][11].run()  ;
            end
            begin
              drv[32][11].run()  ;
            end
            begin
              mem_check[32][11].run()  ;
            end
            begin
              rf_driver[32][11].run()  ;
            end

            begin
              gen[32][12].run()  ;
            end
            begin
              drv[32][12].run()  ;
            end
            begin
              mem_check[32][12].run()  ;
            end
            begin
              rf_driver[32][12].run()  ;
            end

            begin
              gen[32][13].run()  ;
            end
            begin
              drv[32][13].run()  ;
            end
            begin
              mem_check[32][13].run()  ;
            end
            begin
              rf_driver[32][13].run()  ;
            end

            begin
              gen[32][14].run()  ;
            end
            begin
              drv[32][14].run()  ;
            end
            begin
              mem_check[32][14].run()  ;
            end
            begin
              rf_driver[32][14].run()  ;
            end

            begin
              gen[32][15].run()  ;
            end
            begin
              drv[32][15].run()  ;
            end
            begin
              mem_check[32][15].run()  ;
            end
            begin
              rf_driver[32][15].run()  ;
            end

            begin
              gen[32][16].run()  ;
            end
            begin
              drv[32][16].run()  ;
            end
            begin
              mem_check[32][16].run()  ;
            end
            begin
              rf_driver[32][16].run()  ;
            end

            begin
              gen[32][17].run()  ;
            end
            begin
              drv[32][17].run()  ;
            end
            begin
              mem_check[32][17].run()  ;
            end
            begin
              rf_driver[32][17].run()  ;
            end

            begin
              gen[32][18].run()  ;
            end
            begin
              drv[32][18].run()  ;
            end
            begin
              mem_check[32][18].run()  ;
            end
            begin
              rf_driver[32][18].run()  ;
            end

            begin
              gen[32][19].run()  ;
            end
            begin
              drv[32][19].run()  ;
            end
            begin
              mem_check[32][19].run()  ;
            end
            begin
              rf_driver[32][19].run()  ;
            end

            begin
              gen[32][20].run()  ;
            end
            begin
              drv[32][20].run()  ;
            end
            begin
              mem_check[32][20].run()  ;
            end
            begin
              rf_driver[32][20].run()  ;
            end

            begin
              gen[32][21].run()  ;
            end
            begin
              drv[32][21].run()  ;
            end
            begin
              mem_check[32][21].run()  ;
            end
            begin
              rf_driver[32][21].run()  ;
            end

            begin
              gen[32][22].run()  ;
            end
            begin
              drv[32][22].run()  ;
            end
            begin
              mem_check[32][22].run()  ;
            end
            begin
              rf_driver[32][22].run()  ;
            end

            begin
              gen[32][23].run()  ;
            end
            begin
              drv[32][23].run()  ;
            end
            begin
              mem_check[32][23].run()  ;
            end
            begin
              rf_driver[32][23].run()  ;
            end

            begin
              gen[32][24].run()  ;
            end
            begin
              drv[32][24].run()  ;
            end
            begin
              mem_check[32][24].run()  ;
            end
            begin
              rf_driver[32][24].run()  ;
            end

            begin
              gen[32][25].run()  ;
            end
            begin
              drv[32][25].run()  ;
            end
            begin
              mem_check[32][25].run()  ;
            end
            begin
              rf_driver[32][25].run()  ;
            end

            begin
              gen[32][26].run()  ;
            end
            begin
              drv[32][26].run()  ;
            end
            begin
              mem_check[32][26].run()  ;
            end
            begin
              rf_driver[32][26].run()  ;
            end

            begin
              gen[32][27].run()  ;
            end
            begin
              drv[32][27].run()  ;
            end
            begin
              mem_check[32][27].run()  ;
            end
            begin
              rf_driver[32][27].run()  ;
            end

            begin
              gen[32][28].run()  ;
            end
            begin
              drv[32][28].run()  ;
            end
            begin
              mem_check[32][28].run()  ;
            end
            begin
              rf_driver[32][28].run()  ;
            end

            begin
              gen[32][29].run()  ;
            end
            begin
              drv[32][29].run()  ;
            end
            begin
              mem_check[32][29].run()  ;
            end
            begin
              rf_driver[32][29].run()  ;
            end

            begin
              gen[32][30].run()  ;
            end
            begin
              drv[32][30].run()  ;
            end
            begin
              mem_check[32][30].run()  ;
            end
            begin
              rf_driver[32][30].run()  ;
            end

            begin
              gen[32][31].run()  ;
            end
            begin
              drv[32][31].run()  ;
            end
            begin
              mem_check[32][31].run()  ;
            end
            begin
              rf_driver[32][31].run()  ;
            end

            begin
              ldst_driver[33].run()  ;
            end
            begin
              mgr[33].run()  ;
            end
            begin
              oob_drv[33].run()  ;
            end
            begin
              up_check[33].run()  ;
            end
            begin
              gen[33][0].run()  ;
            end
            begin
              drv[33][0].run()  ;
            end
            begin
              mem_check[33][0].run()  ;
            end
            begin
              rf_driver[33][0].run()  ;
            end

            begin
              gen[33][1].run()  ;
            end
            begin
              drv[33][1].run()  ;
            end
            begin
              mem_check[33][1].run()  ;
            end
            begin
              rf_driver[33][1].run()  ;
            end

            begin
              gen[33][2].run()  ;
            end
            begin
              drv[33][2].run()  ;
            end
            begin
              mem_check[33][2].run()  ;
            end
            begin
              rf_driver[33][2].run()  ;
            end

            begin
              gen[33][3].run()  ;
            end
            begin
              drv[33][3].run()  ;
            end
            begin
              mem_check[33][3].run()  ;
            end
            begin
              rf_driver[33][3].run()  ;
            end

            begin
              gen[33][4].run()  ;
            end
            begin
              drv[33][4].run()  ;
            end
            begin
              mem_check[33][4].run()  ;
            end
            begin
              rf_driver[33][4].run()  ;
            end

            begin
              gen[33][5].run()  ;
            end
            begin
              drv[33][5].run()  ;
            end
            begin
              mem_check[33][5].run()  ;
            end
            begin
              rf_driver[33][5].run()  ;
            end

            begin
              gen[33][6].run()  ;
            end
            begin
              drv[33][6].run()  ;
            end
            begin
              mem_check[33][6].run()  ;
            end
            begin
              rf_driver[33][6].run()  ;
            end

            begin
              gen[33][7].run()  ;
            end
            begin
              drv[33][7].run()  ;
            end
            begin
              mem_check[33][7].run()  ;
            end
            begin
              rf_driver[33][7].run()  ;
            end

            begin
              gen[33][8].run()  ;
            end
            begin
              drv[33][8].run()  ;
            end
            begin
              mem_check[33][8].run()  ;
            end
            begin
              rf_driver[33][8].run()  ;
            end

            begin
              gen[33][9].run()  ;
            end
            begin
              drv[33][9].run()  ;
            end
            begin
              mem_check[33][9].run()  ;
            end
            begin
              rf_driver[33][9].run()  ;
            end

            begin
              gen[33][10].run()  ;
            end
            begin
              drv[33][10].run()  ;
            end
            begin
              mem_check[33][10].run()  ;
            end
            begin
              rf_driver[33][10].run()  ;
            end

            begin
              gen[33][11].run()  ;
            end
            begin
              drv[33][11].run()  ;
            end
            begin
              mem_check[33][11].run()  ;
            end
            begin
              rf_driver[33][11].run()  ;
            end

            begin
              gen[33][12].run()  ;
            end
            begin
              drv[33][12].run()  ;
            end
            begin
              mem_check[33][12].run()  ;
            end
            begin
              rf_driver[33][12].run()  ;
            end

            begin
              gen[33][13].run()  ;
            end
            begin
              drv[33][13].run()  ;
            end
            begin
              mem_check[33][13].run()  ;
            end
            begin
              rf_driver[33][13].run()  ;
            end

            begin
              gen[33][14].run()  ;
            end
            begin
              drv[33][14].run()  ;
            end
            begin
              mem_check[33][14].run()  ;
            end
            begin
              rf_driver[33][14].run()  ;
            end

            begin
              gen[33][15].run()  ;
            end
            begin
              drv[33][15].run()  ;
            end
            begin
              mem_check[33][15].run()  ;
            end
            begin
              rf_driver[33][15].run()  ;
            end

            begin
              gen[33][16].run()  ;
            end
            begin
              drv[33][16].run()  ;
            end
            begin
              mem_check[33][16].run()  ;
            end
            begin
              rf_driver[33][16].run()  ;
            end

            begin
              gen[33][17].run()  ;
            end
            begin
              drv[33][17].run()  ;
            end
            begin
              mem_check[33][17].run()  ;
            end
            begin
              rf_driver[33][17].run()  ;
            end

            begin
              gen[33][18].run()  ;
            end
            begin
              drv[33][18].run()  ;
            end
            begin
              mem_check[33][18].run()  ;
            end
            begin
              rf_driver[33][18].run()  ;
            end

            begin
              gen[33][19].run()  ;
            end
            begin
              drv[33][19].run()  ;
            end
            begin
              mem_check[33][19].run()  ;
            end
            begin
              rf_driver[33][19].run()  ;
            end

            begin
              gen[33][20].run()  ;
            end
            begin
              drv[33][20].run()  ;
            end
            begin
              mem_check[33][20].run()  ;
            end
            begin
              rf_driver[33][20].run()  ;
            end

            begin
              gen[33][21].run()  ;
            end
            begin
              drv[33][21].run()  ;
            end
            begin
              mem_check[33][21].run()  ;
            end
            begin
              rf_driver[33][21].run()  ;
            end

            begin
              gen[33][22].run()  ;
            end
            begin
              drv[33][22].run()  ;
            end
            begin
              mem_check[33][22].run()  ;
            end
            begin
              rf_driver[33][22].run()  ;
            end

            begin
              gen[33][23].run()  ;
            end
            begin
              drv[33][23].run()  ;
            end
            begin
              mem_check[33][23].run()  ;
            end
            begin
              rf_driver[33][23].run()  ;
            end

            begin
              gen[33][24].run()  ;
            end
            begin
              drv[33][24].run()  ;
            end
            begin
              mem_check[33][24].run()  ;
            end
            begin
              rf_driver[33][24].run()  ;
            end

            begin
              gen[33][25].run()  ;
            end
            begin
              drv[33][25].run()  ;
            end
            begin
              mem_check[33][25].run()  ;
            end
            begin
              rf_driver[33][25].run()  ;
            end

            begin
              gen[33][26].run()  ;
            end
            begin
              drv[33][26].run()  ;
            end
            begin
              mem_check[33][26].run()  ;
            end
            begin
              rf_driver[33][26].run()  ;
            end

            begin
              gen[33][27].run()  ;
            end
            begin
              drv[33][27].run()  ;
            end
            begin
              mem_check[33][27].run()  ;
            end
            begin
              rf_driver[33][27].run()  ;
            end

            begin
              gen[33][28].run()  ;
            end
            begin
              drv[33][28].run()  ;
            end
            begin
              mem_check[33][28].run()  ;
            end
            begin
              rf_driver[33][28].run()  ;
            end

            begin
              gen[33][29].run()  ;
            end
            begin
              drv[33][29].run()  ;
            end
            begin
              mem_check[33][29].run()  ;
            end
            begin
              rf_driver[33][29].run()  ;
            end

            begin
              gen[33][30].run()  ;
            end
            begin
              drv[33][30].run()  ;
            end
            begin
              mem_check[33][30].run()  ;
            end
            begin
              rf_driver[33][30].run()  ;
            end

            begin
              gen[33][31].run()  ;
            end
            begin
              drv[33][31].run()  ;
            end
            begin
              mem_check[33][31].run()  ;
            end
            begin
              rf_driver[33][31].run()  ;
            end

            begin
              ldst_driver[34].run()  ;
            end
            begin
              mgr[34].run()  ;
            end
            begin
              oob_drv[34].run()  ;
            end
            begin
              up_check[34].run()  ;
            end
            begin
              gen[34][0].run()  ;
            end
            begin
              drv[34][0].run()  ;
            end
            begin
              mem_check[34][0].run()  ;
            end
            begin
              rf_driver[34][0].run()  ;
            end

            begin
              gen[34][1].run()  ;
            end
            begin
              drv[34][1].run()  ;
            end
            begin
              mem_check[34][1].run()  ;
            end
            begin
              rf_driver[34][1].run()  ;
            end

            begin
              gen[34][2].run()  ;
            end
            begin
              drv[34][2].run()  ;
            end
            begin
              mem_check[34][2].run()  ;
            end
            begin
              rf_driver[34][2].run()  ;
            end

            begin
              gen[34][3].run()  ;
            end
            begin
              drv[34][3].run()  ;
            end
            begin
              mem_check[34][3].run()  ;
            end
            begin
              rf_driver[34][3].run()  ;
            end

            begin
              gen[34][4].run()  ;
            end
            begin
              drv[34][4].run()  ;
            end
            begin
              mem_check[34][4].run()  ;
            end
            begin
              rf_driver[34][4].run()  ;
            end

            begin
              gen[34][5].run()  ;
            end
            begin
              drv[34][5].run()  ;
            end
            begin
              mem_check[34][5].run()  ;
            end
            begin
              rf_driver[34][5].run()  ;
            end

            begin
              gen[34][6].run()  ;
            end
            begin
              drv[34][6].run()  ;
            end
            begin
              mem_check[34][6].run()  ;
            end
            begin
              rf_driver[34][6].run()  ;
            end

            begin
              gen[34][7].run()  ;
            end
            begin
              drv[34][7].run()  ;
            end
            begin
              mem_check[34][7].run()  ;
            end
            begin
              rf_driver[34][7].run()  ;
            end

            begin
              gen[34][8].run()  ;
            end
            begin
              drv[34][8].run()  ;
            end
            begin
              mem_check[34][8].run()  ;
            end
            begin
              rf_driver[34][8].run()  ;
            end

            begin
              gen[34][9].run()  ;
            end
            begin
              drv[34][9].run()  ;
            end
            begin
              mem_check[34][9].run()  ;
            end
            begin
              rf_driver[34][9].run()  ;
            end

            begin
              gen[34][10].run()  ;
            end
            begin
              drv[34][10].run()  ;
            end
            begin
              mem_check[34][10].run()  ;
            end
            begin
              rf_driver[34][10].run()  ;
            end

            begin
              gen[34][11].run()  ;
            end
            begin
              drv[34][11].run()  ;
            end
            begin
              mem_check[34][11].run()  ;
            end
            begin
              rf_driver[34][11].run()  ;
            end

            begin
              gen[34][12].run()  ;
            end
            begin
              drv[34][12].run()  ;
            end
            begin
              mem_check[34][12].run()  ;
            end
            begin
              rf_driver[34][12].run()  ;
            end

            begin
              gen[34][13].run()  ;
            end
            begin
              drv[34][13].run()  ;
            end
            begin
              mem_check[34][13].run()  ;
            end
            begin
              rf_driver[34][13].run()  ;
            end

            begin
              gen[34][14].run()  ;
            end
            begin
              drv[34][14].run()  ;
            end
            begin
              mem_check[34][14].run()  ;
            end
            begin
              rf_driver[34][14].run()  ;
            end

            begin
              gen[34][15].run()  ;
            end
            begin
              drv[34][15].run()  ;
            end
            begin
              mem_check[34][15].run()  ;
            end
            begin
              rf_driver[34][15].run()  ;
            end

            begin
              gen[34][16].run()  ;
            end
            begin
              drv[34][16].run()  ;
            end
            begin
              mem_check[34][16].run()  ;
            end
            begin
              rf_driver[34][16].run()  ;
            end

            begin
              gen[34][17].run()  ;
            end
            begin
              drv[34][17].run()  ;
            end
            begin
              mem_check[34][17].run()  ;
            end
            begin
              rf_driver[34][17].run()  ;
            end

            begin
              gen[34][18].run()  ;
            end
            begin
              drv[34][18].run()  ;
            end
            begin
              mem_check[34][18].run()  ;
            end
            begin
              rf_driver[34][18].run()  ;
            end

            begin
              gen[34][19].run()  ;
            end
            begin
              drv[34][19].run()  ;
            end
            begin
              mem_check[34][19].run()  ;
            end
            begin
              rf_driver[34][19].run()  ;
            end

            begin
              gen[34][20].run()  ;
            end
            begin
              drv[34][20].run()  ;
            end
            begin
              mem_check[34][20].run()  ;
            end
            begin
              rf_driver[34][20].run()  ;
            end

            begin
              gen[34][21].run()  ;
            end
            begin
              drv[34][21].run()  ;
            end
            begin
              mem_check[34][21].run()  ;
            end
            begin
              rf_driver[34][21].run()  ;
            end

            begin
              gen[34][22].run()  ;
            end
            begin
              drv[34][22].run()  ;
            end
            begin
              mem_check[34][22].run()  ;
            end
            begin
              rf_driver[34][22].run()  ;
            end

            begin
              gen[34][23].run()  ;
            end
            begin
              drv[34][23].run()  ;
            end
            begin
              mem_check[34][23].run()  ;
            end
            begin
              rf_driver[34][23].run()  ;
            end

            begin
              gen[34][24].run()  ;
            end
            begin
              drv[34][24].run()  ;
            end
            begin
              mem_check[34][24].run()  ;
            end
            begin
              rf_driver[34][24].run()  ;
            end

            begin
              gen[34][25].run()  ;
            end
            begin
              drv[34][25].run()  ;
            end
            begin
              mem_check[34][25].run()  ;
            end
            begin
              rf_driver[34][25].run()  ;
            end

            begin
              gen[34][26].run()  ;
            end
            begin
              drv[34][26].run()  ;
            end
            begin
              mem_check[34][26].run()  ;
            end
            begin
              rf_driver[34][26].run()  ;
            end

            begin
              gen[34][27].run()  ;
            end
            begin
              drv[34][27].run()  ;
            end
            begin
              mem_check[34][27].run()  ;
            end
            begin
              rf_driver[34][27].run()  ;
            end

            begin
              gen[34][28].run()  ;
            end
            begin
              drv[34][28].run()  ;
            end
            begin
              mem_check[34][28].run()  ;
            end
            begin
              rf_driver[34][28].run()  ;
            end

            begin
              gen[34][29].run()  ;
            end
            begin
              drv[34][29].run()  ;
            end
            begin
              mem_check[34][29].run()  ;
            end
            begin
              rf_driver[34][29].run()  ;
            end

            begin
              gen[34][30].run()  ;
            end
            begin
              drv[34][30].run()  ;
            end
            begin
              mem_check[34][30].run()  ;
            end
            begin
              rf_driver[34][30].run()  ;
            end

            begin
              gen[34][31].run()  ;
            end
            begin
              drv[34][31].run()  ;
            end
            begin
              mem_check[34][31].run()  ;
            end
            begin
              rf_driver[34][31].run()  ;
            end

            begin
              ldst_driver[35].run()  ;
            end
            begin
              mgr[35].run()  ;
            end
            begin
              oob_drv[35].run()  ;
            end
            begin
              up_check[35].run()  ;
            end
            begin
              gen[35][0].run()  ;
            end
            begin
              drv[35][0].run()  ;
            end
            begin
              mem_check[35][0].run()  ;
            end
            begin
              rf_driver[35][0].run()  ;
            end

            begin
              gen[35][1].run()  ;
            end
            begin
              drv[35][1].run()  ;
            end
            begin
              mem_check[35][1].run()  ;
            end
            begin
              rf_driver[35][1].run()  ;
            end

            begin
              gen[35][2].run()  ;
            end
            begin
              drv[35][2].run()  ;
            end
            begin
              mem_check[35][2].run()  ;
            end
            begin
              rf_driver[35][2].run()  ;
            end

            begin
              gen[35][3].run()  ;
            end
            begin
              drv[35][3].run()  ;
            end
            begin
              mem_check[35][3].run()  ;
            end
            begin
              rf_driver[35][3].run()  ;
            end

            begin
              gen[35][4].run()  ;
            end
            begin
              drv[35][4].run()  ;
            end
            begin
              mem_check[35][4].run()  ;
            end
            begin
              rf_driver[35][4].run()  ;
            end

            begin
              gen[35][5].run()  ;
            end
            begin
              drv[35][5].run()  ;
            end
            begin
              mem_check[35][5].run()  ;
            end
            begin
              rf_driver[35][5].run()  ;
            end

            begin
              gen[35][6].run()  ;
            end
            begin
              drv[35][6].run()  ;
            end
            begin
              mem_check[35][6].run()  ;
            end
            begin
              rf_driver[35][6].run()  ;
            end

            begin
              gen[35][7].run()  ;
            end
            begin
              drv[35][7].run()  ;
            end
            begin
              mem_check[35][7].run()  ;
            end
            begin
              rf_driver[35][7].run()  ;
            end

            begin
              gen[35][8].run()  ;
            end
            begin
              drv[35][8].run()  ;
            end
            begin
              mem_check[35][8].run()  ;
            end
            begin
              rf_driver[35][8].run()  ;
            end

            begin
              gen[35][9].run()  ;
            end
            begin
              drv[35][9].run()  ;
            end
            begin
              mem_check[35][9].run()  ;
            end
            begin
              rf_driver[35][9].run()  ;
            end

            begin
              gen[35][10].run()  ;
            end
            begin
              drv[35][10].run()  ;
            end
            begin
              mem_check[35][10].run()  ;
            end
            begin
              rf_driver[35][10].run()  ;
            end

            begin
              gen[35][11].run()  ;
            end
            begin
              drv[35][11].run()  ;
            end
            begin
              mem_check[35][11].run()  ;
            end
            begin
              rf_driver[35][11].run()  ;
            end

            begin
              gen[35][12].run()  ;
            end
            begin
              drv[35][12].run()  ;
            end
            begin
              mem_check[35][12].run()  ;
            end
            begin
              rf_driver[35][12].run()  ;
            end

            begin
              gen[35][13].run()  ;
            end
            begin
              drv[35][13].run()  ;
            end
            begin
              mem_check[35][13].run()  ;
            end
            begin
              rf_driver[35][13].run()  ;
            end

            begin
              gen[35][14].run()  ;
            end
            begin
              drv[35][14].run()  ;
            end
            begin
              mem_check[35][14].run()  ;
            end
            begin
              rf_driver[35][14].run()  ;
            end

            begin
              gen[35][15].run()  ;
            end
            begin
              drv[35][15].run()  ;
            end
            begin
              mem_check[35][15].run()  ;
            end
            begin
              rf_driver[35][15].run()  ;
            end

            begin
              gen[35][16].run()  ;
            end
            begin
              drv[35][16].run()  ;
            end
            begin
              mem_check[35][16].run()  ;
            end
            begin
              rf_driver[35][16].run()  ;
            end

            begin
              gen[35][17].run()  ;
            end
            begin
              drv[35][17].run()  ;
            end
            begin
              mem_check[35][17].run()  ;
            end
            begin
              rf_driver[35][17].run()  ;
            end

            begin
              gen[35][18].run()  ;
            end
            begin
              drv[35][18].run()  ;
            end
            begin
              mem_check[35][18].run()  ;
            end
            begin
              rf_driver[35][18].run()  ;
            end

            begin
              gen[35][19].run()  ;
            end
            begin
              drv[35][19].run()  ;
            end
            begin
              mem_check[35][19].run()  ;
            end
            begin
              rf_driver[35][19].run()  ;
            end

            begin
              gen[35][20].run()  ;
            end
            begin
              drv[35][20].run()  ;
            end
            begin
              mem_check[35][20].run()  ;
            end
            begin
              rf_driver[35][20].run()  ;
            end

            begin
              gen[35][21].run()  ;
            end
            begin
              drv[35][21].run()  ;
            end
            begin
              mem_check[35][21].run()  ;
            end
            begin
              rf_driver[35][21].run()  ;
            end

            begin
              gen[35][22].run()  ;
            end
            begin
              drv[35][22].run()  ;
            end
            begin
              mem_check[35][22].run()  ;
            end
            begin
              rf_driver[35][22].run()  ;
            end

            begin
              gen[35][23].run()  ;
            end
            begin
              drv[35][23].run()  ;
            end
            begin
              mem_check[35][23].run()  ;
            end
            begin
              rf_driver[35][23].run()  ;
            end

            begin
              gen[35][24].run()  ;
            end
            begin
              drv[35][24].run()  ;
            end
            begin
              mem_check[35][24].run()  ;
            end
            begin
              rf_driver[35][24].run()  ;
            end

            begin
              gen[35][25].run()  ;
            end
            begin
              drv[35][25].run()  ;
            end
            begin
              mem_check[35][25].run()  ;
            end
            begin
              rf_driver[35][25].run()  ;
            end

            begin
              gen[35][26].run()  ;
            end
            begin
              drv[35][26].run()  ;
            end
            begin
              mem_check[35][26].run()  ;
            end
            begin
              rf_driver[35][26].run()  ;
            end

            begin
              gen[35][27].run()  ;
            end
            begin
              drv[35][27].run()  ;
            end
            begin
              mem_check[35][27].run()  ;
            end
            begin
              rf_driver[35][27].run()  ;
            end

            begin
              gen[35][28].run()  ;
            end
            begin
              drv[35][28].run()  ;
            end
            begin
              mem_check[35][28].run()  ;
            end
            begin
              rf_driver[35][28].run()  ;
            end

            begin
              gen[35][29].run()  ;
            end
            begin
              drv[35][29].run()  ;
            end
            begin
              mem_check[35][29].run()  ;
            end
            begin
              rf_driver[35][29].run()  ;
            end

            begin
              gen[35][30].run()  ;
            end
            begin
              drv[35][30].run()  ;
            end
            begin
              mem_check[35][30].run()  ;
            end
            begin
              rf_driver[35][30].run()  ;
            end

            begin
              gen[35][31].run()  ;
            end
            begin
              drv[35][31].run()  ;
            end
            begin
              mem_check[35][31].run()  ;
            end
            begin
              rf_driver[35][31].run()  ;
            end

            begin
              ldst_driver[36].run()  ;
            end
            begin
              mgr[36].run()  ;
            end
            begin
              oob_drv[36].run()  ;
            end
            begin
              up_check[36].run()  ;
            end
            begin
              gen[36][0].run()  ;
            end
            begin
              drv[36][0].run()  ;
            end
            begin
              mem_check[36][0].run()  ;
            end
            begin
              rf_driver[36][0].run()  ;
            end

            begin
              gen[36][1].run()  ;
            end
            begin
              drv[36][1].run()  ;
            end
            begin
              mem_check[36][1].run()  ;
            end
            begin
              rf_driver[36][1].run()  ;
            end

            begin
              gen[36][2].run()  ;
            end
            begin
              drv[36][2].run()  ;
            end
            begin
              mem_check[36][2].run()  ;
            end
            begin
              rf_driver[36][2].run()  ;
            end

            begin
              gen[36][3].run()  ;
            end
            begin
              drv[36][3].run()  ;
            end
            begin
              mem_check[36][3].run()  ;
            end
            begin
              rf_driver[36][3].run()  ;
            end

            begin
              gen[36][4].run()  ;
            end
            begin
              drv[36][4].run()  ;
            end
            begin
              mem_check[36][4].run()  ;
            end
            begin
              rf_driver[36][4].run()  ;
            end

            begin
              gen[36][5].run()  ;
            end
            begin
              drv[36][5].run()  ;
            end
            begin
              mem_check[36][5].run()  ;
            end
            begin
              rf_driver[36][5].run()  ;
            end

            begin
              gen[36][6].run()  ;
            end
            begin
              drv[36][6].run()  ;
            end
            begin
              mem_check[36][6].run()  ;
            end
            begin
              rf_driver[36][6].run()  ;
            end

            begin
              gen[36][7].run()  ;
            end
            begin
              drv[36][7].run()  ;
            end
            begin
              mem_check[36][7].run()  ;
            end
            begin
              rf_driver[36][7].run()  ;
            end

            begin
              gen[36][8].run()  ;
            end
            begin
              drv[36][8].run()  ;
            end
            begin
              mem_check[36][8].run()  ;
            end
            begin
              rf_driver[36][8].run()  ;
            end

            begin
              gen[36][9].run()  ;
            end
            begin
              drv[36][9].run()  ;
            end
            begin
              mem_check[36][9].run()  ;
            end
            begin
              rf_driver[36][9].run()  ;
            end

            begin
              gen[36][10].run()  ;
            end
            begin
              drv[36][10].run()  ;
            end
            begin
              mem_check[36][10].run()  ;
            end
            begin
              rf_driver[36][10].run()  ;
            end

            begin
              gen[36][11].run()  ;
            end
            begin
              drv[36][11].run()  ;
            end
            begin
              mem_check[36][11].run()  ;
            end
            begin
              rf_driver[36][11].run()  ;
            end

            begin
              gen[36][12].run()  ;
            end
            begin
              drv[36][12].run()  ;
            end
            begin
              mem_check[36][12].run()  ;
            end
            begin
              rf_driver[36][12].run()  ;
            end

            begin
              gen[36][13].run()  ;
            end
            begin
              drv[36][13].run()  ;
            end
            begin
              mem_check[36][13].run()  ;
            end
            begin
              rf_driver[36][13].run()  ;
            end

            begin
              gen[36][14].run()  ;
            end
            begin
              drv[36][14].run()  ;
            end
            begin
              mem_check[36][14].run()  ;
            end
            begin
              rf_driver[36][14].run()  ;
            end

            begin
              gen[36][15].run()  ;
            end
            begin
              drv[36][15].run()  ;
            end
            begin
              mem_check[36][15].run()  ;
            end
            begin
              rf_driver[36][15].run()  ;
            end

            begin
              gen[36][16].run()  ;
            end
            begin
              drv[36][16].run()  ;
            end
            begin
              mem_check[36][16].run()  ;
            end
            begin
              rf_driver[36][16].run()  ;
            end

            begin
              gen[36][17].run()  ;
            end
            begin
              drv[36][17].run()  ;
            end
            begin
              mem_check[36][17].run()  ;
            end
            begin
              rf_driver[36][17].run()  ;
            end

            begin
              gen[36][18].run()  ;
            end
            begin
              drv[36][18].run()  ;
            end
            begin
              mem_check[36][18].run()  ;
            end
            begin
              rf_driver[36][18].run()  ;
            end

            begin
              gen[36][19].run()  ;
            end
            begin
              drv[36][19].run()  ;
            end
            begin
              mem_check[36][19].run()  ;
            end
            begin
              rf_driver[36][19].run()  ;
            end

            begin
              gen[36][20].run()  ;
            end
            begin
              drv[36][20].run()  ;
            end
            begin
              mem_check[36][20].run()  ;
            end
            begin
              rf_driver[36][20].run()  ;
            end

            begin
              gen[36][21].run()  ;
            end
            begin
              drv[36][21].run()  ;
            end
            begin
              mem_check[36][21].run()  ;
            end
            begin
              rf_driver[36][21].run()  ;
            end

            begin
              gen[36][22].run()  ;
            end
            begin
              drv[36][22].run()  ;
            end
            begin
              mem_check[36][22].run()  ;
            end
            begin
              rf_driver[36][22].run()  ;
            end

            begin
              gen[36][23].run()  ;
            end
            begin
              drv[36][23].run()  ;
            end
            begin
              mem_check[36][23].run()  ;
            end
            begin
              rf_driver[36][23].run()  ;
            end

            begin
              gen[36][24].run()  ;
            end
            begin
              drv[36][24].run()  ;
            end
            begin
              mem_check[36][24].run()  ;
            end
            begin
              rf_driver[36][24].run()  ;
            end

            begin
              gen[36][25].run()  ;
            end
            begin
              drv[36][25].run()  ;
            end
            begin
              mem_check[36][25].run()  ;
            end
            begin
              rf_driver[36][25].run()  ;
            end

            begin
              gen[36][26].run()  ;
            end
            begin
              drv[36][26].run()  ;
            end
            begin
              mem_check[36][26].run()  ;
            end
            begin
              rf_driver[36][26].run()  ;
            end

            begin
              gen[36][27].run()  ;
            end
            begin
              drv[36][27].run()  ;
            end
            begin
              mem_check[36][27].run()  ;
            end
            begin
              rf_driver[36][27].run()  ;
            end

            begin
              gen[36][28].run()  ;
            end
            begin
              drv[36][28].run()  ;
            end
            begin
              mem_check[36][28].run()  ;
            end
            begin
              rf_driver[36][28].run()  ;
            end

            begin
              gen[36][29].run()  ;
            end
            begin
              drv[36][29].run()  ;
            end
            begin
              mem_check[36][29].run()  ;
            end
            begin
              rf_driver[36][29].run()  ;
            end

            begin
              gen[36][30].run()  ;
            end
            begin
              drv[36][30].run()  ;
            end
            begin
              mem_check[36][30].run()  ;
            end
            begin
              rf_driver[36][30].run()  ;
            end

            begin
              gen[36][31].run()  ;
            end
            begin
              drv[36][31].run()  ;
            end
            begin
              mem_check[36][31].run()  ;
            end
            begin
              rf_driver[36][31].run()  ;
            end

            begin
              ldst_driver[37].run()  ;
            end
            begin
              mgr[37].run()  ;
            end
            begin
              oob_drv[37].run()  ;
            end
            begin
              up_check[37].run()  ;
            end
            begin
              gen[37][0].run()  ;
            end
            begin
              drv[37][0].run()  ;
            end
            begin
              mem_check[37][0].run()  ;
            end
            begin
              rf_driver[37][0].run()  ;
            end

            begin
              gen[37][1].run()  ;
            end
            begin
              drv[37][1].run()  ;
            end
            begin
              mem_check[37][1].run()  ;
            end
            begin
              rf_driver[37][1].run()  ;
            end

            begin
              gen[37][2].run()  ;
            end
            begin
              drv[37][2].run()  ;
            end
            begin
              mem_check[37][2].run()  ;
            end
            begin
              rf_driver[37][2].run()  ;
            end

            begin
              gen[37][3].run()  ;
            end
            begin
              drv[37][3].run()  ;
            end
            begin
              mem_check[37][3].run()  ;
            end
            begin
              rf_driver[37][3].run()  ;
            end

            begin
              gen[37][4].run()  ;
            end
            begin
              drv[37][4].run()  ;
            end
            begin
              mem_check[37][4].run()  ;
            end
            begin
              rf_driver[37][4].run()  ;
            end

            begin
              gen[37][5].run()  ;
            end
            begin
              drv[37][5].run()  ;
            end
            begin
              mem_check[37][5].run()  ;
            end
            begin
              rf_driver[37][5].run()  ;
            end

            begin
              gen[37][6].run()  ;
            end
            begin
              drv[37][6].run()  ;
            end
            begin
              mem_check[37][6].run()  ;
            end
            begin
              rf_driver[37][6].run()  ;
            end

            begin
              gen[37][7].run()  ;
            end
            begin
              drv[37][7].run()  ;
            end
            begin
              mem_check[37][7].run()  ;
            end
            begin
              rf_driver[37][7].run()  ;
            end

            begin
              gen[37][8].run()  ;
            end
            begin
              drv[37][8].run()  ;
            end
            begin
              mem_check[37][8].run()  ;
            end
            begin
              rf_driver[37][8].run()  ;
            end

            begin
              gen[37][9].run()  ;
            end
            begin
              drv[37][9].run()  ;
            end
            begin
              mem_check[37][9].run()  ;
            end
            begin
              rf_driver[37][9].run()  ;
            end

            begin
              gen[37][10].run()  ;
            end
            begin
              drv[37][10].run()  ;
            end
            begin
              mem_check[37][10].run()  ;
            end
            begin
              rf_driver[37][10].run()  ;
            end

            begin
              gen[37][11].run()  ;
            end
            begin
              drv[37][11].run()  ;
            end
            begin
              mem_check[37][11].run()  ;
            end
            begin
              rf_driver[37][11].run()  ;
            end

            begin
              gen[37][12].run()  ;
            end
            begin
              drv[37][12].run()  ;
            end
            begin
              mem_check[37][12].run()  ;
            end
            begin
              rf_driver[37][12].run()  ;
            end

            begin
              gen[37][13].run()  ;
            end
            begin
              drv[37][13].run()  ;
            end
            begin
              mem_check[37][13].run()  ;
            end
            begin
              rf_driver[37][13].run()  ;
            end

            begin
              gen[37][14].run()  ;
            end
            begin
              drv[37][14].run()  ;
            end
            begin
              mem_check[37][14].run()  ;
            end
            begin
              rf_driver[37][14].run()  ;
            end

            begin
              gen[37][15].run()  ;
            end
            begin
              drv[37][15].run()  ;
            end
            begin
              mem_check[37][15].run()  ;
            end
            begin
              rf_driver[37][15].run()  ;
            end

            begin
              gen[37][16].run()  ;
            end
            begin
              drv[37][16].run()  ;
            end
            begin
              mem_check[37][16].run()  ;
            end
            begin
              rf_driver[37][16].run()  ;
            end

            begin
              gen[37][17].run()  ;
            end
            begin
              drv[37][17].run()  ;
            end
            begin
              mem_check[37][17].run()  ;
            end
            begin
              rf_driver[37][17].run()  ;
            end

            begin
              gen[37][18].run()  ;
            end
            begin
              drv[37][18].run()  ;
            end
            begin
              mem_check[37][18].run()  ;
            end
            begin
              rf_driver[37][18].run()  ;
            end

            begin
              gen[37][19].run()  ;
            end
            begin
              drv[37][19].run()  ;
            end
            begin
              mem_check[37][19].run()  ;
            end
            begin
              rf_driver[37][19].run()  ;
            end

            begin
              gen[37][20].run()  ;
            end
            begin
              drv[37][20].run()  ;
            end
            begin
              mem_check[37][20].run()  ;
            end
            begin
              rf_driver[37][20].run()  ;
            end

            begin
              gen[37][21].run()  ;
            end
            begin
              drv[37][21].run()  ;
            end
            begin
              mem_check[37][21].run()  ;
            end
            begin
              rf_driver[37][21].run()  ;
            end

            begin
              gen[37][22].run()  ;
            end
            begin
              drv[37][22].run()  ;
            end
            begin
              mem_check[37][22].run()  ;
            end
            begin
              rf_driver[37][22].run()  ;
            end

            begin
              gen[37][23].run()  ;
            end
            begin
              drv[37][23].run()  ;
            end
            begin
              mem_check[37][23].run()  ;
            end
            begin
              rf_driver[37][23].run()  ;
            end

            begin
              gen[37][24].run()  ;
            end
            begin
              drv[37][24].run()  ;
            end
            begin
              mem_check[37][24].run()  ;
            end
            begin
              rf_driver[37][24].run()  ;
            end

            begin
              gen[37][25].run()  ;
            end
            begin
              drv[37][25].run()  ;
            end
            begin
              mem_check[37][25].run()  ;
            end
            begin
              rf_driver[37][25].run()  ;
            end

            begin
              gen[37][26].run()  ;
            end
            begin
              drv[37][26].run()  ;
            end
            begin
              mem_check[37][26].run()  ;
            end
            begin
              rf_driver[37][26].run()  ;
            end

            begin
              gen[37][27].run()  ;
            end
            begin
              drv[37][27].run()  ;
            end
            begin
              mem_check[37][27].run()  ;
            end
            begin
              rf_driver[37][27].run()  ;
            end

            begin
              gen[37][28].run()  ;
            end
            begin
              drv[37][28].run()  ;
            end
            begin
              mem_check[37][28].run()  ;
            end
            begin
              rf_driver[37][28].run()  ;
            end

            begin
              gen[37][29].run()  ;
            end
            begin
              drv[37][29].run()  ;
            end
            begin
              mem_check[37][29].run()  ;
            end
            begin
              rf_driver[37][29].run()  ;
            end

            begin
              gen[37][30].run()  ;
            end
            begin
              drv[37][30].run()  ;
            end
            begin
              mem_check[37][30].run()  ;
            end
            begin
              rf_driver[37][30].run()  ;
            end

            begin
              gen[37][31].run()  ;
            end
            begin
              drv[37][31].run()  ;
            end
            begin
              mem_check[37][31].run()  ;
            end
            begin
              rf_driver[37][31].run()  ;
            end

            begin
              ldst_driver[38].run()  ;
            end
            begin
              mgr[38].run()  ;
            end
            begin
              oob_drv[38].run()  ;
            end
            begin
              up_check[38].run()  ;
            end
            begin
              gen[38][0].run()  ;
            end
            begin
              drv[38][0].run()  ;
            end
            begin
              mem_check[38][0].run()  ;
            end
            begin
              rf_driver[38][0].run()  ;
            end

            begin
              gen[38][1].run()  ;
            end
            begin
              drv[38][1].run()  ;
            end
            begin
              mem_check[38][1].run()  ;
            end
            begin
              rf_driver[38][1].run()  ;
            end

            begin
              gen[38][2].run()  ;
            end
            begin
              drv[38][2].run()  ;
            end
            begin
              mem_check[38][2].run()  ;
            end
            begin
              rf_driver[38][2].run()  ;
            end

            begin
              gen[38][3].run()  ;
            end
            begin
              drv[38][3].run()  ;
            end
            begin
              mem_check[38][3].run()  ;
            end
            begin
              rf_driver[38][3].run()  ;
            end

            begin
              gen[38][4].run()  ;
            end
            begin
              drv[38][4].run()  ;
            end
            begin
              mem_check[38][4].run()  ;
            end
            begin
              rf_driver[38][4].run()  ;
            end

            begin
              gen[38][5].run()  ;
            end
            begin
              drv[38][5].run()  ;
            end
            begin
              mem_check[38][5].run()  ;
            end
            begin
              rf_driver[38][5].run()  ;
            end

            begin
              gen[38][6].run()  ;
            end
            begin
              drv[38][6].run()  ;
            end
            begin
              mem_check[38][6].run()  ;
            end
            begin
              rf_driver[38][6].run()  ;
            end

            begin
              gen[38][7].run()  ;
            end
            begin
              drv[38][7].run()  ;
            end
            begin
              mem_check[38][7].run()  ;
            end
            begin
              rf_driver[38][7].run()  ;
            end

            begin
              gen[38][8].run()  ;
            end
            begin
              drv[38][8].run()  ;
            end
            begin
              mem_check[38][8].run()  ;
            end
            begin
              rf_driver[38][8].run()  ;
            end

            begin
              gen[38][9].run()  ;
            end
            begin
              drv[38][9].run()  ;
            end
            begin
              mem_check[38][9].run()  ;
            end
            begin
              rf_driver[38][9].run()  ;
            end

            begin
              gen[38][10].run()  ;
            end
            begin
              drv[38][10].run()  ;
            end
            begin
              mem_check[38][10].run()  ;
            end
            begin
              rf_driver[38][10].run()  ;
            end

            begin
              gen[38][11].run()  ;
            end
            begin
              drv[38][11].run()  ;
            end
            begin
              mem_check[38][11].run()  ;
            end
            begin
              rf_driver[38][11].run()  ;
            end

            begin
              gen[38][12].run()  ;
            end
            begin
              drv[38][12].run()  ;
            end
            begin
              mem_check[38][12].run()  ;
            end
            begin
              rf_driver[38][12].run()  ;
            end

            begin
              gen[38][13].run()  ;
            end
            begin
              drv[38][13].run()  ;
            end
            begin
              mem_check[38][13].run()  ;
            end
            begin
              rf_driver[38][13].run()  ;
            end

            begin
              gen[38][14].run()  ;
            end
            begin
              drv[38][14].run()  ;
            end
            begin
              mem_check[38][14].run()  ;
            end
            begin
              rf_driver[38][14].run()  ;
            end

            begin
              gen[38][15].run()  ;
            end
            begin
              drv[38][15].run()  ;
            end
            begin
              mem_check[38][15].run()  ;
            end
            begin
              rf_driver[38][15].run()  ;
            end

            begin
              gen[38][16].run()  ;
            end
            begin
              drv[38][16].run()  ;
            end
            begin
              mem_check[38][16].run()  ;
            end
            begin
              rf_driver[38][16].run()  ;
            end

            begin
              gen[38][17].run()  ;
            end
            begin
              drv[38][17].run()  ;
            end
            begin
              mem_check[38][17].run()  ;
            end
            begin
              rf_driver[38][17].run()  ;
            end

            begin
              gen[38][18].run()  ;
            end
            begin
              drv[38][18].run()  ;
            end
            begin
              mem_check[38][18].run()  ;
            end
            begin
              rf_driver[38][18].run()  ;
            end

            begin
              gen[38][19].run()  ;
            end
            begin
              drv[38][19].run()  ;
            end
            begin
              mem_check[38][19].run()  ;
            end
            begin
              rf_driver[38][19].run()  ;
            end

            begin
              gen[38][20].run()  ;
            end
            begin
              drv[38][20].run()  ;
            end
            begin
              mem_check[38][20].run()  ;
            end
            begin
              rf_driver[38][20].run()  ;
            end

            begin
              gen[38][21].run()  ;
            end
            begin
              drv[38][21].run()  ;
            end
            begin
              mem_check[38][21].run()  ;
            end
            begin
              rf_driver[38][21].run()  ;
            end

            begin
              gen[38][22].run()  ;
            end
            begin
              drv[38][22].run()  ;
            end
            begin
              mem_check[38][22].run()  ;
            end
            begin
              rf_driver[38][22].run()  ;
            end

            begin
              gen[38][23].run()  ;
            end
            begin
              drv[38][23].run()  ;
            end
            begin
              mem_check[38][23].run()  ;
            end
            begin
              rf_driver[38][23].run()  ;
            end

            begin
              gen[38][24].run()  ;
            end
            begin
              drv[38][24].run()  ;
            end
            begin
              mem_check[38][24].run()  ;
            end
            begin
              rf_driver[38][24].run()  ;
            end

            begin
              gen[38][25].run()  ;
            end
            begin
              drv[38][25].run()  ;
            end
            begin
              mem_check[38][25].run()  ;
            end
            begin
              rf_driver[38][25].run()  ;
            end

            begin
              gen[38][26].run()  ;
            end
            begin
              drv[38][26].run()  ;
            end
            begin
              mem_check[38][26].run()  ;
            end
            begin
              rf_driver[38][26].run()  ;
            end

            begin
              gen[38][27].run()  ;
            end
            begin
              drv[38][27].run()  ;
            end
            begin
              mem_check[38][27].run()  ;
            end
            begin
              rf_driver[38][27].run()  ;
            end

            begin
              gen[38][28].run()  ;
            end
            begin
              drv[38][28].run()  ;
            end
            begin
              mem_check[38][28].run()  ;
            end
            begin
              rf_driver[38][28].run()  ;
            end

            begin
              gen[38][29].run()  ;
            end
            begin
              drv[38][29].run()  ;
            end
            begin
              mem_check[38][29].run()  ;
            end
            begin
              rf_driver[38][29].run()  ;
            end

            begin
              gen[38][30].run()  ;
            end
            begin
              drv[38][30].run()  ;
            end
            begin
              mem_check[38][30].run()  ;
            end
            begin
              rf_driver[38][30].run()  ;
            end

            begin
              gen[38][31].run()  ;
            end
            begin
              drv[38][31].run()  ;
            end
            begin
              mem_check[38][31].run()  ;
            end
            begin
              rf_driver[38][31].run()  ;
            end

            begin
              ldst_driver[39].run()  ;
            end
            begin
              mgr[39].run()  ;
            end
            begin
              oob_drv[39].run()  ;
            end
            begin
              up_check[39].run()  ;
            end
            begin
              gen[39][0].run()  ;
            end
            begin
              drv[39][0].run()  ;
            end
            begin
              mem_check[39][0].run()  ;
            end
            begin
              rf_driver[39][0].run()  ;
            end

            begin
              gen[39][1].run()  ;
            end
            begin
              drv[39][1].run()  ;
            end
            begin
              mem_check[39][1].run()  ;
            end
            begin
              rf_driver[39][1].run()  ;
            end

            begin
              gen[39][2].run()  ;
            end
            begin
              drv[39][2].run()  ;
            end
            begin
              mem_check[39][2].run()  ;
            end
            begin
              rf_driver[39][2].run()  ;
            end

            begin
              gen[39][3].run()  ;
            end
            begin
              drv[39][3].run()  ;
            end
            begin
              mem_check[39][3].run()  ;
            end
            begin
              rf_driver[39][3].run()  ;
            end

            begin
              gen[39][4].run()  ;
            end
            begin
              drv[39][4].run()  ;
            end
            begin
              mem_check[39][4].run()  ;
            end
            begin
              rf_driver[39][4].run()  ;
            end

            begin
              gen[39][5].run()  ;
            end
            begin
              drv[39][5].run()  ;
            end
            begin
              mem_check[39][5].run()  ;
            end
            begin
              rf_driver[39][5].run()  ;
            end

            begin
              gen[39][6].run()  ;
            end
            begin
              drv[39][6].run()  ;
            end
            begin
              mem_check[39][6].run()  ;
            end
            begin
              rf_driver[39][6].run()  ;
            end

            begin
              gen[39][7].run()  ;
            end
            begin
              drv[39][7].run()  ;
            end
            begin
              mem_check[39][7].run()  ;
            end
            begin
              rf_driver[39][7].run()  ;
            end

            begin
              gen[39][8].run()  ;
            end
            begin
              drv[39][8].run()  ;
            end
            begin
              mem_check[39][8].run()  ;
            end
            begin
              rf_driver[39][8].run()  ;
            end

            begin
              gen[39][9].run()  ;
            end
            begin
              drv[39][9].run()  ;
            end
            begin
              mem_check[39][9].run()  ;
            end
            begin
              rf_driver[39][9].run()  ;
            end

            begin
              gen[39][10].run()  ;
            end
            begin
              drv[39][10].run()  ;
            end
            begin
              mem_check[39][10].run()  ;
            end
            begin
              rf_driver[39][10].run()  ;
            end

            begin
              gen[39][11].run()  ;
            end
            begin
              drv[39][11].run()  ;
            end
            begin
              mem_check[39][11].run()  ;
            end
            begin
              rf_driver[39][11].run()  ;
            end

            begin
              gen[39][12].run()  ;
            end
            begin
              drv[39][12].run()  ;
            end
            begin
              mem_check[39][12].run()  ;
            end
            begin
              rf_driver[39][12].run()  ;
            end

            begin
              gen[39][13].run()  ;
            end
            begin
              drv[39][13].run()  ;
            end
            begin
              mem_check[39][13].run()  ;
            end
            begin
              rf_driver[39][13].run()  ;
            end

            begin
              gen[39][14].run()  ;
            end
            begin
              drv[39][14].run()  ;
            end
            begin
              mem_check[39][14].run()  ;
            end
            begin
              rf_driver[39][14].run()  ;
            end

            begin
              gen[39][15].run()  ;
            end
            begin
              drv[39][15].run()  ;
            end
            begin
              mem_check[39][15].run()  ;
            end
            begin
              rf_driver[39][15].run()  ;
            end

            begin
              gen[39][16].run()  ;
            end
            begin
              drv[39][16].run()  ;
            end
            begin
              mem_check[39][16].run()  ;
            end
            begin
              rf_driver[39][16].run()  ;
            end

            begin
              gen[39][17].run()  ;
            end
            begin
              drv[39][17].run()  ;
            end
            begin
              mem_check[39][17].run()  ;
            end
            begin
              rf_driver[39][17].run()  ;
            end

            begin
              gen[39][18].run()  ;
            end
            begin
              drv[39][18].run()  ;
            end
            begin
              mem_check[39][18].run()  ;
            end
            begin
              rf_driver[39][18].run()  ;
            end

            begin
              gen[39][19].run()  ;
            end
            begin
              drv[39][19].run()  ;
            end
            begin
              mem_check[39][19].run()  ;
            end
            begin
              rf_driver[39][19].run()  ;
            end

            begin
              gen[39][20].run()  ;
            end
            begin
              drv[39][20].run()  ;
            end
            begin
              mem_check[39][20].run()  ;
            end
            begin
              rf_driver[39][20].run()  ;
            end

            begin
              gen[39][21].run()  ;
            end
            begin
              drv[39][21].run()  ;
            end
            begin
              mem_check[39][21].run()  ;
            end
            begin
              rf_driver[39][21].run()  ;
            end

            begin
              gen[39][22].run()  ;
            end
            begin
              drv[39][22].run()  ;
            end
            begin
              mem_check[39][22].run()  ;
            end
            begin
              rf_driver[39][22].run()  ;
            end

            begin
              gen[39][23].run()  ;
            end
            begin
              drv[39][23].run()  ;
            end
            begin
              mem_check[39][23].run()  ;
            end
            begin
              rf_driver[39][23].run()  ;
            end

            begin
              gen[39][24].run()  ;
            end
            begin
              drv[39][24].run()  ;
            end
            begin
              mem_check[39][24].run()  ;
            end
            begin
              rf_driver[39][24].run()  ;
            end

            begin
              gen[39][25].run()  ;
            end
            begin
              drv[39][25].run()  ;
            end
            begin
              mem_check[39][25].run()  ;
            end
            begin
              rf_driver[39][25].run()  ;
            end

            begin
              gen[39][26].run()  ;
            end
            begin
              drv[39][26].run()  ;
            end
            begin
              mem_check[39][26].run()  ;
            end
            begin
              rf_driver[39][26].run()  ;
            end

            begin
              gen[39][27].run()  ;
            end
            begin
              drv[39][27].run()  ;
            end
            begin
              mem_check[39][27].run()  ;
            end
            begin
              rf_driver[39][27].run()  ;
            end

            begin
              gen[39][28].run()  ;
            end
            begin
              drv[39][28].run()  ;
            end
            begin
              mem_check[39][28].run()  ;
            end
            begin
              rf_driver[39][28].run()  ;
            end

            begin
              gen[39][29].run()  ;
            end
            begin
              drv[39][29].run()  ;
            end
            begin
              mem_check[39][29].run()  ;
            end
            begin
              rf_driver[39][29].run()  ;
            end

            begin
              gen[39][30].run()  ;
            end
            begin
              drv[39][30].run()  ;
            end
            begin
              mem_check[39][30].run()  ;
            end
            begin
              rf_driver[39][30].run()  ;
            end

            begin
              gen[39][31].run()  ;
            end
            begin
              drv[39][31].run()  ;
            end
            begin
              mem_check[39][31].run()  ;
            end
            begin
              rf_driver[39][31].run()  ;
            end

            begin
              ldst_driver[40].run()  ;
            end
            begin
              mgr[40].run()  ;
            end
            begin
              oob_drv[40].run()  ;
            end
            begin
              up_check[40].run()  ;
            end
            begin
              gen[40][0].run()  ;
            end
            begin
              drv[40][0].run()  ;
            end
            begin
              mem_check[40][0].run()  ;
            end
            begin
              rf_driver[40][0].run()  ;
            end

            begin
              gen[40][1].run()  ;
            end
            begin
              drv[40][1].run()  ;
            end
            begin
              mem_check[40][1].run()  ;
            end
            begin
              rf_driver[40][1].run()  ;
            end

            begin
              gen[40][2].run()  ;
            end
            begin
              drv[40][2].run()  ;
            end
            begin
              mem_check[40][2].run()  ;
            end
            begin
              rf_driver[40][2].run()  ;
            end

            begin
              gen[40][3].run()  ;
            end
            begin
              drv[40][3].run()  ;
            end
            begin
              mem_check[40][3].run()  ;
            end
            begin
              rf_driver[40][3].run()  ;
            end

            begin
              gen[40][4].run()  ;
            end
            begin
              drv[40][4].run()  ;
            end
            begin
              mem_check[40][4].run()  ;
            end
            begin
              rf_driver[40][4].run()  ;
            end

            begin
              gen[40][5].run()  ;
            end
            begin
              drv[40][5].run()  ;
            end
            begin
              mem_check[40][5].run()  ;
            end
            begin
              rf_driver[40][5].run()  ;
            end

            begin
              gen[40][6].run()  ;
            end
            begin
              drv[40][6].run()  ;
            end
            begin
              mem_check[40][6].run()  ;
            end
            begin
              rf_driver[40][6].run()  ;
            end

            begin
              gen[40][7].run()  ;
            end
            begin
              drv[40][7].run()  ;
            end
            begin
              mem_check[40][7].run()  ;
            end
            begin
              rf_driver[40][7].run()  ;
            end

            begin
              gen[40][8].run()  ;
            end
            begin
              drv[40][8].run()  ;
            end
            begin
              mem_check[40][8].run()  ;
            end
            begin
              rf_driver[40][8].run()  ;
            end

            begin
              gen[40][9].run()  ;
            end
            begin
              drv[40][9].run()  ;
            end
            begin
              mem_check[40][9].run()  ;
            end
            begin
              rf_driver[40][9].run()  ;
            end

            begin
              gen[40][10].run()  ;
            end
            begin
              drv[40][10].run()  ;
            end
            begin
              mem_check[40][10].run()  ;
            end
            begin
              rf_driver[40][10].run()  ;
            end

            begin
              gen[40][11].run()  ;
            end
            begin
              drv[40][11].run()  ;
            end
            begin
              mem_check[40][11].run()  ;
            end
            begin
              rf_driver[40][11].run()  ;
            end

            begin
              gen[40][12].run()  ;
            end
            begin
              drv[40][12].run()  ;
            end
            begin
              mem_check[40][12].run()  ;
            end
            begin
              rf_driver[40][12].run()  ;
            end

            begin
              gen[40][13].run()  ;
            end
            begin
              drv[40][13].run()  ;
            end
            begin
              mem_check[40][13].run()  ;
            end
            begin
              rf_driver[40][13].run()  ;
            end

            begin
              gen[40][14].run()  ;
            end
            begin
              drv[40][14].run()  ;
            end
            begin
              mem_check[40][14].run()  ;
            end
            begin
              rf_driver[40][14].run()  ;
            end

            begin
              gen[40][15].run()  ;
            end
            begin
              drv[40][15].run()  ;
            end
            begin
              mem_check[40][15].run()  ;
            end
            begin
              rf_driver[40][15].run()  ;
            end

            begin
              gen[40][16].run()  ;
            end
            begin
              drv[40][16].run()  ;
            end
            begin
              mem_check[40][16].run()  ;
            end
            begin
              rf_driver[40][16].run()  ;
            end

            begin
              gen[40][17].run()  ;
            end
            begin
              drv[40][17].run()  ;
            end
            begin
              mem_check[40][17].run()  ;
            end
            begin
              rf_driver[40][17].run()  ;
            end

            begin
              gen[40][18].run()  ;
            end
            begin
              drv[40][18].run()  ;
            end
            begin
              mem_check[40][18].run()  ;
            end
            begin
              rf_driver[40][18].run()  ;
            end

            begin
              gen[40][19].run()  ;
            end
            begin
              drv[40][19].run()  ;
            end
            begin
              mem_check[40][19].run()  ;
            end
            begin
              rf_driver[40][19].run()  ;
            end

            begin
              gen[40][20].run()  ;
            end
            begin
              drv[40][20].run()  ;
            end
            begin
              mem_check[40][20].run()  ;
            end
            begin
              rf_driver[40][20].run()  ;
            end

            begin
              gen[40][21].run()  ;
            end
            begin
              drv[40][21].run()  ;
            end
            begin
              mem_check[40][21].run()  ;
            end
            begin
              rf_driver[40][21].run()  ;
            end

            begin
              gen[40][22].run()  ;
            end
            begin
              drv[40][22].run()  ;
            end
            begin
              mem_check[40][22].run()  ;
            end
            begin
              rf_driver[40][22].run()  ;
            end

            begin
              gen[40][23].run()  ;
            end
            begin
              drv[40][23].run()  ;
            end
            begin
              mem_check[40][23].run()  ;
            end
            begin
              rf_driver[40][23].run()  ;
            end

            begin
              gen[40][24].run()  ;
            end
            begin
              drv[40][24].run()  ;
            end
            begin
              mem_check[40][24].run()  ;
            end
            begin
              rf_driver[40][24].run()  ;
            end

            begin
              gen[40][25].run()  ;
            end
            begin
              drv[40][25].run()  ;
            end
            begin
              mem_check[40][25].run()  ;
            end
            begin
              rf_driver[40][25].run()  ;
            end

            begin
              gen[40][26].run()  ;
            end
            begin
              drv[40][26].run()  ;
            end
            begin
              mem_check[40][26].run()  ;
            end
            begin
              rf_driver[40][26].run()  ;
            end

            begin
              gen[40][27].run()  ;
            end
            begin
              drv[40][27].run()  ;
            end
            begin
              mem_check[40][27].run()  ;
            end
            begin
              rf_driver[40][27].run()  ;
            end

            begin
              gen[40][28].run()  ;
            end
            begin
              drv[40][28].run()  ;
            end
            begin
              mem_check[40][28].run()  ;
            end
            begin
              rf_driver[40][28].run()  ;
            end

            begin
              gen[40][29].run()  ;
            end
            begin
              drv[40][29].run()  ;
            end
            begin
              mem_check[40][29].run()  ;
            end
            begin
              rf_driver[40][29].run()  ;
            end

            begin
              gen[40][30].run()  ;
            end
            begin
              drv[40][30].run()  ;
            end
            begin
              mem_check[40][30].run()  ;
            end
            begin
              rf_driver[40][30].run()  ;
            end

            begin
              gen[40][31].run()  ;
            end
            begin
              drv[40][31].run()  ;
            end
            begin
              mem_check[40][31].run()  ;
            end
            begin
              rf_driver[40][31].run()  ;
            end

            begin
              ldst_driver[41].run()  ;
            end
            begin
              mgr[41].run()  ;
            end
            begin
              oob_drv[41].run()  ;
            end
            begin
              up_check[41].run()  ;
            end
            begin
              gen[41][0].run()  ;
            end
            begin
              drv[41][0].run()  ;
            end
            begin
              mem_check[41][0].run()  ;
            end
            begin
              rf_driver[41][0].run()  ;
            end

            begin
              gen[41][1].run()  ;
            end
            begin
              drv[41][1].run()  ;
            end
            begin
              mem_check[41][1].run()  ;
            end
            begin
              rf_driver[41][1].run()  ;
            end

            begin
              gen[41][2].run()  ;
            end
            begin
              drv[41][2].run()  ;
            end
            begin
              mem_check[41][2].run()  ;
            end
            begin
              rf_driver[41][2].run()  ;
            end

            begin
              gen[41][3].run()  ;
            end
            begin
              drv[41][3].run()  ;
            end
            begin
              mem_check[41][3].run()  ;
            end
            begin
              rf_driver[41][3].run()  ;
            end

            begin
              gen[41][4].run()  ;
            end
            begin
              drv[41][4].run()  ;
            end
            begin
              mem_check[41][4].run()  ;
            end
            begin
              rf_driver[41][4].run()  ;
            end

            begin
              gen[41][5].run()  ;
            end
            begin
              drv[41][5].run()  ;
            end
            begin
              mem_check[41][5].run()  ;
            end
            begin
              rf_driver[41][5].run()  ;
            end

            begin
              gen[41][6].run()  ;
            end
            begin
              drv[41][6].run()  ;
            end
            begin
              mem_check[41][6].run()  ;
            end
            begin
              rf_driver[41][6].run()  ;
            end

            begin
              gen[41][7].run()  ;
            end
            begin
              drv[41][7].run()  ;
            end
            begin
              mem_check[41][7].run()  ;
            end
            begin
              rf_driver[41][7].run()  ;
            end

            begin
              gen[41][8].run()  ;
            end
            begin
              drv[41][8].run()  ;
            end
            begin
              mem_check[41][8].run()  ;
            end
            begin
              rf_driver[41][8].run()  ;
            end

            begin
              gen[41][9].run()  ;
            end
            begin
              drv[41][9].run()  ;
            end
            begin
              mem_check[41][9].run()  ;
            end
            begin
              rf_driver[41][9].run()  ;
            end

            begin
              gen[41][10].run()  ;
            end
            begin
              drv[41][10].run()  ;
            end
            begin
              mem_check[41][10].run()  ;
            end
            begin
              rf_driver[41][10].run()  ;
            end

            begin
              gen[41][11].run()  ;
            end
            begin
              drv[41][11].run()  ;
            end
            begin
              mem_check[41][11].run()  ;
            end
            begin
              rf_driver[41][11].run()  ;
            end

            begin
              gen[41][12].run()  ;
            end
            begin
              drv[41][12].run()  ;
            end
            begin
              mem_check[41][12].run()  ;
            end
            begin
              rf_driver[41][12].run()  ;
            end

            begin
              gen[41][13].run()  ;
            end
            begin
              drv[41][13].run()  ;
            end
            begin
              mem_check[41][13].run()  ;
            end
            begin
              rf_driver[41][13].run()  ;
            end

            begin
              gen[41][14].run()  ;
            end
            begin
              drv[41][14].run()  ;
            end
            begin
              mem_check[41][14].run()  ;
            end
            begin
              rf_driver[41][14].run()  ;
            end

            begin
              gen[41][15].run()  ;
            end
            begin
              drv[41][15].run()  ;
            end
            begin
              mem_check[41][15].run()  ;
            end
            begin
              rf_driver[41][15].run()  ;
            end

            begin
              gen[41][16].run()  ;
            end
            begin
              drv[41][16].run()  ;
            end
            begin
              mem_check[41][16].run()  ;
            end
            begin
              rf_driver[41][16].run()  ;
            end

            begin
              gen[41][17].run()  ;
            end
            begin
              drv[41][17].run()  ;
            end
            begin
              mem_check[41][17].run()  ;
            end
            begin
              rf_driver[41][17].run()  ;
            end

            begin
              gen[41][18].run()  ;
            end
            begin
              drv[41][18].run()  ;
            end
            begin
              mem_check[41][18].run()  ;
            end
            begin
              rf_driver[41][18].run()  ;
            end

            begin
              gen[41][19].run()  ;
            end
            begin
              drv[41][19].run()  ;
            end
            begin
              mem_check[41][19].run()  ;
            end
            begin
              rf_driver[41][19].run()  ;
            end

            begin
              gen[41][20].run()  ;
            end
            begin
              drv[41][20].run()  ;
            end
            begin
              mem_check[41][20].run()  ;
            end
            begin
              rf_driver[41][20].run()  ;
            end

            begin
              gen[41][21].run()  ;
            end
            begin
              drv[41][21].run()  ;
            end
            begin
              mem_check[41][21].run()  ;
            end
            begin
              rf_driver[41][21].run()  ;
            end

            begin
              gen[41][22].run()  ;
            end
            begin
              drv[41][22].run()  ;
            end
            begin
              mem_check[41][22].run()  ;
            end
            begin
              rf_driver[41][22].run()  ;
            end

            begin
              gen[41][23].run()  ;
            end
            begin
              drv[41][23].run()  ;
            end
            begin
              mem_check[41][23].run()  ;
            end
            begin
              rf_driver[41][23].run()  ;
            end

            begin
              gen[41][24].run()  ;
            end
            begin
              drv[41][24].run()  ;
            end
            begin
              mem_check[41][24].run()  ;
            end
            begin
              rf_driver[41][24].run()  ;
            end

            begin
              gen[41][25].run()  ;
            end
            begin
              drv[41][25].run()  ;
            end
            begin
              mem_check[41][25].run()  ;
            end
            begin
              rf_driver[41][25].run()  ;
            end

            begin
              gen[41][26].run()  ;
            end
            begin
              drv[41][26].run()  ;
            end
            begin
              mem_check[41][26].run()  ;
            end
            begin
              rf_driver[41][26].run()  ;
            end

            begin
              gen[41][27].run()  ;
            end
            begin
              drv[41][27].run()  ;
            end
            begin
              mem_check[41][27].run()  ;
            end
            begin
              rf_driver[41][27].run()  ;
            end

            begin
              gen[41][28].run()  ;
            end
            begin
              drv[41][28].run()  ;
            end
            begin
              mem_check[41][28].run()  ;
            end
            begin
              rf_driver[41][28].run()  ;
            end

            begin
              gen[41][29].run()  ;
            end
            begin
              drv[41][29].run()  ;
            end
            begin
              mem_check[41][29].run()  ;
            end
            begin
              rf_driver[41][29].run()  ;
            end

            begin
              gen[41][30].run()  ;
            end
            begin
              drv[41][30].run()  ;
            end
            begin
              mem_check[41][30].run()  ;
            end
            begin
              rf_driver[41][30].run()  ;
            end

            begin
              gen[41][31].run()  ;
            end
            begin
              drv[41][31].run()  ;
            end
            begin
              mem_check[41][31].run()  ;
            end
            begin
              rf_driver[41][31].run()  ;
            end

            begin
              ldst_driver[42].run()  ;
            end
            begin
              mgr[42].run()  ;
            end
            begin
              oob_drv[42].run()  ;
            end
            begin
              up_check[42].run()  ;
            end
            begin
              gen[42][0].run()  ;
            end
            begin
              drv[42][0].run()  ;
            end
            begin
              mem_check[42][0].run()  ;
            end
            begin
              rf_driver[42][0].run()  ;
            end

            begin
              gen[42][1].run()  ;
            end
            begin
              drv[42][1].run()  ;
            end
            begin
              mem_check[42][1].run()  ;
            end
            begin
              rf_driver[42][1].run()  ;
            end

            begin
              gen[42][2].run()  ;
            end
            begin
              drv[42][2].run()  ;
            end
            begin
              mem_check[42][2].run()  ;
            end
            begin
              rf_driver[42][2].run()  ;
            end

            begin
              gen[42][3].run()  ;
            end
            begin
              drv[42][3].run()  ;
            end
            begin
              mem_check[42][3].run()  ;
            end
            begin
              rf_driver[42][3].run()  ;
            end

            begin
              gen[42][4].run()  ;
            end
            begin
              drv[42][4].run()  ;
            end
            begin
              mem_check[42][4].run()  ;
            end
            begin
              rf_driver[42][4].run()  ;
            end

            begin
              gen[42][5].run()  ;
            end
            begin
              drv[42][5].run()  ;
            end
            begin
              mem_check[42][5].run()  ;
            end
            begin
              rf_driver[42][5].run()  ;
            end

            begin
              gen[42][6].run()  ;
            end
            begin
              drv[42][6].run()  ;
            end
            begin
              mem_check[42][6].run()  ;
            end
            begin
              rf_driver[42][6].run()  ;
            end

            begin
              gen[42][7].run()  ;
            end
            begin
              drv[42][7].run()  ;
            end
            begin
              mem_check[42][7].run()  ;
            end
            begin
              rf_driver[42][7].run()  ;
            end

            begin
              gen[42][8].run()  ;
            end
            begin
              drv[42][8].run()  ;
            end
            begin
              mem_check[42][8].run()  ;
            end
            begin
              rf_driver[42][8].run()  ;
            end

            begin
              gen[42][9].run()  ;
            end
            begin
              drv[42][9].run()  ;
            end
            begin
              mem_check[42][9].run()  ;
            end
            begin
              rf_driver[42][9].run()  ;
            end

            begin
              gen[42][10].run()  ;
            end
            begin
              drv[42][10].run()  ;
            end
            begin
              mem_check[42][10].run()  ;
            end
            begin
              rf_driver[42][10].run()  ;
            end

            begin
              gen[42][11].run()  ;
            end
            begin
              drv[42][11].run()  ;
            end
            begin
              mem_check[42][11].run()  ;
            end
            begin
              rf_driver[42][11].run()  ;
            end

            begin
              gen[42][12].run()  ;
            end
            begin
              drv[42][12].run()  ;
            end
            begin
              mem_check[42][12].run()  ;
            end
            begin
              rf_driver[42][12].run()  ;
            end

            begin
              gen[42][13].run()  ;
            end
            begin
              drv[42][13].run()  ;
            end
            begin
              mem_check[42][13].run()  ;
            end
            begin
              rf_driver[42][13].run()  ;
            end

            begin
              gen[42][14].run()  ;
            end
            begin
              drv[42][14].run()  ;
            end
            begin
              mem_check[42][14].run()  ;
            end
            begin
              rf_driver[42][14].run()  ;
            end

            begin
              gen[42][15].run()  ;
            end
            begin
              drv[42][15].run()  ;
            end
            begin
              mem_check[42][15].run()  ;
            end
            begin
              rf_driver[42][15].run()  ;
            end

            begin
              gen[42][16].run()  ;
            end
            begin
              drv[42][16].run()  ;
            end
            begin
              mem_check[42][16].run()  ;
            end
            begin
              rf_driver[42][16].run()  ;
            end

            begin
              gen[42][17].run()  ;
            end
            begin
              drv[42][17].run()  ;
            end
            begin
              mem_check[42][17].run()  ;
            end
            begin
              rf_driver[42][17].run()  ;
            end

            begin
              gen[42][18].run()  ;
            end
            begin
              drv[42][18].run()  ;
            end
            begin
              mem_check[42][18].run()  ;
            end
            begin
              rf_driver[42][18].run()  ;
            end

            begin
              gen[42][19].run()  ;
            end
            begin
              drv[42][19].run()  ;
            end
            begin
              mem_check[42][19].run()  ;
            end
            begin
              rf_driver[42][19].run()  ;
            end

            begin
              gen[42][20].run()  ;
            end
            begin
              drv[42][20].run()  ;
            end
            begin
              mem_check[42][20].run()  ;
            end
            begin
              rf_driver[42][20].run()  ;
            end

            begin
              gen[42][21].run()  ;
            end
            begin
              drv[42][21].run()  ;
            end
            begin
              mem_check[42][21].run()  ;
            end
            begin
              rf_driver[42][21].run()  ;
            end

            begin
              gen[42][22].run()  ;
            end
            begin
              drv[42][22].run()  ;
            end
            begin
              mem_check[42][22].run()  ;
            end
            begin
              rf_driver[42][22].run()  ;
            end

            begin
              gen[42][23].run()  ;
            end
            begin
              drv[42][23].run()  ;
            end
            begin
              mem_check[42][23].run()  ;
            end
            begin
              rf_driver[42][23].run()  ;
            end

            begin
              gen[42][24].run()  ;
            end
            begin
              drv[42][24].run()  ;
            end
            begin
              mem_check[42][24].run()  ;
            end
            begin
              rf_driver[42][24].run()  ;
            end

            begin
              gen[42][25].run()  ;
            end
            begin
              drv[42][25].run()  ;
            end
            begin
              mem_check[42][25].run()  ;
            end
            begin
              rf_driver[42][25].run()  ;
            end

            begin
              gen[42][26].run()  ;
            end
            begin
              drv[42][26].run()  ;
            end
            begin
              mem_check[42][26].run()  ;
            end
            begin
              rf_driver[42][26].run()  ;
            end

            begin
              gen[42][27].run()  ;
            end
            begin
              drv[42][27].run()  ;
            end
            begin
              mem_check[42][27].run()  ;
            end
            begin
              rf_driver[42][27].run()  ;
            end

            begin
              gen[42][28].run()  ;
            end
            begin
              drv[42][28].run()  ;
            end
            begin
              mem_check[42][28].run()  ;
            end
            begin
              rf_driver[42][28].run()  ;
            end

            begin
              gen[42][29].run()  ;
            end
            begin
              drv[42][29].run()  ;
            end
            begin
              mem_check[42][29].run()  ;
            end
            begin
              rf_driver[42][29].run()  ;
            end

            begin
              gen[42][30].run()  ;
            end
            begin
              drv[42][30].run()  ;
            end
            begin
              mem_check[42][30].run()  ;
            end
            begin
              rf_driver[42][30].run()  ;
            end

            begin
              gen[42][31].run()  ;
            end
            begin
              drv[42][31].run()  ;
            end
            begin
              mem_check[42][31].run()  ;
            end
            begin
              rf_driver[42][31].run()  ;
            end

            begin
              ldst_driver[43].run()  ;
            end
            begin
              mgr[43].run()  ;
            end
            begin
              oob_drv[43].run()  ;
            end
            begin
              up_check[43].run()  ;
            end
            begin
              gen[43][0].run()  ;
            end
            begin
              drv[43][0].run()  ;
            end
            begin
              mem_check[43][0].run()  ;
            end
            begin
              rf_driver[43][0].run()  ;
            end

            begin
              gen[43][1].run()  ;
            end
            begin
              drv[43][1].run()  ;
            end
            begin
              mem_check[43][1].run()  ;
            end
            begin
              rf_driver[43][1].run()  ;
            end

            begin
              gen[43][2].run()  ;
            end
            begin
              drv[43][2].run()  ;
            end
            begin
              mem_check[43][2].run()  ;
            end
            begin
              rf_driver[43][2].run()  ;
            end

            begin
              gen[43][3].run()  ;
            end
            begin
              drv[43][3].run()  ;
            end
            begin
              mem_check[43][3].run()  ;
            end
            begin
              rf_driver[43][3].run()  ;
            end

            begin
              gen[43][4].run()  ;
            end
            begin
              drv[43][4].run()  ;
            end
            begin
              mem_check[43][4].run()  ;
            end
            begin
              rf_driver[43][4].run()  ;
            end

            begin
              gen[43][5].run()  ;
            end
            begin
              drv[43][5].run()  ;
            end
            begin
              mem_check[43][5].run()  ;
            end
            begin
              rf_driver[43][5].run()  ;
            end

            begin
              gen[43][6].run()  ;
            end
            begin
              drv[43][6].run()  ;
            end
            begin
              mem_check[43][6].run()  ;
            end
            begin
              rf_driver[43][6].run()  ;
            end

            begin
              gen[43][7].run()  ;
            end
            begin
              drv[43][7].run()  ;
            end
            begin
              mem_check[43][7].run()  ;
            end
            begin
              rf_driver[43][7].run()  ;
            end

            begin
              gen[43][8].run()  ;
            end
            begin
              drv[43][8].run()  ;
            end
            begin
              mem_check[43][8].run()  ;
            end
            begin
              rf_driver[43][8].run()  ;
            end

            begin
              gen[43][9].run()  ;
            end
            begin
              drv[43][9].run()  ;
            end
            begin
              mem_check[43][9].run()  ;
            end
            begin
              rf_driver[43][9].run()  ;
            end

            begin
              gen[43][10].run()  ;
            end
            begin
              drv[43][10].run()  ;
            end
            begin
              mem_check[43][10].run()  ;
            end
            begin
              rf_driver[43][10].run()  ;
            end

            begin
              gen[43][11].run()  ;
            end
            begin
              drv[43][11].run()  ;
            end
            begin
              mem_check[43][11].run()  ;
            end
            begin
              rf_driver[43][11].run()  ;
            end

            begin
              gen[43][12].run()  ;
            end
            begin
              drv[43][12].run()  ;
            end
            begin
              mem_check[43][12].run()  ;
            end
            begin
              rf_driver[43][12].run()  ;
            end

            begin
              gen[43][13].run()  ;
            end
            begin
              drv[43][13].run()  ;
            end
            begin
              mem_check[43][13].run()  ;
            end
            begin
              rf_driver[43][13].run()  ;
            end

            begin
              gen[43][14].run()  ;
            end
            begin
              drv[43][14].run()  ;
            end
            begin
              mem_check[43][14].run()  ;
            end
            begin
              rf_driver[43][14].run()  ;
            end

            begin
              gen[43][15].run()  ;
            end
            begin
              drv[43][15].run()  ;
            end
            begin
              mem_check[43][15].run()  ;
            end
            begin
              rf_driver[43][15].run()  ;
            end

            begin
              gen[43][16].run()  ;
            end
            begin
              drv[43][16].run()  ;
            end
            begin
              mem_check[43][16].run()  ;
            end
            begin
              rf_driver[43][16].run()  ;
            end

            begin
              gen[43][17].run()  ;
            end
            begin
              drv[43][17].run()  ;
            end
            begin
              mem_check[43][17].run()  ;
            end
            begin
              rf_driver[43][17].run()  ;
            end

            begin
              gen[43][18].run()  ;
            end
            begin
              drv[43][18].run()  ;
            end
            begin
              mem_check[43][18].run()  ;
            end
            begin
              rf_driver[43][18].run()  ;
            end

            begin
              gen[43][19].run()  ;
            end
            begin
              drv[43][19].run()  ;
            end
            begin
              mem_check[43][19].run()  ;
            end
            begin
              rf_driver[43][19].run()  ;
            end

            begin
              gen[43][20].run()  ;
            end
            begin
              drv[43][20].run()  ;
            end
            begin
              mem_check[43][20].run()  ;
            end
            begin
              rf_driver[43][20].run()  ;
            end

            begin
              gen[43][21].run()  ;
            end
            begin
              drv[43][21].run()  ;
            end
            begin
              mem_check[43][21].run()  ;
            end
            begin
              rf_driver[43][21].run()  ;
            end

            begin
              gen[43][22].run()  ;
            end
            begin
              drv[43][22].run()  ;
            end
            begin
              mem_check[43][22].run()  ;
            end
            begin
              rf_driver[43][22].run()  ;
            end

            begin
              gen[43][23].run()  ;
            end
            begin
              drv[43][23].run()  ;
            end
            begin
              mem_check[43][23].run()  ;
            end
            begin
              rf_driver[43][23].run()  ;
            end

            begin
              gen[43][24].run()  ;
            end
            begin
              drv[43][24].run()  ;
            end
            begin
              mem_check[43][24].run()  ;
            end
            begin
              rf_driver[43][24].run()  ;
            end

            begin
              gen[43][25].run()  ;
            end
            begin
              drv[43][25].run()  ;
            end
            begin
              mem_check[43][25].run()  ;
            end
            begin
              rf_driver[43][25].run()  ;
            end

            begin
              gen[43][26].run()  ;
            end
            begin
              drv[43][26].run()  ;
            end
            begin
              mem_check[43][26].run()  ;
            end
            begin
              rf_driver[43][26].run()  ;
            end

            begin
              gen[43][27].run()  ;
            end
            begin
              drv[43][27].run()  ;
            end
            begin
              mem_check[43][27].run()  ;
            end
            begin
              rf_driver[43][27].run()  ;
            end

            begin
              gen[43][28].run()  ;
            end
            begin
              drv[43][28].run()  ;
            end
            begin
              mem_check[43][28].run()  ;
            end
            begin
              rf_driver[43][28].run()  ;
            end

            begin
              gen[43][29].run()  ;
            end
            begin
              drv[43][29].run()  ;
            end
            begin
              mem_check[43][29].run()  ;
            end
            begin
              rf_driver[43][29].run()  ;
            end

            begin
              gen[43][30].run()  ;
            end
            begin
              drv[43][30].run()  ;
            end
            begin
              mem_check[43][30].run()  ;
            end
            begin
              rf_driver[43][30].run()  ;
            end

            begin
              gen[43][31].run()  ;
            end
            begin
              drv[43][31].run()  ;
            end
            begin
              mem_check[43][31].run()  ;
            end
            begin
              rf_driver[43][31].run()  ;
            end

            begin
              ldst_driver[44].run()  ;
            end
            begin
              mgr[44].run()  ;
            end
            begin
              oob_drv[44].run()  ;
            end
            begin
              up_check[44].run()  ;
            end
            begin
              gen[44][0].run()  ;
            end
            begin
              drv[44][0].run()  ;
            end
            begin
              mem_check[44][0].run()  ;
            end
            begin
              rf_driver[44][0].run()  ;
            end

            begin
              gen[44][1].run()  ;
            end
            begin
              drv[44][1].run()  ;
            end
            begin
              mem_check[44][1].run()  ;
            end
            begin
              rf_driver[44][1].run()  ;
            end

            begin
              gen[44][2].run()  ;
            end
            begin
              drv[44][2].run()  ;
            end
            begin
              mem_check[44][2].run()  ;
            end
            begin
              rf_driver[44][2].run()  ;
            end

            begin
              gen[44][3].run()  ;
            end
            begin
              drv[44][3].run()  ;
            end
            begin
              mem_check[44][3].run()  ;
            end
            begin
              rf_driver[44][3].run()  ;
            end

            begin
              gen[44][4].run()  ;
            end
            begin
              drv[44][4].run()  ;
            end
            begin
              mem_check[44][4].run()  ;
            end
            begin
              rf_driver[44][4].run()  ;
            end

            begin
              gen[44][5].run()  ;
            end
            begin
              drv[44][5].run()  ;
            end
            begin
              mem_check[44][5].run()  ;
            end
            begin
              rf_driver[44][5].run()  ;
            end

            begin
              gen[44][6].run()  ;
            end
            begin
              drv[44][6].run()  ;
            end
            begin
              mem_check[44][6].run()  ;
            end
            begin
              rf_driver[44][6].run()  ;
            end

            begin
              gen[44][7].run()  ;
            end
            begin
              drv[44][7].run()  ;
            end
            begin
              mem_check[44][7].run()  ;
            end
            begin
              rf_driver[44][7].run()  ;
            end

            begin
              gen[44][8].run()  ;
            end
            begin
              drv[44][8].run()  ;
            end
            begin
              mem_check[44][8].run()  ;
            end
            begin
              rf_driver[44][8].run()  ;
            end

            begin
              gen[44][9].run()  ;
            end
            begin
              drv[44][9].run()  ;
            end
            begin
              mem_check[44][9].run()  ;
            end
            begin
              rf_driver[44][9].run()  ;
            end

            begin
              gen[44][10].run()  ;
            end
            begin
              drv[44][10].run()  ;
            end
            begin
              mem_check[44][10].run()  ;
            end
            begin
              rf_driver[44][10].run()  ;
            end

            begin
              gen[44][11].run()  ;
            end
            begin
              drv[44][11].run()  ;
            end
            begin
              mem_check[44][11].run()  ;
            end
            begin
              rf_driver[44][11].run()  ;
            end

            begin
              gen[44][12].run()  ;
            end
            begin
              drv[44][12].run()  ;
            end
            begin
              mem_check[44][12].run()  ;
            end
            begin
              rf_driver[44][12].run()  ;
            end

            begin
              gen[44][13].run()  ;
            end
            begin
              drv[44][13].run()  ;
            end
            begin
              mem_check[44][13].run()  ;
            end
            begin
              rf_driver[44][13].run()  ;
            end

            begin
              gen[44][14].run()  ;
            end
            begin
              drv[44][14].run()  ;
            end
            begin
              mem_check[44][14].run()  ;
            end
            begin
              rf_driver[44][14].run()  ;
            end

            begin
              gen[44][15].run()  ;
            end
            begin
              drv[44][15].run()  ;
            end
            begin
              mem_check[44][15].run()  ;
            end
            begin
              rf_driver[44][15].run()  ;
            end

            begin
              gen[44][16].run()  ;
            end
            begin
              drv[44][16].run()  ;
            end
            begin
              mem_check[44][16].run()  ;
            end
            begin
              rf_driver[44][16].run()  ;
            end

            begin
              gen[44][17].run()  ;
            end
            begin
              drv[44][17].run()  ;
            end
            begin
              mem_check[44][17].run()  ;
            end
            begin
              rf_driver[44][17].run()  ;
            end

            begin
              gen[44][18].run()  ;
            end
            begin
              drv[44][18].run()  ;
            end
            begin
              mem_check[44][18].run()  ;
            end
            begin
              rf_driver[44][18].run()  ;
            end

            begin
              gen[44][19].run()  ;
            end
            begin
              drv[44][19].run()  ;
            end
            begin
              mem_check[44][19].run()  ;
            end
            begin
              rf_driver[44][19].run()  ;
            end

            begin
              gen[44][20].run()  ;
            end
            begin
              drv[44][20].run()  ;
            end
            begin
              mem_check[44][20].run()  ;
            end
            begin
              rf_driver[44][20].run()  ;
            end

            begin
              gen[44][21].run()  ;
            end
            begin
              drv[44][21].run()  ;
            end
            begin
              mem_check[44][21].run()  ;
            end
            begin
              rf_driver[44][21].run()  ;
            end

            begin
              gen[44][22].run()  ;
            end
            begin
              drv[44][22].run()  ;
            end
            begin
              mem_check[44][22].run()  ;
            end
            begin
              rf_driver[44][22].run()  ;
            end

            begin
              gen[44][23].run()  ;
            end
            begin
              drv[44][23].run()  ;
            end
            begin
              mem_check[44][23].run()  ;
            end
            begin
              rf_driver[44][23].run()  ;
            end

            begin
              gen[44][24].run()  ;
            end
            begin
              drv[44][24].run()  ;
            end
            begin
              mem_check[44][24].run()  ;
            end
            begin
              rf_driver[44][24].run()  ;
            end

            begin
              gen[44][25].run()  ;
            end
            begin
              drv[44][25].run()  ;
            end
            begin
              mem_check[44][25].run()  ;
            end
            begin
              rf_driver[44][25].run()  ;
            end

            begin
              gen[44][26].run()  ;
            end
            begin
              drv[44][26].run()  ;
            end
            begin
              mem_check[44][26].run()  ;
            end
            begin
              rf_driver[44][26].run()  ;
            end

            begin
              gen[44][27].run()  ;
            end
            begin
              drv[44][27].run()  ;
            end
            begin
              mem_check[44][27].run()  ;
            end
            begin
              rf_driver[44][27].run()  ;
            end

            begin
              gen[44][28].run()  ;
            end
            begin
              drv[44][28].run()  ;
            end
            begin
              mem_check[44][28].run()  ;
            end
            begin
              rf_driver[44][28].run()  ;
            end

            begin
              gen[44][29].run()  ;
            end
            begin
              drv[44][29].run()  ;
            end
            begin
              mem_check[44][29].run()  ;
            end
            begin
              rf_driver[44][29].run()  ;
            end

            begin
              gen[44][30].run()  ;
            end
            begin
              drv[44][30].run()  ;
            end
            begin
              mem_check[44][30].run()  ;
            end
            begin
              rf_driver[44][30].run()  ;
            end

            begin
              gen[44][31].run()  ;
            end
            begin
              drv[44][31].run()  ;
            end
            begin
              mem_check[44][31].run()  ;
            end
            begin
              rf_driver[44][31].run()  ;
            end

            begin
              ldst_driver[45].run()  ;
            end
            begin
              mgr[45].run()  ;
            end
            begin
              oob_drv[45].run()  ;
            end
            begin
              up_check[45].run()  ;
            end
            begin
              gen[45][0].run()  ;
            end
            begin
              drv[45][0].run()  ;
            end
            begin
              mem_check[45][0].run()  ;
            end
            begin
              rf_driver[45][0].run()  ;
            end

            begin
              gen[45][1].run()  ;
            end
            begin
              drv[45][1].run()  ;
            end
            begin
              mem_check[45][1].run()  ;
            end
            begin
              rf_driver[45][1].run()  ;
            end

            begin
              gen[45][2].run()  ;
            end
            begin
              drv[45][2].run()  ;
            end
            begin
              mem_check[45][2].run()  ;
            end
            begin
              rf_driver[45][2].run()  ;
            end

            begin
              gen[45][3].run()  ;
            end
            begin
              drv[45][3].run()  ;
            end
            begin
              mem_check[45][3].run()  ;
            end
            begin
              rf_driver[45][3].run()  ;
            end

            begin
              gen[45][4].run()  ;
            end
            begin
              drv[45][4].run()  ;
            end
            begin
              mem_check[45][4].run()  ;
            end
            begin
              rf_driver[45][4].run()  ;
            end

            begin
              gen[45][5].run()  ;
            end
            begin
              drv[45][5].run()  ;
            end
            begin
              mem_check[45][5].run()  ;
            end
            begin
              rf_driver[45][5].run()  ;
            end

            begin
              gen[45][6].run()  ;
            end
            begin
              drv[45][6].run()  ;
            end
            begin
              mem_check[45][6].run()  ;
            end
            begin
              rf_driver[45][6].run()  ;
            end

            begin
              gen[45][7].run()  ;
            end
            begin
              drv[45][7].run()  ;
            end
            begin
              mem_check[45][7].run()  ;
            end
            begin
              rf_driver[45][7].run()  ;
            end

            begin
              gen[45][8].run()  ;
            end
            begin
              drv[45][8].run()  ;
            end
            begin
              mem_check[45][8].run()  ;
            end
            begin
              rf_driver[45][8].run()  ;
            end

            begin
              gen[45][9].run()  ;
            end
            begin
              drv[45][9].run()  ;
            end
            begin
              mem_check[45][9].run()  ;
            end
            begin
              rf_driver[45][9].run()  ;
            end

            begin
              gen[45][10].run()  ;
            end
            begin
              drv[45][10].run()  ;
            end
            begin
              mem_check[45][10].run()  ;
            end
            begin
              rf_driver[45][10].run()  ;
            end

            begin
              gen[45][11].run()  ;
            end
            begin
              drv[45][11].run()  ;
            end
            begin
              mem_check[45][11].run()  ;
            end
            begin
              rf_driver[45][11].run()  ;
            end

            begin
              gen[45][12].run()  ;
            end
            begin
              drv[45][12].run()  ;
            end
            begin
              mem_check[45][12].run()  ;
            end
            begin
              rf_driver[45][12].run()  ;
            end

            begin
              gen[45][13].run()  ;
            end
            begin
              drv[45][13].run()  ;
            end
            begin
              mem_check[45][13].run()  ;
            end
            begin
              rf_driver[45][13].run()  ;
            end

            begin
              gen[45][14].run()  ;
            end
            begin
              drv[45][14].run()  ;
            end
            begin
              mem_check[45][14].run()  ;
            end
            begin
              rf_driver[45][14].run()  ;
            end

            begin
              gen[45][15].run()  ;
            end
            begin
              drv[45][15].run()  ;
            end
            begin
              mem_check[45][15].run()  ;
            end
            begin
              rf_driver[45][15].run()  ;
            end

            begin
              gen[45][16].run()  ;
            end
            begin
              drv[45][16].run()  ;
            end
            begin
              mem_check[45][16].run()  ;
            end
            begin
              rf_driver[45][16].run()  ;
            end

            begin
              gen[45][17].run()  ;
            end
            begin
              drv[45][17].run()  ;
            end
            begin
              mem_check[45][17].run()  ;
            end
            begin
              rf_driver[45][17].run()  ;
            end

            begin
              gen[45][18].run()  ;
            end
            begin
              drv[45][18].run()  ;
            end
            begin
              mem_check[45][18].run()  ;
            end
            begin
              rf_driver[45][18].run()  ;
            end

            begin
              gen[45][19].run()  ;
            end
            begin
              drv[45][19].run()  ;
            end
            begin
              mem_check[45][19].run()  ;
            end
            begin
              rf_driver[45][19].run()  ;
            end

            begin
              gen[45][20].run()  ;
            end
            begin
              drv[45][20].run()  ;
            end
            begin
              mem_check[45][20].run()  ;
            end
            begin
              rf_driver[45][20].run()  ;
            end

            begin
              gen[45][21].run()  ;
            end
            begin
              drv[45][21].run()  ;
            end
            begin
              mem_check[45][21].run()  ;
            end
            begin
              rf_driver[45][21].run()  ;
            end

            begin
              gen[45][22].run()  ;
            end
            begin
              drv[45][22].run()  ;
            end
            begin
              mem_check[45][22].run()  ;
            end
            begin
              rf_driver[45][22].run()  ;
            end

            begin
              gen[45][23].run()  ;
            end
            begin
              drv[45][23].run()  ;
            end
            begin
              mem_check[45][23].run()  ;
            end
            begin
              rf_driver[45][23].run()  ;
            end

            begin
              gen[45][24].run()  ;
            end
            begin
              drv[45][24].run()  ;
            end
            begin
              mem_check[45][24].run()  ;
            end
            begin
              rf_driver[45][24].run()  ;
            end

            begin
              gen[45][25].run()  ;
            end
            begin
              drv[45][25].run()  ;
            end
            begin
              mem_check[45][25].run()  ;
            end
            begin
              rf_driver[45][25].run()  ;
            end

            begin
              gen[45][26].run()  ;
            end
            begin
              drv[45][26].run()  ;
            end
            begin
              mem_check[45][26].run()  ;
            end
            begin
              rf_driver[45][26].run()  ;
            end

            begin
              gen[45][27].run()  ;
            end
            begin
              drv[45][27].run()  ;
            end
            begin
              mem_check[45][27].run()  ;
            end
            begin
              rf_driver[45][27].run()  ;
            end

            begin
              gen[45][28].run()  ;
            end
            begin
              drv[45][28].run()  ;
            end
            begin
              mem_check[45][28].run()  ;
            end
            begin
              rf_driver[45][28].run()  ;
            end

            begin
              gen[45][29].run()  ;
            end
            begin
              drv[45][29].run()  ;
            end
            begin
              mem_check[45][29].run()  ;
            end
            begin
              rf_driver[45][29].run()  ;
            end

            begin
              gen[45][30].run()  ;
            end
            begin
              drv[45][30].run()  ;
            end
            begin
              mem_check[45][30].run()  ;
            end
            begin
              rf_driver[45][30].run()  ;
            end

            begin
              gen[45][31].run()  ;
            end
            begin
              drv[45][31].run()  ;
            end
            begin
              mem_check[45][31].run()  ;
            end
            begin
              rf_driver[45][31].run()  ;
            end

            begin
              ldst_driver[46].run()  ;
            end
            begin
              mgr[46].run()  ;
            end
            begin
              oob_drv[46].run()  ;
            end
            begin
              up_check[46].run()  ;
            end
            begin
              gen[46][0].run()  ;
            end
            begin
              drv[46][0].run()  ;
            end
            begin
              mem_check[46][0].run()  ;
            end
            begin
              rf_driver[46][0].run()  ;
            end

            begin
              gen[46][1].run()  ;
            end
            begin
              drv[46][1].run()  ;
            end
            begin
              mem_check[46][1].run()  ;
            end
            begin
              rf_driver[46][1].run()  ;
            end

            begin
              gen[46][2].run()  ;
            end
            begin
              drv[46][2].run()  ;
            end
            begin
              mem_check[46][2].run()  ;
            end
            begin
              rf_driver[46][2].run()  ;
            end

            begin
              gen[46][3].run()  ;
            end
            begin
              drv[46][3].run()  ;
            end
            begin
              mem_check[46][3].run()  ;
            end
            begin
              rf_driver[46][3].run()  ;
            end

            begin
              gen[46][4].run()  ;
            end
            begin
              drv[46][4].run()  ;
            end
            begin
              mem_check[46][4].run()  ;
            end
            begin
              rf_driver[46][4].run()  ;
            end

            begin
              gen[46][5].run()  ;
            end
            begin
              drv[46][5].run()  ;
            end
            begin
              mem_check[46][5].run()  ;
            end
            begin
              rf_driver[46][5].run()  ;
            end

            begin
              gen[46][6].run()  ;
            end
            begin
              drv[46][6].run()  ;
            end
            begin
              mem_check[46][6].run()  ;
            end
            begin
              rf_driver[46][6].run()  ;
            end

            begin
              gen[46][7].run()  ;
            end
            begin
              drv[46][7].run()  ;
            end
            begin
              mem_check[46][7].run()  ;
            end
            begin
              rf_driver[46][7].run()  ;
            end

            begin
              gen[46][8].run()  ;
            end
            begin
              drv[46][8].run()  ;
            end
            begin
              mem_check[46][8].run()  ;
            end
            begin
              rf_driver[46][8].run()  ;
            end

            begin
              gen[46][9].run()  ;
            end
            begin
              drv[46][9].run()  ;
            end
            begin
              mem_check[46][9].run()  ;
            end
            begin
              rf_driver[46][9].run()  ;
            end

            begin
              gen[46][10].run()  ;
            end
            begin
              drv[46][10].run()  ;
            end
            begin
              mem_check[46][10].run()  ;
            end
            begin
              rf_driver[46][10].run()  ;
            end

            begin
              gen[46][11].run()  ;
            end
            begin
              drv[46][11].run()  ;
            end
            begin
              mem_check[46][11].run()  ;
            end
            begin
              rf_driver[46][11].run()  ;
            end

            begin
              gen[46][12].run()  ;
            end
            begin
              drv[46][12].run()  ;
            end
            begin
              mem_check[46][12].run()  ;
            end
            begin
              rf_driver[46][12].run()  ;
            end

            begin
              gen[46][13].run()  ;
            end
            begin
              drv[46][13].run()  ;
            end
            begin
              mem_check[46][13].run()  ;
            end
            begin
              rf_driver[46][13].run()  ;
            end

            begin
              gen[46][14].run()  ;
            end
            begin
              drv[46][14].run()  ;
            end
            begin
              mem_check[46][14].run()  ;
            end
            begin
              rf_driver[46][14].run()  ;
            end

            begin
              gen[46][15].run()  ;
            end
            begin
              drv[46][15].run()  ;
            end
            begin
              mem_check[46][15].run()  ;
            end
            begin
              rf_driver[46][15].run()  ;
            end

            begin
              gen[46][16].run()  ;
            end
            begin
              drv[46][16].run()  ;
            end
            begin
              mem_check[46][16].run()  ;
            end
            begin
              rf_driver[46][16].run()  ;
            end

            begin
              gen[46][17].run()  ;
            end
            begin
              drv[46][17].run()  ;
            end
            begin
              mem_check[46][17].run()  ;
            end
            begin
              rf_driver[46][17].run()  ;
            end

            begin
              gen[46][18].run()  ;
            end
            begin
              drv[46][18].run()  ;
            end
            begin
              mem_check[46][18].run()  ;
            end
            begin
              rf_driver[46][18].run()  ;
            end

            begin
              gen[46][19].run()  ;
            end
            begin
              drv[46][19].run()  ;
            end
            begin
              mem_check[46][19].run()  ;
            end
            begin
              rf_driver[46][19].run()  ;
            end

            begin
              gen[46][20].run()  ;
            end
            begin
              drv[46][20].run()  ;
            end
            begin
              mem_check[46][20].run()  ;
            end
            begin
              rf_driver[46][20].run()  ;
            end

            begin
              gen[46][21].run()  ;
            end
            begin
              drv[46][21].run()  ;
            end
            begin
              mem_check[46][21].run()  ;
            end
            begin
              rf_driver[46][21].run()  ;
            end

            begin
              gen[46][22].run()  ;
            end
            begin
              drv[46][22].run()  ;
            end
            begin
              mem_check[46][22].run()  ;
            end
            begin
              rf_driver[46][22].run()  ;
            end

            begin
              gen[46][23].run()  ;
            end
            begin
              drv[46][23].run()  ;
            end
            begin
              mem_check[46][23].run()  ;
            end
            begin
              rf_driver[46][23].run()  ;
            end

            begin
              gen[46][24].run()  ;
            end
            begin
              drv[46][24].run()  ;
            end
            begin
              mem_check[46][24].run()  ;
            end
            begin
              rf_driver[46][24].run()  ;
            end

            begin
              gen[46][25].run()  ;
            end
            begin
              drv[46][25].run()  ;
            end
            begin
              mem_check[46][25].run()  ;
            end
            begin
              rf_driver[46][25].run()  ;
            end

            begin
              gen[46][26].run()  ;
            end
            begin
              drv[46][26].run()  ;
            end
            begin
              mem_check[46][26].run()  ;
            end
            begin
              rf_driver[46][26].run()  ;
            end

            begin
              gen[46][27].run()  ;
            end
            begin
              drv[46][27].run()  ;
            end
            begin
              mem_check[46][27].run()  ;
            end
            begin
              rf_driver[46][27].run()  ;
            end

            begin
              gen[46][28].run()  ;
            end
            begin
              drv[46][28].run()  ;
            end
            begin
              mem_check[46][28].run()  ;
            end
            begin
              rf_driver[46][28].run()  ;
            end

            begin
              gen[46][29].run()  ;
            end
            begin
              drv[46][29].run()  ;
            end
            begin
              mem_check[46][29].run()  ;
            end
            begin
              rf_driver[46][29].run()  ;
            end

            begin
              gen[46][30].run()  ;
            end
            begin
              drv[46][30].run()  ;
            end
            begin
              mem_check[46][30].run()  ;
            end
            begin
              rf_driver[46][30].run()  ;
            end

            begin
              gen[46][31].run()  ;
            end
            begin
              drv[46][31].run()  ;
            end
            begin
              mem_check[46][31].run()  ;
            end
            begin
              rf_driver[46][31].run()  ;
            end

            begin
              ldst_driver[47].run()  ;
            end
            begin
              mgr[47].run()  ;
            end
            begin
              oob_drv[47].run()  ;
            end
            begin
              up_check[47].run()  ;
            end
            begin
              gen[47][0].run()  ;
            end
            begin
              drv[47][0].run()  ;
            end
            begin
              mem_check[47][0].run()  ;
            end
            begin
              rf_driver[47][0].run()  ;
            end

            begin
              gen[47][1].run()  ;
            end
            begin
              drv[47][1].run()  ;
            end
            begin
              mem_check[47][1].run()  ;
            end
            begin
              rf_driver[47][1].run()  ;
            end

            begin
              gen[47][2].run()  ;
            end
            begin
              drv[47][2].run()  ;
            end
            begin
              mem_check[47][2].run()  ;
            end
            begin
              rf_driver[47][2].run()  ;
            end

            begin
              gen[47][3].run()  ;
            end
            begin
              drv[47][3].run()  ;
            end
            begin
              mem_check[47][3].run()  ;
            end
            begin
              rf_driver[47][3].run()  ;
            end

            begin
              gen[47][4].run()  ;
            end
            begin
              drv[47][4].run()  ;
            end
            begin
              mem_check[47][4].run()  ;
            end
            begin
              rf_driver[47][4].run()  ;
            end

            begin
              gen[47][5].run()  ;
            end
            begin
              drv[47][5].run()  ;
            end
            begin
              mem_check[47][5].run()  ;
            end
            begin
              rf_driver[47][5].run()  ;
            end

            begin
              gen[47][6].run()  ;
            end
            begin
              drv[47][6].run()  ;
            end
            begin
              mem_check[47][6].run()  ;
            end
            begin
              rf_driver[47][6].run()  ;
            end

            begin
              gen[47][7].run()  ;
            end
            begin
              drv[47][7].run()  ;
            end
            begin
              mem_check[47][7].run()  ;
            end
            begin
              rf_driver[47][7].run()  ;
            end

            begin
              gen[47][8].run()  ;
            end
            begin
              drv[47][8].run()  ;
            end
            begin
              mem_check[47][8].run()  ;
            end
            begin
              rf_driver[47][8].run()  ;
            end

            begin
              gen[47][9].run()  ;
            end
            begin
              drv[47][9].run()  ;
            end
            begin
              mem_check[47][9].run()  ;
            end
            begin
              rf_driver[47][9].run()  ;
            end

            begin
              gen[47][10].run()  ;
            end
            begin
              drv[47][10].run()  ;
            end
            begin
              mem_check[47][10].run()  ;
            end
            begin
              rf_driver[47][10].run()  ;
            end

            begin
              gen[47][11].run()  ;
            end
            begin
              drv[47][11].run()  ;
            end
            begin
              mem_check[47][11].run()  ;
            end
            begin
              rf_driver[47][11].run()  ;
            end

            begin
              gen[47][12].run()  ;
            end
            begin
              drv[47][12].run()  ;
            end
            begin
              mem_check[47][12].run()  ;
            end
            begin
              rf_driver[47][12].run()  ;
            end

            begin
              gen[47][13].run()  ;
            end
            begin
              drv[47][13].run()  ;
            end
            begin
              mem_check[47][13].run()  ;
            end
            begin
              rf_driver[47][13].run()  ;
            end

            begin
              gen[47][14].run()  ;
            end
            begin
              drv[47][14].run()  ;
            end
            begin
              mem_check[47][14].run()  ;
            end
            begin
              rf_driver[47][14].run()  ;
            end

            begin
              gen[47][15].run()  ;
            end
            begin
              drv[47][15].run()  ;
            end
            begin
              mem_check[47][15].run()  ;
            end
            begin
              rf_driver[47][15].run()  ;
            end

            begin
              gen[47][16].run()  ;
            end
            begin
              drv[47][16].run()  ;
            end
            begin
              mem_check[47][16].run()  ;
            end
            begin
              rf_driver[47][16].run()  ;
            end

            begin
              gen[47][17].run()  ;
            end
            begin
              drv[47][17].run()  ;
            end
            begin
              mem_check[47][17].run()  ;
            end
            begin
              rf_driver[47][17].run()  ;
            end

            begin
              gen[47][18].run()  ;
            end
            begin
              drv[47][18].run()  ;
            end
            begin
              mem_check[47][18].run()  ;
            end
            begin
              rf_driver[47][18].run()  ;
            end

            begin
              gen[47][19].run()  ;
            end
            begin
              drv[47][19].run()  ;
            end
            begin
              mem_check[47][19].run()  ;
            end
            begin
              rf_driver[47][19].run()  ;
            end

            begin
              gen[47][20].run()  ;
            end
            begin
              drv[47][20].run()  ;
            end
            begin
              mem_check[47][20].run()  ;
            end
            begin
              rf_driver[47][20].run()  ;
            end

            begin
              gen[47][21].run()  ;
            end
            begin
              drv[47][21].run()  ;
            end
            begin
              mem_check[47][21].run()  ;
            end
            begin
              rf_driver[47][21].run()  ;
            end

            begin
              gen[47][22].run()  ;
            end
            begin
              drv[47][22].run()  ;
            end
            begin
              mem_check[47][22].run()  ;
            end
            begin
              rf_driver[47][22].run()  ;
            end

            begin
              gen[47][23].run()  ;
            end
            begin
              drv[47][23].run()  ;
            end
            begin
              mem_check[47][23].run()  ;
            end
            begin
              rf_driver[47][23].run()  ;
            end

            begin
              gen[47][24].run()  ;
            end
            begin
              drv[47][24].run()  ;
            end
            begin
              mem_check[47][24].run()  ;
            end
            begin
              rf_driver[47][24].run()  ;
            end

            begin
              gen[47][25].run()  ;
            end
            begin
              drv[47][25].run()  ;
            end
            begin
              mem_check[47][25].run()  ;
            end
            begin
              rf_driver[47][25].run()  ;
            end

            begin
              gen[47][26].run()  ;
            end
            begin
              drv[47][26].run()  ;
            end
            begin
              mem_check[47][26].run()  ;
            end
            begin
              rf_driver[47][26].run()  ;
            end

            begin
              gen[47][27].run()  ;
            end
            begin
              drv[47][27].run()  ;
            end
            begin
              mem_check[47][27].run()  ;
            end
            begin
              rf_driver[47][27].run()  ;
            end

            begin
              gen[47][28].run()  ;
            end
            begin
              drv[47][28].run()  ;
            end
            begin
              mem_check[47][28].run()  ;
            end
            begin
              rf_driver[47][28].run()  ;
            end

            begin
              gen[47][29].run()  ;
            end
            begin
              drv[47][29].run()  ;
            end
            begin
              mem_check[47][29].run()  ;
            end
            begin
              rf_driver[47][29].run()  ;
            end

            begin
              gen[47][30].run()  ;
            end
            begin
              drv[47][30].run()  ;
            end
            begin
              mem_check[47][30].run()  ;
            end
            begin
              rf_driver[47][30].run()  ;
            end

            begin
              gen[47][31].run()  ;
            end
            begin
              drv[47][31].run()  ;
            end
            begin
              mem_check[47][31].run()  ;
            end
            begin
              rf_driver[47][31].run()  ;
            end

            begin
              ldst_driver[48].run()  ;
            end
            begin
              mgr[48].run()  ;
            end
            begin
              oob_drv[48].run()  ;
            end
            begin
              up_check[48].run()  ;
            end
            begin
              gen[48][0].run()  ;
            end
            begin
              drv[48][0].run()  ;
            end
            begin
              mem_check[48][0].run()  ;
            end
            begin
              rf_driver[48][0].run()  ;
            end

            begin
              gen[48][1].run()  ;
            end
            begin
              drv[48][1].run()  ;
            end
            begin
              mem_check[48][1].run()  ;
            end
            begin
              rf_driver[48][1].run()  ;
            end

            begin
              gen[48][2].run()  ;
            end
            begin
              drv[48][2].run()  ;
            end
            begin
              mem_check[48][2].run()  ;
            end
            begin
              rf_driver[48][2].run()  ;
            end

            begin
              gen[48][3].run()  ;
            end
            begin
              drv[48][3].run()  ;
            end
            begin
              mem_check[48][3].run()  ;
            end
            begin
              rf_driver[48][3].run()  ;
            end

            begin
              gen[48][4].run()  ;
            end
            begin
              drv[48][4].run()  ;
            end
            begin
              mem_check[48][4].run()  ;
            end
            begin
              rf_driver[48][4].run()  ;
            end

            begin
              gen[48][5].run()  ;
            end
            begin
              drv[48][5].run()  ;
            end
            begin
              mem_check[48][5].run()  ;
            end
            begin
              rf_driver[48][5].run()  ;
            end

            begin
              gen[48][6].run()  ;
            end
            begin
              drv[48][6].run()  ;
            end
            begin
              mem_check[48][6].run()  ;
            end
            begin
              rf_driver[48][6].run()  ;
            end

            begin
              gen[48][7].run()  ;
            end
            begin
              drv[48][7].run()  ;
            end
            begin
              mem_check[48][7].run()  ;
            end
            begin
              rf_driver[48][7].run()  ;
            end

            begin
              gen[48][8].run()  ;
            end
            begin
              drv[48][8].run()  ;
            end
            begin
              mem_check[48][8].run()  ;
            end
            begin
              rf_driver[48][8].run()  ;
            end

            begin
              gen[48][9].run()  ;
            end
            begin
              drv[48][9].run()  ;
            end
            begin
              mem_check[48][9].run()  ;
            end
            begin
              rf_driver[48][9].run()  ;
            end

            begin
              gen[48][10].run()  ;
            end
            begin
              drv[48][10].run()  ;
            end
            begin
              mem_check[48][10].run()  ;
            end
            begin
              rf_driver[48][10].run()  ;
            end

            begin
              gen[48][11].run()  ;
            end
            begin
              drv[48][11].run()  ;
            end
            begin
              mem_check[48][11].run()  ;
            end
            begin
              rf_driver[48][11].run()  ;
            end

            begin
              gen[48][12].run()  ;
            end
            begin
              drv[48][12].run()  ;
            end
            begin
              mem_check[48][12].run()  ;
            end
            begin
              rf_driver[48][12].run()  ;
            end

            begin
              gen[48][13].run()  ;
            end
            begin
              drv[48][13].run()  ;
            end
            begin
              mem_check[48][13].run()  ;
            end
            begin
              rf_driver[48][13].run()  ;
            end

            begin
              gen[48][14].run()  ;
            end
            begin
              drv[48][14].run()  ;
            end
            begin
              mem_check[48][14].run()  ;
            end
            begin
              rf_driver[48][14].run()  ;
            end

            begin
              gen[48][15].run()  ;
            end
            begin
              drv[48][15].run()  ;
            end
            begin
              mem_check[48][15].run()  ;
            end
            begin
              rf_driver[48][15].run()  ;
            end

            begin
              gen[48][16].run()  ;
            end
            begin
              drv[48][16].run()  ;
            end
            begin
              mem_check[48][16].run()  ;
            end
            begin
              rf_driver[48][16].run()  ;
            end

            begin
              gen[48][17].run()  ;
            end
            begin
              drv[48][17].run()  ;
            end
            begin
              mem_check[48][17].run()  ;
            end
            begin
              rf_driver[48][17].run()  ;
            end

            begin
              gen[48][18].run()  ;
            end
            begin
              drv[48][18].run()  ;
            end
            begin
              mem_check[48][18].run()  ;
            end
            begin
              rf_driver[48][18].run()  ;
            end

            begin
              gen[48][19].run()  ;
            end
            begin
              drv[48][19].run()  ;
            end
            begin
              mem_check[48][19].run()  ;
            end
            begin
              rf_driver[48][19].run()  ;
            end

            begin
              gen[48][20].run()  ;
            end
            begin
              drv[48][20].run()  ;
            end
            begin
              mem_check[48][20].run()  ;
            end
            begin
              rf_driver[48][20].run()  ;
            end

            begin
              gen[48][21].run()  ;
            end
            begin
              drv[48][21].run()  ;
            end
            begin
              mem_check[48][21].run()  ;
            end
            begin
              rf_driver[48][21].run()  ;
            end

            begin
              gen[48][22].run()  ;
            end
            begin
              drv[48][22].run()  ;
            end
            begin
              mem_check[48][22].run()  ;
            end
            begin
              rf_driver[48][22].run()  ;
            end

            begin
              gen[48][23].run()  ;
            end
            begin
              drv[48][23].run()  ;
            end
            begin
              mem_check[48][23].run()  ;
            end
            begin
              rf_driver[48][23].run()  ;
            end

            begin
              gen[48][24].run()  ;
            end
            begin
              drv[48][24].run()  ;
            end
            begin
              mem_check[48][24].run()  ;
            end
            begin
              rf_driver[48][24].run()  ;
            end

            begin
              gen[48][25].run()  ;
            end
            begin
              drv[48][25].run()  ;
            end
            begin
              mem_check[48][25].run()  ;
            end
            begin
              rf_driver[48][25].run()  ;
            end

            begin
              gen[48][26].run()  ;
            end
            begin
              drv[48][26].run()  ;
            end
            begin
              mem_check[48][26].run()  ;
            end
            begin
              rf_driver[48][26].run()  ;
            end

            begin
              gen[48][27].run()  ;
            end
            begin
              drv[48][27].run()  ;
            end
            begin
              mem_check[48][27].run()  ;
            end
            begin
              rf_driver[48][27].run()  ;
            end

            begin
              gen[48][28].run()  ;
            end
            begin
              drv[48][28].run()  ;
            end
            begin
              mem_check[48][28].run()  ;
            end
            begin
              rf_driver[48][28].run()  ;
            end

            begin
              gen[48][29].run()  ;
            end
            begin
              drv[48][29].run()  ;
            end
            begin
              mem_check[48][29].run()  ;
            end
            begin
              rf_driver[48][29].run()  ;
            end

            begin
              gen[48][30].run()  ;
            end
            begin
              drv[48][30].run()  ;
            end
            begin
              mem_check[48][30].run()  ;
            end
            begin
              rf_driver[48][30].run()  ;
            end

            begin
              gen[48][31].run()  ;
            end
            begin
              drv[48][31].run()  ;
            end
            begin
              mem_check[48][31].run()  ;
            end
            begin
              rf_driver[48][31].run()  ;
            end

            begin
              ldst_driver[49].run()  ;
            end
            begin
              mgr[49].run()  ;
            end
            begin
              oob_drv[49].run()  ;
            end
            begin
              up_check[49].run()  ;
            end
            begin
              gen[49][0].run()  ;
            end
            begin
              drv[49][0].run()  ;
            end
            begin
              mem_check[49][0].run()  ;
            end
            begin
              rf_driver[49][0].run()  ;
            end

            begin
              gen[49][1].run()  ;
            end
            begin
              drv[49][1].run()  ;
            end
            begin
              mem_check[49][1].run()  ;
            end
            begin
              rf_driver[49][1].run()  ;
            end

            begin
              gen[49][2].run()  ;
            end
            begin
              drv[49][2].run()  ;
            end
            begin
              mem_check[49][2].run()  ;
            end
            begin
              rf_driver[49][2].run()  ;
            end

            begin
              gen[49][3].run()  ;
            end
            begin
              drv[49][3].run()  ;
            end
            begin
              mem_check[49][3].run()  ;
            end
            begin
              rf_driver[49][3].run()  ;
            end

            begin
              gen[49][4].run()  ;
            end
            begin
              drv[49][4].run()  ;
            end
            begin
              mem_check[49][4].run()  ;
            end
            begin
              rf_driver[49][4].run()  ;
            end

            begin
              gen[49][5].run()  ;
            end
            begin
              drv[49][5].run()  ;
            end
            begin
              mem_check[49][5].run()  ;
            end
            begin
              rf_driver[49][5].run()  ;
            end

            begin
              gen[49][6].run()  ;
            end
            begin
              drv[49][6].run()  ;
            end
            begin
              mem_check[49][6].run()  ;
            end
            begin
              rf_driver[49][6].run()  ;
            end

            begin
              gen[49][7].run()  ;
            end
            begin
              drv[49][7].run()  ;
            end
            begin
              mem_check[49][7].run()  ;
            end
            begin
              rf_driver[49][7].run()  ;
            end

            begin
              gen[49][8].run()  ;
            end
            begin
              drv[49][8].run()  ;
            end
            begin
              mem_check[49][8].run()  ;
            end
            begin
              rf_driver[49][8].run()  ;
            end

            begin
              gen[49][9].run()  ;
            end
            begin
              drv[49][9].run()  ;
            end
            begin
              mem_check[49][9].run()  ;
            end
            begin
              rf_driver[49][9].run()  ;
            end

            begin
              gen[49][10].run()  ;
            end
            begin
              drv[49][10].run()  ;
            end
            begin
              mem_check[49][10].run()  ;
            end
            begin
              rf_driver[49][10].run()  ;
            end

            begin
              gen[49][11].run()  ;
            end
            begin
              drv[49][11].run()  ;
            end
            begin
              mem_check[49][11].run()  ;
            end
            begin
              rf_driver[49][11].run()  ;
            end

            begin
              gen[49][12].run()  ;
            end
            begin
              drv[49][12].run()  ;
            end
            begin
              mem_check[49][12].run()  ;
            end
            begin
              rf_driver[49][12].run()  ;
            end

            begin
              gen[49][13].run()  ;
            end
            begin
              drv[49][13].run()  ;
            end
            begin
              mem_check[49][13].run()  ;
            end
            begin
              rf_driver[49][13].run()  ;
            end

            begin
              gen[49][14].run()  ;
            end
            begin
              drv[49][14].run()  ;
            end
            begin
              mem_check[49][14].run()  ;
            end
            begin
              rf_driver[49][14].run()  ;
            end

            begin
              gen[49][15].run()  ;
            end
            begin
              drv[49][15].run()  ;
            end
            begin
              mem_check[49][15].run()  ;
            end
            begin
              rf_driver[49][15].run()  ;
            end

            begin
              gen[49][16].run()  ;
            end
            begin
              drv[49][16].run()  ;
            end
            begin
              mem_check[49][16].run()  ;
            end
            begin
              rf_driver[49][16].run()  ;
            end

            begin
              gen[49][17].run()  ;
            end
            begin
              drv[49][17].run()  ;
            end
            begin
              mem_check[49][17].run()  ;
            end
            begin
              rf_driver[49][17].run()  ;
            end

            begin
              gen[49][18].run()  ;
            end
            begin
              drv[49][18].run()  ;
            end
            begin
              mem_check[49][18].run()  ;
            end
            begin
              rf_driver[49][18].run()  ;
            end

            begin
              gen[49][19].run()  ;
            end
            begin
              drv[49][19].run()  ;
            end
            begin
              mem_check[49][19].run()  ;
            end
            begin
              rf_driver[49][19].run()  ;
            end

            begin
              gen[49][20].run()  ;
            end
            begin
              drv[49][20].run()  ;
            end
            begin
              mem_check[49][20].run()  ;
            end
            begin
              rf_driver[49][20].run()  ;
            end

            begin
              gen[49][21].run()  ;
            end
            begin
              drv[49][21].run()  ;
            end
            begin
              mem_check[49][21].run()  ;
            end
            begin
              rf_driver[49][21].run()  ;
            end

            begin
              gen[49][22].run()  ;
            end
            begin
              drv[49][22].run()  ;
            end
            begin
              mem_check[49][22].run()  ;
            end
            begin
              rf_driver[49][22].run()  ;
            end

            begin
              gen[49][23].run()  ;
            end
            begin
              drv[49][23].run()  ;
            end
            begin
              mem_check[49][23].run()  ;
            end
            begin
              rf_driver[49][23].run()  ;
            end

            begin
              gen[49][24].run()  ;
            end
            begin
              drv[49][24].run()  ;
            end
            begin
              mem_check[49][24].run()  ;
            end
            begin
              rf_driver[49][24].run()  ;
            end

            begin
              gen[49][25].run()  ;
            end
            begin
              drv[49][25].run()  ;
            end
            begin
              mem_check[49][25].run()  ;
            end
            begin
              rf_driver[49][25].run()  ;
            end

            begin
              gen[49][26].run()  ;
            end
            begin
              drv[49][26].run()  ;
            end
            begin
              mem_check[49][26].run()  ;
            end
            begin
              rf_driver[49][26].run()  ;
            end

            begin
              gen[49][27].run()  ;
            end
            begin
              drv[49][27].run()  ;
            end
            begin
              mem_check[49][27].run()  ;
            end
            begin
              rf_driver[49][27].run()  ;
            end

            begin
              gen[49][28].run()  ;
            end
            begin
              drv[49][28].run()  ;
            end
            begin
              mem_check[49][28].run()  ;
            end
            begin
              rf_driver[49][28].run()  ;
            end

            begin
              gen[49][29].run()  ;
            end
            begin
              drv[49][29].run()  ;
            end
            begin
              mem_check[49][29].run()  ;
            end
            begin
              rf_driver[49][29].run()  ;
            end

            begin
              gen[49][30].run()  ;
            end
            begin
              drv[49][30].run()  ;
            end
            begin
              mem_check[49][30].run()  ;
            end
            begin
              rf_driver[49][30].run()  ;
            end

            begin
              gen[49][31].run()  ;
            end
            begin
              drv[49][31].run()  ;
            end
            begin
              mem_check[49][31].run()  ;
            end
            begin
              rf_driver[49][31].run()  ;
            end

            begin
              ldst_driver[50].run()  ;
            end
            begin
              mgr[50].run()  ;
            end
            begin
              oob_drv[50].run()  ;
            end
            begin
              up_check[50].run()  ;
            end
            begin
              gen[50][0].run()  ;
            end
            begin
              drv[50][0].run()  ;
            end
            begin
              mem_check[50][0].run()  ;
            end
            begin
              rf_driver[50][0].run()  ;
            end

            begin
              gen[50][1].run()  ;
            end
            begin
              drv[50][1].run()  ;
            end
            begin
              mem_check[50][1].run()  ;
            end
            begin
              rf_driver[50][1].run()  ;
            end

            begin
              gen[50][2].run()  ;
            end
            begin
              drv[50][2].run()  ;
            end
            begin
              mem_check[50][2].run()  ;
            end
            begin
              rf_driver[50][2].run()  ;
            end

            begin
              gen[50][3].run()  ;
            end
            begin
              drv[50][3].run()  ;
            end
            begin
              mem_check[50][3].run()  ;
            end
            begin
              rf_driver[50][3].run()  ;
            end

            begin
              gen[50][4].run()  ;
            end
            begin
              drv[50][4].run()  ;
            end
            begin
              mem_check[50][4].run()  ;
            end
            begin
              rf_driver[50][4].run()  ;
            end

            begin
              gen[50][5].run()  ;
            end
            begin
              drv[50][5].run()  ;
            end
            begin
              mem_check[50][5].run()  ;
            end
            begin
              rf_driver[50][5].run()  ;
            end

            begin
              gen[50][6].run()  ;
            end
            begin
              drv[50][6].run()  ;
            end
            begin
              mem_check[50][6].run()  ;
            end
            begin
              rf_driver[50][6].run()  ;
            end

            begin
              gen[50][7].run()  ;
            end
            begin
              drv[50][7].run()  ;
            end
            begin
              mem_check[50][7].run()  ;
            end
            begin
              rf_driver[50][7].run()  ;
            end

            begin
              gen[50][8].run()  ;
            end
            begin
              drv[50][8].run()  ;
            end
            begin
              mem_check[50][8].run()  ;
            end
            begin
              rf_driver[50][8].run()  ;
            end

            begin
              gen[50][9].run()  ;
            end
            begin
              drv[50][9].run()  ;
            end
            begin
              mem_check[50][9].run()  ;
            end
            begin
              rf_driver[50][9].run()  ;
            end

            begin
              gen[50][10].run()  ;
            end
            begin
              drv[50][10].run()  ;
            end
            begin
              mem_check[50][10].run()  ;
            end
            begin
              rf_driver[50][10].run()  ;
            end

            begin
              gen[50][11].run()  ;
            end
            begin
              drv[50][11].run()  ;
            end
            begin
              mem_check[50][11].run()  ;
            end
            begin
              rf_driver[50][11].run()  ;
            end

            begin
              gen[50][12].run()  ;
            end
            begin
              drv[50][12].run()  ;
            end
            begin
              mem_check[50][12].run()  ;
            end
            begin
              rf_driver[50][12].run()  ;
            end

            begin
              gen[50][13].run()  ;
            end
            begin
              drv[50][13].run()  ;
            end
            begin
              mem_check[50][13].run()  ;
            end
            begin
              rf_driver[50][13].run()  ;
            end

            begin
              gen[50][14].run()  ;
            end
            begin
              drv[50][14].run()  ;
            end
            begin
              mem_check[50][14].run()  ;
            end
            begin
              rf_driver[50][14].run()  ;
            end

            begin
              gen[50][15].run()  ;
            end
            begin
              drv[50][15].run()  ;
            end
            begin
              mem_check[50][15].run()  ;
            end
            begin
              rf_driver[50][15].run()  ;
            end

            begin
              gen[50][16].run()  ;
            end
            begin
              drv[50][16].run()  ;
            end
            begin
              mem_check[50][16].run()  ;
            end
            begin
              rf_driver[50][16].run()  ;
            end

            begin
              gen[50][17].run()  ;
            end
            begin
              drv[50][17].run()  ;
            end
            begin
              mem_check[50][17].run()  ;
            end
            begin
              rf_driver[50][17].run()  ;
            end

            begin
              gen[50][18].run()  ;
            end
            begin
              drv[50][18].run()  ;
            end
            begin
              mem_check[50][18].run()  ;
            end
            begin
              rf_driver[50][18].run()  ;
            end

            begin
              gen[50][19].run()  ;
            end
            begin
              drv[50][19].run()  ;
            end
            begin
              mem_check[50][19].run()  ;
            end
            begin
              rf_driver[50][19].run()  ;
            end

            begin
              gen[50][20].run()  ;
            end
            begin
              drv[50][20].run()  ;
            end
            begin
              mem_check[50][20].run()  ;
            end
            begin
              rf_driver[50][20].run()  ;
            end

            begin
              gen[50][21].run()  ;
            end
            begin
              drv[50][21].run()  ;
            end
            begin
              mem_check[50][21].run()  ;
            end
            begin
              rf_driver[50][21].run()  ;
            end

            begin
              gen[50][22].run()  ;
            end
            begin
              drv[50][22].run()  ;
            end
            begin
              mem_check[50][22].run()  ;
            end
            begin
              rf_driver[50][22].run()  ;
            end

            begin
              gen[50][23].run()  ;
            end
            begin
              drv[50][23].run()  ;
            end
            begin
              mem_check[50][23].run()  ;
            end
            begin
              rf_driver[50][23].run()  ;
            end

            begin
              gen[50][24].run()  ;
            end
            begin
              drv[50][24].run()  ;
            end
            begin
              mem_check[50][24].run()  ;
            end
            begin
              rf_driver[50][24].run()  ;
            end

            begin
              gen[50][25].run()  ;
            end
            begin
              drv[50][25].run()  ;
            end
            begin
              mem_check[50][25].run()  ;
            end
            begin
              rf_driver[50][25].run()  ;
            end

            begin
              gen[50][26].run()  ;
            end
            begin
              drv[50][26].run()  ;
            end
            begin
              mem_check[50][26].run()  ;
            end
            begin
              rf_driver[50][26].run()  ;
            end

            begin
              gen[50][27].run()  ;
            end
            begin
              drv[50][27].run()  ;
            end
            begin
              mem_check[50][27].run()  ;
            end
            begin
              rf_driver[50][27].run()  ;
            end

            begin
              gen[50][28].run()  ;
            end
            begin
              drv[50][28].run()  ;
            end
            begin
              mem_check[50][28].run()  ;
            end
            begin
              rf_driver[50][28].run()  ;
            end

            begin
              gen[50][29].run()  ;
            end
            begin
              drv[50][29].run()  ;
            end
            begin
              mem_check[50][29].run()  ;
            end
            begin
              rf_driver[50][29].run()  ;
            end

            begin
              gen[50][30].run()  ;
            end
            begin
              drv[50][30].run()  ;
            end
            begin
              mem_check[50][30].run()  ;
            end
            begin
              rf_driver[50][30].run()  ;
            end

            begin
              gen[50][31].run()  ;
            end
            begin
              drv[50][31].run()  ;
            end
            begin
              mem_check[50][31].run()  ;
            end
            begin
              rf_driver[50][31].run()  ;
            end

            begin
              ldst_driver[51].run()  ;
            end
            begin
              mgr[51].run()  ;
            end
            begin
              oob_drv[51].run()  ;
            end
            begin
              up_check[51].run()  ;
            end
            begin
              gen[51][0].run()  ;
            end
            begin
              drv[51][0].run()  ;
            end
            begin
              mem_check[51][0].run()  ;
            end
            begin
              rf_driver[51][0].run()  ;
            end

            begin
              gen[51][1].run()  ;
            end
            begin
              drv[51][1].run()  ;
            end
            begin
              mem_check[51][1].run()  ;
            end
            begin
              rf_driver[51][1].run()  ;
            end

            begin
              gen[51][2].run()  ;
            end
            begin
              drv[51][2].run()  ;
            end
            begin
              mem_check[51][2].run()  ;
            end
            begin
              rf_driver[51][2].run()  ;
            end

            begin
              gen[51][3].run()  ;
            end
            begin
              drv[51][3].run()  ;
            end
            begin
              mem_check[51][3].run()  ;
            end
            begin
              rf_driver[51][3].run()  ;
            end

            begin
              gen[51][4].run()  ;
            end
            begin
              drv[51][4].run()  ;
            end
            begin
              mem_check[51][4].run()  ;
            end
            begin
              rf_driver[51][4].run()  ;
            end

            begin
              gen[51][5].run()  ;
            end
            begin
              drv[51][5].run()  ;
            end
            begin
              mem_check[51][5].run()  ;
            end
            begin
              rf_driver[51][5].run()  ;
            end

            begin
              gen[51][6].run()  ;
            end
            begin
              drv[51][6].run()  ;
            end
            begin
              mem_check[51][6].run()  ;
            end
            begin
              rf_driver[51][6].run()  ;
            end

            begin
              gen[51][7].run()  ;
            end
            begin
              drv[51][7].run()  ;
            end
            begin
              mem_check[51][7].run()  ;
            end
            begin
              rf_driver[51][7].run()  ;
            end

            begin
              gen[51][8].run()  ;
            end
            begin
              drv[51][8].run()  ;
            end
            begin
              mem_check[51][8].run()  ;
            end
            begin
              rf_driver[51][8].run()  ;
            end

            begin
              gen[51][9].run()  ;
            end
            begin
              drv[51][9].run()  ;
            end
            begin
              mem_check[51][9].run()  ;
            end
            begin
              rf_driver[51][9].run()  ;
            end

            begin
              gen[51][10].run()  ;
            end
            begin
              drv[51][10].run()  ;
            end
            begin
              mem_check[51][10].run()  ;
            end
            begin
              rf_driver[51][10].run()  ;
            end

            begin
              gen[51][11].run()  ;
            end
            begin
              drv[51][11].run()  ;
            end
            begin
              mem_check[51][11].run()  ;
            end
            begin
              rf_driver[51][11].run()  ;
            end

            begin
              gen[51][12].run()  ;
            end
            begin
              drv[51][12].run()  ;
            end
            begin
              mem_check[51][12].run()  ;
            end
            begin
              rf_driver[51][12].run()  ;
            end

            begin
              gen[51][13].run()  ;
            end
            begin
              drv[51][13].run()  ;
            end
            begin
              mem_check[51][13].run()  ;
            end
            begin
              rf_driver[51][13].run()  ;
            end

            begin
              gen[51][14].run()  ;
            end
            begin
              drv[51][14].run()  ;
            end
            begin
              mem_check[51][14].run()  ;
            end
            begin
              rf_driver[51][14].run()  ;
            end

            begin
              gen[51][15].run()  ;
            end
            begin
              drv[51][15].run()  ;
            end
            begin
              mem_check[51][15].run()  ;
            end
            begin
              rf_driver[51][15].run()  ;
            end

            begin
              gen[51][16].run()  ;
            end
            begin
              drv[51][16].run()  ;
            end
            begin
              mem_check[51][16].run()  ;
            end
            begin
              rf_driver[51][16].run()  ;
            end

            begin
              gen[51][17].run()  ;
            end
            begin
              drv[51][17].run()  ;
            end
            begin
              mem_check[51][17].run()  ;
            end
            begin
              rf_driver[51][17].run()  ;
            end

            begin
              gen[51][18].run()  ;
            end
            begin
              drv[51][18].run()  ;
            end
            begin
              mem_check[51][18].run()  ;
            end
            begin
              rf_driver[51][18].run()  ;
            end

            begin
              gen[51][19].run()  ;
            end
            begin
              drv[51][19].run()  ;
            end
            begin
              mem_check[51][19].run()  ;
            end
            begin
              rf_driver[51][19].run()  ;
            end

            begin
              gen[51][20].run()  ;
            end
            begin
              drv[51][20].run()  ;
            end
            begin
              mem_check[51][20].run()  ;
            end
            begin
              rf_driver[51][20].run()  ;
            end

            begin
              gen[51][21].run()  ;
            end
            begin
              drv[51][21].run()  ;
            end
            begin
              mem_check[51][21].run()  ;
            end
            begin
              rf_driver[51][21].run()  ;
            end

            begin
              gen[51][22].run()  ;
            end
            begin
              drv[51][22].run()  ;
            end
            begin
              mem_check[51][22].run()  ;
            end
            begin
              rf_driver[51][22].run()  ;
            end

            begin
              gen[51][23].run()  ;
            end
            begin
              drv[51][23].run()  ;
            end
            begin
              mem_check[51][23].run()  ;
            end
            begin
              rf_driver[51][23].run()  ;
            end

            begin
              gen[51][24].run()  ;
            end
            begin
              drv[51][24].run()  ;
            end
            begin
              mem_check[51][24].run()  ;
            end
            begin
              rf_driver[51][24].run()  ;
            end

            begin
              gen[51][25].run()  ;
            end
            begin
              drv[51][25].run()  ;
            end
            begin
              mem_check[51][25].run()  ;
            end
            begin
              rf_driver[51][25].run()  ;
            end

            begin
              gen[51][26].run()  ;
            end
            begin
              drv[51][26].run()  ;
            end
            begin
              mem_check[51][26].run()  ;
            end
            begin
              rf_driver[51][26].run()  ;
            end

            begin
              gen[51][27].run()  ;
            end
            begin
              drv[51][27].run()  ;
            end
            begin
              mem_check[51][27].run()  ;
            end
            begin
              rf_driver[51][27].run()  ;
            end

            begin
              gen[51][28].run()  ;
            end
            begin
              drv[51][28].run()  ;
            end
            begin
              mem_check[51][28].run()  ;
            end
            begin
              rf_driver[51][28].run()  ;
            end

            begin
              gen[51][29].run()  ;
            end
            begin
              drv[51][29].run()  ;
            end
            begin
              mem_check[51][29].run()  ;
            end
            begin
              rf_driver[51][29].run()  ;
            end

            begin
              gen[51][30].run()  ;
            end
            begin
              drv[51][30].run()  ;
            end
            begin
              mem_check[51][30].run()  ;
            end
            begin
              rf_driver[51][30].run()  ;
            end

            begin
              gen[51][31].run()  ;
            end
            begin
              drv[51][31].run()  ;
            end
            begin
              mem_check[51][31].run()  ;
            end
            begin
              rf_driver[51][31].run()  ;
            end

            begin
              ldst_driver[52].run()  ;
            end
            begin
              mgr[52].run()  ;
            end
            begin
              oob_drv[52].run()  ;
            end
            begin
              up_check[52].run()  ;
            end
            begin
              gen[52][0].run()  ;
            end
            begin
              drv[52][0].run()  ;
            end
            begin
              mem_check[52][0].run()  ;
            end
            begin
              rf_driver[52][0].run()  ;
            end

            begin
              gen[52][1].run()  ;
            end
            begin
              drv[52][1].run()  ;
            end
            begin
              mem_check[52][1].run()  ;
            end
            begin
              rf_driver[52][1].run()  ;
            end

            begin
              gen[52][2].run()  ;
            end
            begin
              drv[52][2].run()  ;
            end
            begin
              mem_check[52][2].run()  ;
            end
            begin
              rf_driver[52][2].run()  ;
            end

            begin
              gen[52][3].run()  ;
            end
            begin
              drv[52][3].run()  ;
            end
            begin
              mem_check[52][3].run()  ;
            end
            begin
              rf_driver[52][3].run()  ;
            end

            begin
              gen[52][4].run()  ;
            end
            begin
              drv[52][4].run()  ;
            end
            begin
              mem_check[52][4].run()  ;
            end
            begin
              rf_driver[52][4].run()  ;
            end

            begin
              gen[52][5].run()  ;
            end
            begin
              drv[52][5].run()  ;
            end
            begin
              mem_check[52][5].run()  ;
            end
            begin
              rf_driver[52][5].run()  ;
            end

            begin
              gen[52][6].run()  ;
            end
            begin
              drv[52][6].run()  ;
            end
            begin
              mem_check[52][6].run()  ;
            end
            begin
              rf_driver[52][6].run()  ;
            end

            begin
              gen[52][7].run()  ;
            end
            begin
              drv[52][7].run()  ;
            end
            begin
              mem_check[52][7].run()  ;
            end
            begin
              rf_driver[52][7].run()  ;
            end

            begin
              gen[52][8].run()  ;
            end
            begin
              drv[52][8].run()  ;
            end
            begin
              mem_check[52][8].run()  ;
            end
            begin
              rf_driver[52][8].run()  ;
            end

            begin
              gen[52][9].run()  ;
            end
            begin
              drv[52][9].run()  ;
            end
            begin
              mem_check[52][9].run()  ;
            end
            begin
              rf_driver[52][9].run()  ;
            end

            begin
              gen[52][10].run()  ;
            end
            begin
              drv[52][10].run()  ;
            end
            begin
              mem_check[52][10].run()  ;
            end
            begin
              rf_driver[52][10].run()  ;
            end

            begin
              gen[52][11].run()  ;
            end
            begin
              drv[52][11].run()  ;
            end
            begin
              mem_check[52][11].run()  ;
            end
            begin
              rf_driver[52][11].run()  ;
            end

            begin
              gen[52][12].run()  ;
            end
            begin
              drv[52][12].run()  ;
            end
            begin
              mem_check[52][12].run()  ;
            end
            begin
              rf_driver[52][12].run()  ;
            end

            begin
              gen[52][13].run()  ;
            end
            begin
              drv[52][13].run()  ;
            end
            begin
              mem_check[52][13].run()  ;
            end
            begin
              rf_driver[52][13].run()  ;
            end

            begin
              gen[52][14].run()  ;
            end
            begin
              drv[52][14].run()  ;
            end
            begin
              mem_check[52][14].run()  ;
            end
            begin
              rf_driver[52][14].run()  ;
            end

            begin
              gen[52][15].run()  ;
            end
            begin
              drv[52][15].run()  ;
            end
            begin
              mem_check[52][15].run()  ;
            end
            begin
              rf_driver[52][15].run()  ;
            end

            begin
              gen[52][16].run()  ;
            end
            begin
              drv[52][16].run()  ;
            end
            begin
              mem_check[52][16].run()  ;
            end
            begin
              rf_driver[52][16].run()  ;
            end

            begin
              gen[52][17].run()  ;
            end
            begin
              drv[52][17].run()  ;
            end
            begin
              mem_check[52][17].run()  ;
            end
            begin
              rf_driver[52][17].run()  ;
            end

            begin
              gen[52][18].run()  ;
            end
            begin
              drv[52][18].run()  ;
            end
            begin
              mem_check[52][18].run()  ;
            end
            begin
              rf_driver[52][18].run()  ;
            end

            begin
              gen[52][19].run()  ;
            end
            begin
              drv[52][19].run()  ;
            end
            begin
              mem_check[52][19].run()  ;
            end
            begin
              rf_driver[52][19].run()  ;
            end

            begin
              gen[52][20].run()  ;
            end
            begin
              drv[52][20].run()  ;
            end
            begin
              mem_check[52][20].run()  ;
            end
            begin
              rf_driver[52][20].run()  ;
            end

            begin
              gen[52][21].run()  ;
            end
            begin
              drv[52][21].run()  ;
            end
            begin
              mem_check[52][21].run()  ;
            end
            begin
              rf_driver[52][21].run()  ;
            end

            begin
              gen[52][22].run()  ;
            end
            begin
              drv[52][22].run()  ;
            end
            begin
              mem_check[52][22].run()  ;
            end
            begin
              rf_driver[52][22].run()  ;
            end

            begin
              gen[52][23].run()  ;
            end
            begin
              drv[52][23].run()  ;
            end
            begin
              mem_check[52][23].run()  ;
            end
            begin
              rf_driver[52][23].run()  ;
            end

            begin
              gen[52][24].run()  ;
            end
            begin
              drv[52][24].run()  ;
            end
            begin
              mem_check[52][24].run()  ;
            end
            begin
              rf_driver[52][24].run()  ;
            end

            begin
              gen[52][25].run()  ;
            end
            begin
              drv[52][25].run()  ;
            end
            begin
              mem_check[52][25].run()  ;
            end
            begin
              rf_driver[52][25].run()  ;
            end

            begin
              gen[52][26].run()  ;
            end
            begin
              drv[52][26].run()  ;
            end
            begin
              mem_check[52][26].run()  ;
            end
            begin
              rf_driver[52][26].run()  ;
            end

            begin
              gen[52][27].run()  ;
            end
            begin
              drv[52][27].run()  ;
            end
            begin
              mem_check[52][27].run()  ;
            end
            begin
              rf_driver[52][27].run()  ;
            end

            begin
              gen[52][28].run()  ;
            end
            begin
              drv[52][28].run()  ;
            end
            begin
              mem_check[52][28].run()  ;
            end
            begin
              rf_driver[52][28].run()  ;
            end

            begin
              gen[52][29].run()  ;
            end
            begin
              drv[52][29].run()  ;
            end
            begin
              mem_check[52][29].run()  ;
            end
            begin
              rf_driver[52][29].run()  ;
            end

            begin
              gen[52][30].run()  ;
            end
            begin
              drv[52][30].run()  ;
            end
            begin
              mem_check[52][30].run()  ;
            end
            begin
              rf_driver[52][30].run()  ;
            end

            begin
              gen[52][31].run()  ;
            end
            begin
              drv[52][31].run()  ;
            end
            begin
              mem_check[52][31].run()  ;
            end
            begin
              rf_driver[52][31].run()  ;
            end

            begin
              ldst_driver[53].run()  ;
            end
            begin
              mgr[53].run()  ;
            end
            begin
              oob_drv[53].run()  ;
            end
            begin
              up_check[53].run()  ;
            end
            begin
              gen[53][0].run()  ;
            end
            begin
              drv[53][0].run()  ;
            end
            begin
              mem_check[53][0].run()  ;
            end
            begin
              rf_driver[53][0].run()  ;
            end

            begin
              gen[53][1].run()  ;
            end
            begin
              drv[53][1].run()  ;
            end
            begin
              mem_check[53][1].run()  ;
            end
            begin
              rf_driver[53][1].run()  ;
            end

            begin
              gen[53][2].run()  ;
            end
            begin
              drv[53][2].run()  ;
            end
            begin
              mem_check[53][2].run()  ;
            end
            begin
              rf_driver[53][2].run()  ;
            end

            begin
              gen[53][3].run()  ;
            end
            begin
              drv[53][3].run()  ;
            end
            begin
              mem_check[53][3].run()  ;
            end
            begin
              rf_driver[53][3].run()  ;
            end

            begin
              gen[53][4].run()  ;
            end
            begin
              drv[53][4].run()  ;
            end
            begin
              mem_check[53][4].run()  ;
            end
            begin
              rf_driver[53][4].run()  ;
            end

            begin
              gen[53][5].run()  ;
            end
            begin
              drv[53][5].run()  ;
            end
            begin
              mem_check[53][5].run()  ;
            end
            begin
              rf_driver[53][5].run()  ;
            end

            begin
              gen[53][6].run()  ;
            end
            begin
              drv[53][6].run()  ;
            end
            begin
              mem_check[53][6].run()  ;
            end
            begin
              rf_driver[53][6].run()  ;
            end

            begin
              gen[53][7].run()  ;
            end
            begin
              drv[53][7].run()  ;
            end
            begin
              mem_check[53][7].run()  ;
            end
            begin
              rf_driver[53][7].run()  ;
            end

            begin
              gen[53][8].run()  ;
            end
            begin
              drv[53][8].run()  ;
            end
            begin
              mem_check[53][8].run()  ;
            end
            begin
              rf_driver[53][8].run()  ;
            end

            begin
              gen[53][9].run()  ;
            end
            begin
              drv[53][9].run()  ;
            end
            begin
              mem_check[53][9].run()  ;
            end
            begin
              rf_driver[53][9].run()  ;
            end

            begin
              gen[53][10].run()  ;
            end
            begin
              drv[53][10].run()  ;
            end
            begin
              mem_check[53][10].run()  ;
            end
            begin
              rf_driver[53][10].run()  ;
            end

            begin
              gen[53][11].run()  ;
            end
            begin
              drv[53][11].run()  ;
            end
            begin
              mem_check[53][11].run()  ;
            end
            begin
              rf_driver[53][11].run()  ;
            end

            begin
              gen[53][12].run()  ;
            end
            begin
              drv[53][12].run()  ;
            end
            begin
              mem_check[53][12].run()  ;
            end
            begin
              rf_driver[53][12].run()  ;
            end

            begin
              gen[53][13].run()  ;
            end
            begin
              drv[53][13].run()  ;
            end
            begin
              mem_check[53][13].run()  ;
            end
            begin
              rf_driver[53][13].run()  ;
            end

            begin
              gen[53][14].run()  ;
            end
            begin
              drv[53][14].run()  ;
            end
            begin
              mem_check[53][14].run()  ;
            end
            begin
              rf_driver[53][14].run()  ;
            end

            begin
              gen[53][15].run()  ;
            end
            begin
              drv[53][15].run()  ;
            end
            begin
              mem_check[53][15].run()  ;
            end
            begin
              rf_driver[53][15].run()  ;
            end

            begin
              gen[53][16].run()  ;
            end
            begin
              drv[53][16].run()  ;
            end
            begin
              mem_check[53][16].run()  ;
            end
            begin
              rf_driver[53][16].run()  ;
            end

            begin
              gen[53][17].run()  ;
            end
            begin
              drv[53][17].run()  ;
            end
            begin
              mem_check[53][17].run()  ;
            end
            begin
              rf_driver[53][17].run()  ;
            end

            begin
              gen[53][18].run()  ;
            end
            begin
              drv[53][18].run()  ;
            end
            begin
              mem_check[53][18].run()  ;
            end
            begin
              rf_driver[53][18].run()  ;
            end

            begin
              gen[53][19].run()  ;
            end
            begin
              drv[53][19].run()  ;
            end
            begin
              mem_check[53][19].run()  ;
            end
            begin
              rf_driver[53][19].run()  ;
            end

            begin
              gen[53][20].run()  ;
            end
            begin
              drv[53][20].run()  ;
            end
            begin
              mem_check[53][20].run()  ;
            end
            begin
              rf_driver[53][20].run()  ;
            end

            begin
              gen[53][21].run()  ;
            end
            begin
              drv[53][21].run()  ;
            end
            begin
              mem_check[53][21].run()  ;
            end
            begin
              rf_driver[53][21].run()  ;
            end

            begin
              gen[53][22].run()  ;
            end
            begin
              drv[53][22].run()  ;
            end
            begin
              mem_check[53][22].run()  ;
            end
            begin
              rf_driver[53][22].run()  ;
            end

            begin
              gen[53][23].run()  ;
            end
            begin
              drv[53][23].run()  ;
            end
            begin
              mem_check[53][23].run()  ;
            end
            begin
              rf_driver[53][23].run()  ;
            end

            begin
              gen[53][24].run()  ;
            end
            begin
              drv[53][24].run()  ;
            end
            begin
              mem_check[53][24].run()  ;
            end
            begin
              rf_driver[53][24].run()  ;
            end

            begin
              gen[53][25].run()  ;
            end
            begin
              drv[53][25].run()  ;
            end
            begin
              mem_check[53][25].run()  ;
            end
            begin
              rf_driver[53][25].run()  ;
            end

            begin
              gen[53][26].run()  ;
            end
            begin
              drv[53][26].run()  ;
            end
            begin
              mem_check[53][26].run()  ;
            end
            begin
              rf_driver[53][26].run()  ;
            end

            begin
              gen[53][27].run()  ;
            end
            begin
              drv[53][27].run()  ;
            end
            begin
              mem_check[53][27].run()  ;
            end
            begin
              rf_driver[53][27].run()  ;
            end

            begin
              gen[53][28].run()  ;
            end
            begin
              drv[53][28].run()  ;
            end
            begin
              mem_check[53][28].run()  ;
            end
            begin
              rf_driver[53][28].run()  ;
            end

            begin
              gen[53][29].run()  ;
            end
            begin
              drv[53][29].run()  ;
            end
            begin
              mem_check[53][29].run()  ;
            end
            begin
              rf_driver[53][29].run()  ;
            end

            begin
              gen[53][30].run()  ;
            end
            begin
              drv[53][30].run()  ;
            end
            begin
              mem_check[53][30].run()  ;
            end
            begin
              rf_driver[53][30].run()  ;
            end

            begin
              gen[53][31].run()  ;
            end
            begin
              drv[53][31].run()  ;
            end
            begin
              mem_check[53][31].run()  ;
            end
            begin
              rf_driver[53][31].run()  ;
            end

            begin
              ldst_driver[54].run()  ;
            end
            begin
              mgr[54].run()  ;
            end
            begin
              oob_drv[54].run()  ;
            end
            begin
              up_check[54].run()  ;
            end
            begin
              gen[54][0].run()  ;
            end
            begin
              drv[54][0].run()  ;
            end
            begin
              mem_check[54][0].run()  ;
            end
            begin
              rf_driver[54][0].run()  ;
            end

            begin
              gen[54][1].run()  ;
            end
            begin
              drv[54][1].run()  ;
            end
            begin
              mem_check[54][1].run()  ;
            end
            begin
              rf_driver[54][1].run()  ;
            end

            begin
              gen[54][2].run()  ;
            end
            begin
              drv[54][2].run()  ;
            end
            begin
              mem_check[54][2].run()  ;
            end
            begin
              rf_driver[54][2].run()  ;
            end

            begin
              gen[54][3].run()  ;
            end
            begin
              drv[54][3].run()  ;
            end
            begin
              mem_check[54][3].run()  ;
            end
            begin
              rf_driver[54][3].run()  ;
            end

            begin
              gen[54][4].run()  ;
            end
            begin
              drv[54][4].run()  ;
            end
            begin
              mem_check[54][4].run()  ;
            end
            begin
              rf_driver[54][4].run()  ;
            end

            begin
              gen[54][5].run()  ;
            end
            begin
              drv[54][5].run()  ;
            end
            begin
              mem_check[54][5].run()  ;
            end
            begin
              rf_driver[54][5].run()  ;
            end

            begin
              gen[54][6].run()  ;
            end
            begin
              drv[54][6].run()  ;
            end
            begin
              mem_check[54][6].run()  ;
            end
            begin
              rf_driver[54][6].run()  ;
            end

            begin
              gen[54][7].run()  ;
            end
            begin
              drv[54][7].run()  ;
            end
            begin
              mem_check[54][7].run()  ;
            end
            begin
              rf_driver[54][7].run()  ;
            end

            begin
              gen[54][8].run()  ;
            end
            begin
              drv[54][8].run()  ;
            end
            begin
              mem_check[54][8].run()  ;
            end
            begin
              rf_driver[54][8].run()  ;
            end

            begin
              gen[54][9].run()  ;
            end
            begin
              drv[54][9].run()  ;
            end
            begin
              mem_check[54][9].run()  ;
            end
            begin
              rf_driver[54][9].run()  ;
            end

            begin
              gen[54][10].run()  ;
            end
            begin
              drv[54][10].run()  ;
            end
            begin
              mem_check[54][10].run()  ;
            end
            begin
              rf_driver[54][10].run()  ;
            end

            begin
              gen[54][11].run()  ;
            end
            begin
              drv[54][11].run()  ;
            end
            begin
              mem_check[54][11].run()  ;
            end
            begin
              rf_driver[54][11].run()  ;
            end

            begin
              gen[54][12].run()  ;
            end
            begin
              drv[54][12].run()  ;
            end
            begin
              mem_check[54][12].run()  ;
            end
            begin
              rf_driver[54][12].run()  ;
            end

            begin
              gen[54][13].run()  ;
            end
            begin
              drv[54][13].run()  ;
            end
            begin
              mem_check[54][13].run()  ;
            end
            begin
              rf_driver[54][13].run()  ;
            end

            begin
              gen[54][14].run()  ;
            end
            begin
              drv[54][14].run()  ;
            end
            begin
              mem_check[54][14].run()  ;
            end
            begin
              rf_driver[54][14].run()  ;
            end

            begin
              gen[54][15].run()  ;
            end
            begin
              drv[54][15].run()  ;
            end
            begin
              mem_check[54][15].run()  ;
            end
            begin
              rf_driver[54][15].run()  ;
            end

            begin
              gen[54][16].run()  ;
            end
            begin
              drv[54][16].run()  ;
            end
            begin
              mem_check[54][16].run()  ;
            end
            begin
              rf_driver[54][16].run()  ;
            end

            begin
              gen[54][17].run()  ;
            end
            begin
              drv[54][17].run()  ;
            end
            begin
              mem_check[54][17].run()  ;
            end
            begin
              rf_driver[54][17].run()  ;
            end

            begin
              gen[54][18].run()  ;
            end
            begin
              drv[54][18].run()  ;
            end
            begin
              mem_check[54][18].run()  ;
            end
            begin
              rf_driver[54][18].run()  ;
            end

            begin
              gen[54][19].run()  ;
            end
            begin
              drv[54][19].run()  ;
            end
            begin
              mem_check[54][19].run()  ;
            end
            begin
              rf_driver[54][19].run()  ;
            end

            begin
              gen[54][20].run()  ;
            end
            begin
              drv[54][20].run()  ;
            end
            begin
              mem_check[54][20].run()  ;
            end
            begin
              rf_driver[54][20].run()  ;
            end

            begin
              gen[54][21].run()  ;
            end
            begin
              drv[54][21].run()  ;
            end
            begin
              mem_check[54][21].run()  ;
            end
            begin
              rf_driver[54][21].run()  ;
            end

            begin
              gen[54][22].run()  ;
            end
            begin
              drv[54][22].run()  ;
            end
            begin
              mem_check[54][22].run()  ;
            end
            begin
              rf_driver[54][22].run()  ;
            end

            begin
              gen[54][23].run()  ;
            end
            begin
              drv[54][23].run()  ;
            end
            begin
              mem_check[54][23].run()  ;
            end
            begin
              rf_driver[54][23].run()  ;
            end

            begin
              gen[54][24].run()  ;
            end
            begin
              drv[54][24].run()  ;
            end
            begin
              mem_check[54][24].run()  ;
            end
            begin
              rf_driver[54][24].run()  ;
            end

            begin
              gen[54][25].run()  ;
            end
            begin
              drv[54][25].run()  ;
            end
            begin
              mem_check[54][25].run()  ;
            end
            begin
              rf_driver[54][25].run()  ;
            end

            begin
              gen[54][26].run()  ;
            end
            begin
              drv[54][26].run()  ;
            end
            begin
              mem_check[54][26].run()  ;
            end
            begin
              rf_driver[54][26].run()  ;
            end

            begin
              gen[54][27].run()  ;
            end
            begin
              drv[54][27].run()  ;
            end
            begin
              mem_check[54][27].run()  ;
            end
            begin
              rf_driver[54][27].run()  ;
            end

            begin
              gen[54][28].run()  ;
            end
            begin
              drv[54][28].run()  ;
            end
            begin
              mem_check[54][28].run()  ;
            end
            begin
              rf_driver[54][28].run()  ;
            end

            begin
              gen[54][29].run()  ;
            end
            begin
              drv[54][29].run()  ;
            end
            begin
              mem_check[54][29].run()  ;
            end
            begin
              rf_driver[54][29].run()  ;
            end

            begin
              gen[54][30].run()  ;
            end
            begin
              drv[54][30].run()  ;
            end
            begin
              mem_check[54][30].run()  ;
            end
            begin
              rf_driver[54][30].run()  ;
            end

            begin
              gen[54][31].run()  ;
            end
            begin
              drv[54][31].run()  ;
            end
            begin
              mem_check[54][31].run()  ;
            end
            begin
              rf_driver[54][31].run()  ;
            end

            begin
              ldst_driver[55].run()  ;
            end
            begin
              mgr[55].run()  ;
            end
            begin
              oob_drv[55].run()  ;
            end
            begin
              up_check[55].run()  ;
            end
            begin
              gen[55][0].run()  ;
            end
            begin
              drv[55][0].run()  ;
            end
            begin
              mem_check[55][0].run()  ;
            end
            begin
              rf_driver[55][0].run()  ;
            end

            begin
              gen[55][1].run()  ;
            end
            begin
              drv[55][1].run()  ;
            end
            begin
              mem_check[55][1].run()  ;
            end
            begin
              rf_driver[55][1].run()  ;
            end

            begin
              gen[55][2].run()  ;
            end
            begin
              drv[55][2].run()  ;
            end
            begin
              mem_check[55][2].run()  ;
            end
            begin
              rf_driver[55][2].run()  ;
            end

            begin
              gen[55][3].run()  ;
            end
            begin
              drv[55][3].run()  ;
            end
            begin
              mem_check[55][3].run()  ;
            end
            begin
              rf_driver[55][3].run()  ;
            end

            begin
              gen[55][4].run()  ;
            end
            begin
              drv[55][4].run()  ;
            end
            begin
              mem_check[55][4].run()  ;
            end
            begin
              rf_driver[55][4].run()  ;
            end

            begin
              gen[55][5].run()  ;
            end
            begin
              drv[55][5].run()  ;
            end
            begin
              mem_check[55][5].run()  ;
            end
            begin
              rf_driver[55][5].run()  ;
            end

            begin
              gen[55][6].run()  ;
            end
            begin
              drv[55][6].run()  ;
            end
            begin
              mem_check[55][6].run()  ;
            end
            begin
              rf_driver[55][6].run()  ;
            end

            begin
              gen[55][7].run()  ;
            end
            begin
              drv[55][7].run()  ;
            end
            begin
              mem_check[55][7].run()  ;
            end
            begin
              rf_driver[55][7].run()  ;
            end

            begin
              gen[55][8].run()  ;
            end
            begin
              drv[55][8].run()  ;
            end
            begin
              mem_check[55][8].run()  ;
            end
            begin
              rf_driver[55][8].run()  ;
            end

            begin
              gen[55][9].run()  ;
            end
            begin
              drv[55][9].run()  ;
            end
            begin
              mem_check[55][9].run()  ;
            end
            begin
              rf_driver[55][9].run()  ;
            end

            begin
              gen[55][10].run()  ;
            end
            begin
              drv[55][10].run()  ;
            end
            begin
              mem_check[55][10].run()  ;
            end
            begin
              rf_driver[55][10].run()  ;
            end

            begin
              gen[55][11].run()  ;
            end
            begin
              drv[55][11].run()  ;
            end
            begin
              mem_check[55][11].run()  ;
            end
            begin
              rf_driver[55][11].run()  ;
            end

            begin
              gen[55][12].run()  ;
            end
            begin
              drv[55][12].run()  ;
            end
            begin
              mem_check[55][12].run()  ;
            end
            begin
              rf_driver[55][12].run()  ;
            end

            begin
              gen[55][13].run()  ;
            end
            begin
              drv[55][13].run()  ;
            end
            begin
              mem_check[55][13].run()  ;
            end
            begin
              rf_driver[55][13].run()  ;
            end

            begin
              gen[55][14].run()  ;
            end
            begin
              drv[55][14].run()  ;
            end
            begin
              mem_check[55][14].run()  ;
            end
            begin
              rf_driver[55][14].run()  ;
            end

            begin
              gen[55][15].run()  ;
            end
            begin
              drv[55][15].run()  ;
            end
            begin
              mem_check[55][15].run()  ;
            end
            begin
              rf_driver[55][15].run()  ;
            end

            begin
              gen[55][16].run()  ;
            end
            begin
              drv[55][16].run()  ;
            end
            begin
              mem_check[55][16].run()  ;
            end
            begin
              rf_driver[55][16].run()  ;
            end

            begin
              gen[55][17].run()  ;
            end
            begin
              drv[55][17].run()  ;
            end
            begin
              mem_check[55][17].run()  ;
            end
            begin
              rf_driver[55][17].run()  ;
            end

            begin
              gen[55][18].run()  ;
            end
            begin
              drv[55][18].run()  ;
            end
            begin
              mem_check[55][18].run()  ;
            end
            begin
              rf_driver[55][18].run()  ;
            end

            begin
              gen[55][19].run()  ;
            end
            begin
              drv[55][19].run()  ;
            end
            begin
              mem_check[55][19].run()  ;
            end
            begin
              rf_driver[55][19].run()  ;
            end

            begin
              gen[55][20].run()  ;
            end
            begin
              drv[55][20].run()  ;
            end
            begin
              mem_check[55][20].run()  ;
            end
            begin
              rf_driver[55][20].run()  ;
            end

            begin
              gen[55][21].run()  ;
            end
            begin
              drv[55][21].run()  ;
            end
            begin
              mem_check[55][21].run()  ;
            end
            begin
              rf_driver[55][21].run()  ;
            end

            begin
              gen[55][22].run()  ;
            end
            begin
              drv[55][22].run()  ;
            end
            begin
              mem_check[55][22].run()  ;
            end
            begin
              rf_driver[55][22].run()  ;
            end

            begin
              gen[55][23].run()  ;
            end
            begin
              drv[55][23].run()  ;
            end
            begin
              mem_check[55][23].run()  ;
            end
            begin
              rf_driver[55][23].run()  ;
            end

            begin
              gen[55][24].run()  ;
            end
            begin
              drv[55][24].run()  ;
            end
            begin
              mem_check[55][24].run()  ;
            end
            begin
              rf_driver[55][24].run()  ;
            end

            begin
              gen[55][25].run()  ;
            end
            begin
              drv[55][25].run()  ;
            end
            begin
              mem_check[55][25].run()  ;
            end
            begin
              rf_driver[55][25].run()  ;
            end

            begin
              gen[55][26].run()  ;
            end
            begin
              drv[55][26].run()  ;
            end
            begin
              mem_check[55][26].run()  ;
            end
            begin
              rf_driver[55][26].run()  ;
            end

            begin
              gen[55][27].run()  ;
            end
            begin
              drv[55][27].run()  ;
            end
            begin
              mem_check[55][27].run()  ;
            end
            begin
              rf_driver[55][27].run()  ;
            end

            begin
              gen[55][28].run()  ;
            end
            begin
              drv[55][28].run()  ;
            end
            begin
              mem_check[55][28].run()  ;
            end
            begin
              rf_driver[55][28].run()  ;
            end

            begin
              gen[55][29].run()  ;
            end
            begin
              drv[55][29].run()  ;
            end
            begin
              mem_check[55][29].run()  ;
            end
            begin
              rf_driver[55][29].run()  ;
            end

            begin
              gen[55][30].run()  ;
            end
            begin
              drv[55][30].run()  ;
            end
            begin
              mem_check[55][30].run()  ;
            end
            begin
              rf_driver[55][30].run()  ;
            end

            begin
              gen[55][31].run()  ;
            end
            begin
              drv[55][31].run()  ;
            end
            begin
              mem_check[55][31].run()  ;
            end
            begin
              rf_driver[55][31].run()  ;
            end

            begin
              ldst_driver[56].run()  ;
            end
            begin
              mgr[56].run()  ;
            end
            begin
              oob_drv[56].run()  ;
            end
            begin
              up_check[56].run()  ;
            end
            begin
              gen[56][0].run()  ;
            end
            begin
              drv[56][0].run()  ;
            end
            begin
              mem_check[56][0].run()  ;
            end
            begin
              rf_driver[56][0].run()  ;
            end

            begin
              gen[56][1].run()  ;
            end
            begin
              drv[56][1].run()  ;
            end
            begin
              mem_check[56][1].run()  ;
            end
            begin
              rf_driver[56][1].run()  ;
            end

            begin
              gen[56][2].run()  ;
            end
            begin
              drv[56][2].run()  ;
            end
            begin
              mem_check[56][2].run()  ;
            end
            begin
              rf_driver[56][2].run()  ;
            end

            begin
              gen[56][3].run()  ;
            end
            begin
              drv[56][3].run()  ;
            end
            begin
              mem_check[56][3].run()  ;
            end
            begin
              rf_driver[56][3].run()  ;
            end

            begin
              gen[56][4].run()  ;
            end
            begin
              drv[56][4].run()  ;
            end
            begin
              mem_check[56][4].run()  ;
            end
            begin
              rf_driver[56][4].run()  ;
            end

            begin
              gen[56][5].run()  ;
            end
            begin
              drv[56][5].run()  ;
            end
            begin
              mem_check[56][5].run()  ;
            end
            begin
              rf_driver[56][5].run()  ;
            end

            begin
              gen[56][6].run()  ;
            end
            begin
              drv[56][6].run()  ;
            end
            begin
              mem_check[56][6].run()  ;
            end
            begin
              rf_driver[56][6].run()  ;
            end

            begin
              gen[56][7].run()  ;
            end
            begin
              drv[56][7].run()  ;
            end
            begin
              mem_check[56][7].run()  ;
            end
            begin
              rf_driver[56][7].run()  ;
            end

            begin
              gen[56][8].run()  ;
            end
            begin
              drv[56][8].run()  ;
            end
            begin
              mem_check[56][8].run()  ;
            end
            begin
              rf_driver[56][8].run()  ;
            end

            begin
              gen[56][9].run()  ;
            end
            begin
              drv[56][9].run()  ;
            end
            begin
              mem_check[56][9].run()  ;
            end
            begin
              rf_driver[56][9].run()  ;
            end

            begin
              gen[56][10].run()  ;
            end
            begin
              drv[56][10].run()  ;
            end
            begin
              mem_check[56][10].run()  ;
            end
            begin
              rf_driver[56][10].run()  ;
            end

            begin
              gen[56][11].run()  ;
            end
            begin
              drv[56][11].run()  ;
            end
            begin
              mem_check[56][11].run()  ;
            end
            begin
              rf_driver[56][11].run()  ;
            end

            begin
              gen[56][12].run()  ;
            end
            begin
              drv[56][12].run()  ;
            end
            begin
              mem_check[56][12].run()  ;
            end
            begin
              rf_driver[56][12].run()  ;
            end

            begin
              gen[56][13].run()  ;
            end
            begin
              drv[56][13].run()  ;
            end
            begin
              mem_check[56][13].run()  ;
            end
            begin
              rf_driver[56][13].run()  ;
            end

            begin
              gen[56][14].run()  ;
            end
            begin
              drv[56][14].run()  ;
            end
            begin
              mem_check[56][14].run()  ;
            end
            begin
              rf_driver[56][14].run()  ;
            end

            begin
              gen[56][15].run()  ;
            end
            begin
              drv[56][15].run()  ;
            end
            begin
              mem_check[56][15].run()  ;
            end
            begin
              rf_driver[56][15].run()  ;
            end

            begin
              gen[56][16].run()  ;
            end
            begin
              drv[56][16].run()  ;
            end
            begin
              mem_check[56][16].run()  ;
            end
            begin
              rf_driver[56][16].run()  ;
            end

            begin
              gen[56][17].run()  ;
            end
            begin
              drv[56][17].run()  ;
            end
            begin
              mem_check[56][17].run()  ;
            end
            begin
              rf_driver[56][17].run()  ;
            end

            begin
              gen[56][18].run()  ;
            end
            begin
              drv[56][18].run()  ;
            end
            begin
              mem_check[56][18].run()  ;
            end
            begin
              rf_driver[56][18].run()  ;
            end

            begin
              gen[56][19].run()  ;
            end
            begin
              drv[56][19].run()  ;
            end
            begin
              mem_check[56][19].run()  ;
            end
            begin
              rf_driver[56][19].run()  ;
            end

            begin
              gen[56][20].run()  ;
            end
            begin
              drv[56][20].run()  ;
            end
            begin
              mem_check[56][20].run()  ;
            end
            begin
              rf_driver[56][20].run()  ;
            end

            begin
              gen[56][21].run()  ;
            end
            begin
              drv[56][21].run()  ;
            end
            begin
              mem_check[56][21].run()  ;
            end
            begin
              rf_driver[56][21].run()  ;
            end

            begin
              gen[56][22].run()  ;
            end
            begin
              drv[56][22].run()  ;
            end
            begin
              mem_check[56][22].run()  ;
            end
            begin
              rf_driver[56][22].run()  ;
            end

            begin
              gen[56][23].run()  ;
            end
            begin
              drv[56][23].run()  ;
            end
            begin
              mem_check[56][23].run()  ;
            end
            begin
              rf_driver[56][23].run()  ;
            end

            begin
              gen[56][24].run()  ;
            end
            begin
              drv[56][24].run()  ;
            end
            begin
              mem_check[56][24].run()  ;
            end
            begin
              rf_driver[56][24].run()  ;
            end

            begin
              gen[56][25].run()  ;
            end
            begin
              drv[56][25].run()  ;
            end
            begin
              mem_check[56][25].run()  ;
            end
            begin
              rf_driver[56][25].run()  ;
            end

            begin
              gen[56][26].run()  ;
            end
            begin
              drv[56][26].run()  ;
            end
            begin
              mem_check[56][26].run()  ;
            end
            begin
              rf_driver[56][26].run()  ;
            end

            begin
              gen[56][27].run()  ;
            end
            begin
              drv[56][27].run()  ;
            end
            begin
              mem_check[56][27].run()  ;
            end
            begin
              rf_driver[56][27].run()  ;
            end

            begin
              gen[56][28].run()  ;
            end
            begin
              drv[56][28].run()  ;
            end
            begin
              mem_check[56][28].run()  ;
            end
            begin
              rf_driver[56][28].run()  ;
            end

            begin
              gen[56][29].run()  ;
            end
            begin
              drv[56][29].run()  ;
            end
            begin
              mem_check[56][29].run()  ;
            end
            begin
              rf_driver[56][29].run()  ;
            end

            begin
              gen[56][30].run()  ;
            end
            begin
              drv[56][30].run()  ;
            end
            begin
              mem_check[56][30].run()  ;
            end
            begin
              rf_driver[56][30].run()  ;
            end

            begin
              gen[56][31].run()  ;
            end
            begin
              drv[56][31].run()  ;
            end
            begin
              mem_check[56][31].run()  ;
            end
            begin
              rf_driver[56][31].run()  ;
            end

            begin
              ldst_driver[57].run()  ;
            end
            begin
              mgr[57].run()  ;
            end
            begin
              oob_drv[57].run()  ;
            end
            begin
              up_check[57].run()  ;
            end
            begin
              gen[57][0].run()  ;
            end
            begin
              drv[57][0].run()  ;
            end
            begin
              mem_check[57][0].run()  ;
            end
            begin
              rf_driver[57][0].run()  ;
            end

            begin
              gen[57][1].run()  ;
            end
            begin
              drv[57][1].run()  ;
            end
            begin
              mem_check[57][1].run()  ;
            end
            begin
              rf_driver[57][1].run()  ;
            end

            begin
              gen[57][2].run()  ;
            end
            begin
              drv[57][2].run()  ;
            end
            begin
              mem_check[57][2].run()  ;
            end
            begin
              rf_driver[57][2].run()  ;
            end

            begin
              gen[57][3].run()  ;
            end
            begin
              drv[57][3].run()  ;
            end
            begin
              mem_check[57][3].run()  ;
            end
            begin
              rf_driver[57][3].run()  ;
            end

            begin
              gen[57][4].run()  ;
            end
            begin
              drv[57][4].run()  ;
            end
            begin
              mem_check[57][4].run()  ;
            end
            begin
              rf_driver[57][4].run()  ;
            end

            begin
              gen[57][5].run()  ;
            end
            begin
              drv[57][5].run()  ;
            end
            begin
              mem_check[57][5].run()  ;
            end
            begin
              rf_driver[57][5].run()  ;
            end

            begin
              gen[57][6].run()  ;
            end
            begin
              drv[57][6].run()  ;
            end
            begin
              mem_check[57][6].run()  ;
            end
            begin
              rf_driver[57][6].run()  ;
            end

            begin
              gen[57][7].run()  ;
            end
            begin
              drv[57][7].run()  ;
            end
            begin
              mem_check[57][7].run()  ;
            end
            begin
              rf_driver[57][7].run()  ;
            end

            begin
              gen[57][8].run()  ;
            end
            begin
              drv[57][8].run()  ;
            end
            begin
              mem_check[57][8].run()  ;
            end
            begin
              rf_driver[57][8].run()  ;
            end

            begin
              gen[57][9].run()  ;
            end
            begin
              drv[57][9].run()  ;
            end
            begin
              mem_check[57][9].run()  ;
            end
            begin
              rf_driver[57][9].run()  ;
            end

            begin
              gen[57][10].run()  ;
            end
            begin
              drv[57][10].run()  ;
            end
            begin
              mem_check[57][10].run()  ;
            end
            begin
              rf_driver[57][10].run()  ;
            end

            begin
              gen[57][11].run()  ;
            end
            begin
              drv[57][11].run()  ;
            end
            begin
              mem_check[57][11].run()  ;
            end
            begin
              rf_driver[57][11].run()  ;
            end

            begin
              gen[57][12].run()  ;
            end
            begin
              drv[57][12].run()  ;
            end
            begin
              mem_check[57][12].run()  ;
            end
            begin
              rf_driver[57][12].run()  ;
            end

            begin
              gen[57][13].run()  ;
            end
            begin
              drv[57][13].run()  ;
            end
            begin
              mem_check[57][13].run()  ;
            end
            begin
              rf_driver[57][13].run()  ;
            end

            begin
              gen[57][14].run()  ;
            end
            begin
              drv[57][14].run()  ;
            end
            begin
              mem_check[57][14].run()  ;
            end
            begin
              rf_driver[57][14].run()  ;
            end

            begin
              gen[57][15].run()  ;
            end
            begin
              drv[57][15].run()  ;
            end
            begin
              mem_check[57][15].run()  ;
            end
            begin
              rf_driver[57][15].run()  ;
            end

            begin
              gen[57][16].run()  ;
            end
            begin
              drv[57][16].run()  ;
            end
            begin
              mem_check[57][16].run()  ;
            end
            begin
              rf_driver[57][16].run()  ;
            end

            begin
              gen[57][17].run()  ;
            end
            begin
              drv[57][17].run()  ;
            end
            begin
              mem_check[57][17].run()  ;
            end
            begin
              rf_driver[57][17].run()  ;
            end

            begin
              gen[57][18].run()  ;
            end
            begin
              drv[57][18].run()  ;
            end
            begin
              mem_check[57][18].run()  ;
            end
            begin
              rf_driver[57][18].run()  ;
            end

            begin
              gen[57][19].run()  ;
            end
            begin
              drv[57][19].run()  ;
            end
            begin
              mem_check[57][19].run()  ;
            end
            begin
              rf_driver[57][19].run()  ;
            end

            begin
              gen[57][20].run()  ;
            end
            begin
              drv[57][20].run()  ;
            end
            begin
              mem_check[57][20].run()  ;
            end
            begin
              rf_driver[57][20].run()  ;
            end

            begin
              gen[57][21].run()  ;
            end
            begin
              drv[57][21].run()  ;
            end
            begin
              mem_check[57][21].run()  ;
            end
            begin
              rf_driver[57][21].run()  ;
            end

            begin
              gen[57][22].run()  ;
            end
            begin
              drv[57][22].run()  ;
            end
            begin
              mem_check[57][22].run()  ;
            end
            begin
              rf_driver[57][22].run()  ;
            end

            begin
              gen[57][23].run()  ;
            end
            begin
              drv[57][23].run()  ;
            end
            begin
              mem_check[57][23].run()  ;
            end
            begin
              rf_driver[57][23].run()  ;
            end

            begin
              gen[57][24].run()  ;
            end
            begin
              drv[57][24].run()  ;
            end
            begin
              mem_check[57][24].run()  ;
            end
            begin
              rf_driver[57][24].run()  ;
            end

            begin
              gen[57][25].run()  ;
            end
            begin
              drv[57][25].run()  ;
            end
            begin
              mem_check[57][25].run()  ;
            end
            begin
              rf_driver[57][25].run()  ;
            end

            begin
              gen[57][26].run()  ;
            end
            begin
              drv[57][26].run()  ;
            end
            begin
              mem_check[57][26].run()  ;
            end
            begin
              rf_driver[57][26].run()  ;
            end

            begin
              gen[57][27].run()  ;
            end
            begin
              drv[57][27].run()  ;
            end
            begin
              mem_check[57][27].run()  ;
            end
            begin
              rf_driver[57][27].run()  ;
            end

            begin
              gen[57][28].run()  ;
            end
            begin
              drv[57][28].run()  ;
            end
            begin
              mem_check[57][28].run()  ;
            end
            begin
              rf_driver[57][28].run()  ;
            end

            begin
              gen[57][29].run()  ;
            end
            begin
              drv[57][29].run()  ;
            end
            begin
              mem_check[57][29].run()  ;
            end
            begin
              rf_driver[57][29].run()  ;
            end

            begin
              gen[57][30].run()  ;
            end
            begin
              drv[57][30].run()  ;
            end
            begin
              mem_check[57][30].run()  ;
            end
            begin
              rf_driver[57][30].run()  ;
            end

            begin
              gen[57][31].run()  ;
            end
            begin
              drv[57][31].run()  ;
            end
            begin
              mem_check[57][31].run()  ;
            end
            begin
              rf_driver[57][31].run()  ;
            end

            begin
              ldst_driver[58].run()  ;
            end
            begin
              mgr[58].run()  ;
            end
            begin
              oob_drv[58].run()  ;
            end
            begin
              up_check[58].run()  ;
            end
            begin
              gen[58][0].run()  ;
            end
            begin
              drv[58][0].run()  ;
            end
            begin
              mem_check[58][0].run()  ;
            end
            begin
              rf_driver[58][0].run()  ;
            end

            begin
              gen[58][1].run()  ;
            end
            begin
              drv[58][1].run()  ;
            end
            begin
              mem_check[58][1].run()  ;
            end
            begin
              rf_driver[58][1].run()  ;
            end

            begin
              gen[58][2].run()  ;
            end
            begin
              drv[58][2].run()  ;
            end
            begin
              mem_check[58][2].run()  ;
            end
            begin
              rf_driver[58][2].run()  ;
            end

            begin
              gen[58][3].run()  ;
            end
            begin
              drv[58][3].run()  ;
            end
            begin
              mem_check[58][3].run()  ;
            end
            begin
              rf_driver[58][3].run()  ;
            end

            begin
              gen[58][4].run()  ;
            end
            begin
              drv[58][4].run()  ;
            end
            begin
              mem_check[58][4].run()  ;
            end
            begin
              rf_driver[58][4].run()  ;
            end

            begin
              gen[58][5].run()  ;
            end
            begin
              drv[58][5].run()  ;
            end
            begin
              mem_check[58][5].run()  ;
            end
            begin
              rf_driver[58][5].run()  ;
            end

            begin
              gen[58][6].run()  ;
            end
            begin
              drv[58][6].run()  ;
            end
            begin
              mem_check[58][6].run()  ;
            end
            begin
              rf_driver[58][6].run()  ;
            end

            begin
              gen[58][7].run()  ;
            end
            begin
              drv[58][7].run()  ;
            end
            begin
              mem_check[58][7].run()  ;
            end
            begin
              rf_driver[58][7].run()  ;
            end

            begin
              gen[58][8].run()  ;
            end
            begin
              drv[58][8].run()  ;
            end
            begin
              mem_check[58][8].run()  ;
            end
            begin
              rf_driver[58][8].run()  ;
            end

            begin
              gen[58][9].run()  ;
            end
            begin
              drv[58][9].run()  ;
            end
            begin
              mem_check[58][9].run()  ;
            end
            begin
              rf_driver[58][9].run()  ;
            end

            begin
              gen[58][10].run()  ;
            end
            begin
              drv[58][10].run()  ;
            end
            begin
              mem_check[58][10].run()  ;
            end
            begin
              rf_driver[58][10].run()  ;
            end

            begin
              gen[58][11].run()  ;
            end
            begin
              drv[58][11].run()  ;
            end
            begin
              mem_check[58][11].run()  ;
            end
            begin
              rf_driver[58][11].run()  ;
            end

            begin
              gen[58][12].run()  ;
            end
            begin
              drv[58][12].run()  ;
            end
            begin
              mem_check[58][12].run()  ;
            end
            begin
              rf_driver[58][12].run()  ;
            end

            begin
              gen[58][13].run()  ;
            end
            begin
              drv[58][13].run()  ;
            end
            begin
              mem_check[58][13].run()  ;
            end
            begin
              rf_driver[58][13].run()  ;
            end

            begin
              gen[58][14].run()  ;
            end
            begin
              drv[58][14].run()  ;
            end
            begin
              mem_check[58][14].run()  ;
            end
            begin
              rf_driver[58][14].run()  ;
            end

            begin
              gen[58][15].run()  ;
            end
            begin
              drv[58][15].run()  ;
            end
            begin
              mem_check[58][15].run()  ;
            end
            begin
              rf_driver[58][15].run()  ;
            end

            begin
              gen[58][16].run()  ;
            end
            begin
              drv[58][16].run()  ;
            end
            begin
              mem_check[58][16].run()  ;
            end
            begin
              rf_driver[58][16].run()  ;
            end

            begin
              gen[58][17].run()  ;
            end
            begin
              drv[58][17].run()  ;
            end
            begin
              mem_check[58][17].run()  ;
            end
            begin
              rf_driver[58][17].run()  ;
            end

            begin
              gen[58][18].run()  ;
            end
            begin
              drv[58][18].run()  ;
            end
            begin
              mem_check[58][18].run()  ;
            end
            begin
              rf_driver[58][18].run()  ;
            end

            begin
              gen[58][19].run()  ;
            end
            begin
              drv[58][19].run()  ;
            end
            begin
              mem_check[58][19].run()  ;
            end
            begin
              rf_driver[58][19].run()  ;
            end

            begin
              gen[58][20].run()  ;
            end
            begin
              drv[58][20].run()  ;
            end
            begin
              mem_check[58][20].run()  ;
            end
            begin
              rf_driver[58][20].run()  ;
            end

            begin
              gen[58][21].run()  ;
            end
            begin
              drv[58][21].run()  ;
            end
            begin
              mem_check[58][21].run()  ;
            end
            begin
              rf_driver[58][21].run()  ;
            end

            begin
              gen[58][22].run()  ;
            end
            begin
              drv[58][22].run()  ;
            end
            begin
              mem_check[58][22].run()  ;
            end
            begin
              rf_driver[58][22].run()  ;
            end

            begin
              gen[58][23].run()  ;
            end
            begin
              drv[58][23].run()  ;
            end
            begin
              mem_check[58][23].run()  ;
            end
            begin
              rf_driver[58][23].run()  ;
            end

            begin
              gen[58][24].run()  ;
            end
            begin
              drv[58][24].run()  ;
            end
            begin
              mem_check[58][24].run()  ;
            end
            begin
              rf_driver[58][24].run()  ;
            end

            begin
              gen[58][25].run()  ;
            end
            begin
              drv[58][25].run()  ;
            end
            begin
              mem_check[58][25].run()  ;
            end
            begin
              rf_driver[58][25].run()  ;
            end

            begin
              gen[58][26].run()  ;
            end
            begin
              drv[58][26].run()  ;
            end
            begin
              mem_check[58][26].run()  ;
            end
            begin
              rf_driver[58][26].run()  ;
            end

            begin
              gen[58][27].run()  ;
            end
            begin
              drv[58][27].run()  ;
            end
            begin
              mem_check[58][27].run()  ;
            end
            begin
              rf_driver[58][27].run()  ;
            end

            begin
              gen[58][28].run()  ;
            end
            begin
              drv[58][28].run()  ;
            end
            begin
              mem_check[58][28].run()  ;
            end
            begin
              rf_driver[58][28].run()  ;
            end

            begin
              gen[58][29].run()  ;
            end
            begin
              drv[58][29].run()  ;
            end
            begin
              mem_check[58][29].run()  ;
            end
            begin
              rf_driver[58][29].run()  ;
            end

            begin
              gen[58][30].run()  ;
            end
            begin
              drv[58][30].run()  ;
            end
            begin
              mem_check[58][30].run()  ;
            end
            begin
              rf_driver[58][30].run()  ;
            end

            begin
              gen[58][31].run()  ;
            end
            begin
              drv[58][31].run()  ;
            end
            begin
              mem_check[58][31].run()  ;
            end
            begin
              rf_driver[58][31].run()  ;
            end

            begin
              ldst_driver[59].run()  ;
            end
            begin
              mgr[59].run()  ;
            end
            begin
              oob_drv[59].run()  ;
            end
            begin
              up_check[59].run()  ;
            end
            begin
              gen[59][0].run()  ;
            end
            begin
              drv[59][0].run()  ;
            end
            begin
              mem_check[59][0].run()  ;
            end
            begin
              rf_driver[59][0].run()  ;
            end

            begin
              gen[59][1].run()  ;
            end
            begin
              drv[59][1].run()  ;
            end
            begin
              mem_check[59][1].run()  ;
            end
            begin
              rf_driver[59][1].run()  ;
            end

            begin
              gen[59][2].run()  ;
            end
            begin
              drv[59][2].run()  ;
            end
            begin
              mem_check[59][2].run()  ;
            end
            begin
              rf_driver[59][2].run()  ;
            end

            begin
              gen[59][3].run()  ;
            end
            begin
              drv[59][3].run()  ;
            end
            begin
              mem_check[59][3].run()  ;
            end
            begin
              rf_driver[59][3].run()  ;
            end

            begin
              gen[59][4].run()  ;
            end
            begin
              drv[59][4].run()  ;
            end
            begin
              mem_check[59][4].run()  ;
            end
            begin
              rf_driver[59][4].run()  ;
            end

            begin
              gen[59][5].run()  ;
            end
            begin
              drv[59][5].run()  ;
            end
            begin
              mem_check[59][5].run()  ;
            end
            begin
              rf_driver[59][5].run()  ;
            end

            begin
              gen[59][6].run()  ;
            end
            begin
              drv[59][6].run()  ;
            end
            begin
              mem_check[59][6].run()  ;
            end
            begin
              rf_driver[59][6].run()  ;
            end

            begin
              gen[59][7].run()  ;
            end
            begin
              drv[59][7].run()  ;
            end
            begin
              mem_check[59][7].run()  ;
            end
            begin
              rf_driver[59][7].run()  ;
            end

            begin
              gen[59][8].run()  ;
            end
            begin
              drv[59][8].run()  ;
            end
            begin
              mem_check[59][8].run()  ;
            end
            begin
              rf_driver[59][8].run()  ;
            end

            begin
              gen[59][9].run()  ;
            end
            begin
              drv[59][9].run()  ;
            end
            begin
              mem_check[59][9].run()  ;
            end
            begin
              rf_driver[59][9].run()  ;
            end

            begin
              gen[59][10].run()  ;
            end
            begin
              drv[59][10].run()  ;
            end
            begin
              mem_check[59][10].run()  ;
            end
            begin
              rf_driver[59][10].run()  ;
            end

            begin
              gen[59][11].run()  ;
            end
            begin
              drv[59][11].run()  ;
            end
            begin
              mem_check[59][11].run()  ;
            end
            begin
              rf_driver[59][11].run()  ;
            end

            begin
              gen[59][12].run()  ;
            end
            begin
              drv[59][12].run()  ;
            end
            begin
              mem_check[59][12].run()  ;
            end
            begin
              rf_driver[59][12].run()  ;
            end

            begin
              gen[59][13].run()  ;
            end
            begin
              drv[59][13].run()  ;
            end
            begin
              mem_check[59][13].run()  ;
            end
            begin
              rf_driver[59][13].run()  ;
            end

            begin
              gen[59][14].run()  ;
            end
            begin
              drv[59][14].run()  ;
            end
            begin
              mem_check[59][14].run()  ;
            end
            begin
              rf_driver[59][14].run()  ;
            end

            begin
              gen[59][15].run()  ;
            end
            begin
              drv[59][15].run()  ;
            end
            begin
              mem_check[59][15].run()  ;
            end
            begin
              rf_driver[59][15].run()  ;
            end

            begin
              gen[59][16].run()  ;
            end
            begin
              drv[59][16].run()  ;
            end
            begin
              mem_check[59][16].run()  ;
            end
            begin
              rf_driver[59][16].run()  ;
            end

            begin
              gen[59][17].run()  ;
            end
            begin
              drv[59][17].run()  ;
            end
            begin
              mem_check[59][17].run()  ;
            end
            begin
              rf_driver[59][17].run()  ;
            end

            begin
              gen[59][18].run()  ;
            end
            begin
              drv[59][18].run()  ;
            end
            begin
              mem_check[59][18].run()  ;
            end
            begin
              rf_driver[59][18].run()  ;
            end

            begin
              gen[59][19].run()  ;
            end
            begin
              drv[59][19].run()  ;
            end
            begin
              mem_check[59][19].run()  ;
            end
            begin
              rf_driver[59][19].run()  ;
            end

            begin
              gen[59][20].run()  ;
            end
            begin
              drv[59][20].run()  ;
            end
            begin
              mem_check[59][20].run()  ;
            end
            begin
              rf_driver[59][20].run()  ;
            end

            begin
              gen[59][21].run()  ;
            end
            begin
              drv[59][21].run()  ;
            end
            begin
              mem_check[59][21].run()  ;
            end
            begin
              rf_driver[59][21].run()  ;
            end

            begin
              gen[59][22].run()  ;
            end
            begin
              drv[59][22].run()  ;
            end
            begin
              mem_check[59][22].run()  ;
            end
            begin
              rf_driver[59][22].run()  ;
            end

            begin
              gen[59][23].run()  ;
            end
            begin
              drv[59][23].run()  ;
            end
            begin
              mem_check[59][23].run()  ;
            end
            begin
              rf_driver[59][23].run()  ;
            end

            begin
              gen[59][24].run()  ;
            end
            begin
              drv[59][24].run()  ;
            end
            begin
              mem_check[59][24].run()  ;
            end
            begin
              rf_driver[59][24].run()  ;
            end

            begin
              gen[59][25].run()  ;
            end
            begin
              drv[59][25].run()  ;
            end
            begin
              mem_check[59][25].run()  ;
            end
            begin
              rf_driver[59][25].run()  ;
            end

            begin
              gen[59][26].run()  ;
            end
            begin
              drv[59][26].run()  ;
            end
            begin
              mem_check[59][26].run()  ;
            end
            begin
              rf_driver[59][26].run()  ;
            end

            begin
              gen[59][27].run()  ;
            end
            begin
              drv[59][27].run()  ;
            end
            begin
              mem_check[59][27].run()  ;
            end
            begin
              rf_driver[59][27].run()  ;
            end

            begin
              gen[59][28].run()  ;
            end
            begin
              drv[59][28].run()  ;
            end
            begin
              mem_check[59][28].run()  ;
            end
            begin
              rf_driver[59][28].run()  ;
            end

            begin
              gen[59][29].run()  ;
            end
            begin
              drv[59][29].run()  ;
            end
            begin
              mem_check[59][29].run()  ;
            end
            begin
              rf_driver[59][29].run()  ;
            end

            begin
              gen[59][30].run()  ;
            end
            begin
              drv[59][30].run()  ;
            end
            begin
              mem_check[59][30].run()  ;
            end
            begin
              rf_driver[59][30].run()  ;
            end

            begin
              gen[59][31].run()  ;
            end
            begin
              drv[59][31].run()  ;
            end
            begin
              mem_check[59][31].run()  ;
            end
            begin
              rf_driver[59][31].run()  ;
            end

            begin
              ldst_driver[60].run()  ;
            end
            begin
              mgr[60].run()  ;
            end
            begin
              oob_drv[60].run()  ;
            end
            begin
              up_check[60].run()  ;
            end
            begin
              gen[60][0].run()  ;
            end
            begin
              drv[60][0].run()  ;
            end
            begin
              mem_check[60][0].run()  ;
            end
            begin
              rf_driver[60][0].run()  ;
            end

            begin
              gen[60][1].run()  ;
            end
            begin
              drv[60][1].run()  ;
            end
            begin
              mem_check[60][1].run()  ;
            end
            begin
              rf_driver[60][1].run()  ;
            end

            begin
              gen[60][2].run()  ;
            end
            begin
              drv[60][2].run()  ;
            end
            begin
              mem_check[60][2].run()  ;
            end
            begin
              rf_driver[60][2].run()  ;
            end

            begin
              gen[60][3].run()  ;
            end
            begin
              drv[60][3].run()  ;
            end
            begin
              mem_check[60][3].run()  ;
            end
            begin
              rf_driver[60][3].run()  ;
            end

            begin
              gen[60][4].run()  ;
            end
            begin
              drv[60][4].run()  ;
            end
            begin
              mem_check[60][4].run()  ;
            end
            begin
              rf_driver[60][4].run()  ;
            end

            begin
              gen[60][5].run()  ;
            end
            begin
              drv[60][5].run()  ;
            end
            begin
              mem_check[60][5].run()  ;
            end
            begin
              rf_driver[60][5].run()  ;
            end

            begin
              gen[60][6].run()  ;
            end
            begin
              drv[60][6].run()  ;
            end
            begin
              mem_check[60][6].run()  ;
            end
            begin
              rf_driver[60][6].run()  ;
            end

            begin
              gen[60][7].run()  ;
            end
            begin
              drv[60][7].run()  ;
            end
            begin
              mem_check[60][7].run()  ;
            end
            begin
              rf_driver[60][7].run()  ;
            end

            begin
              gen[60][8].run()  ;
            end
            begin
              drv[60][8].run()  ;
            end
            begin
              mem_check[60][8].run()  ;
            end
            begin
              rf_driver[60][8].run()  ;
            end

            begin
              gen[60][9].run()  ;
            end
            begin
              drv[60][9].run()  ;
            end
            begin
              mem_check[60][9].run()  ;
            end
            begin
              rf_driver[60][9].run()  ;
            end

            begin
              gen[60][10].run()  ;
            end
            begin
              drv[60][10].run()  ;
            end
            begin
              mem_check[60][10].run()  ;
            end
            begin
              rf_driver[60][10].run()  ;
            end

            begin
              gen[60][11].run()  ;
            end
            begin
              drv[60][11].run()  ;
            end
            begin
              mem_check[60][11].run()  ;
            end
            begin
              rf_driver[60][11].run()  ;
            end

            begin
              gen[60][12].run()  ;
            end
            begin
              drv[60][12].run()  ;
            end
            begin
              mem_check[60][12].run()  ;
            end
            begin
              rf_driver[60][12].run()  ;
            end

            begin
              gen[60][13].run()  ;
            end
            begin
              drv[60][13].run()  ;
            end
            begin
              mem_check[60][13].run()  ;
            end
            begin
              rf_driver[60][13].run()  ;
            end

            begin
              gen[60][14].run()  ;
            end
            begin
              drv[60][14].run()  ;
            end
            begin
              mem_check[60][14].run()  ;
            end
            begin
              rf_driver[60][14].run()  ;
            end

            begin
              gen[60][15].run()  ;
            end
            begin
              drv[60][15].run()  ;
            end
            begin
              mem_check[60][15].run()  ;
            end
            begin
              rf_driver[60][15].run()  ;
            end

            begin
              gen[60][16].run()  ;
            end
            begin
              drv[60][16].run()  ;
            end
            begin
              mem_check[60][16].run()  ;
            end
            begin
              rf_driver[60][16].run()  ;
            end

            begin
              gen[60][17].run()  ;
            end
            begin
              drv[60][17].run()  ;
            end
            begin
              mem_check[60][17].run()  ;
            end
            begin
              rf_driver[60][17].run()  ;
            end

            begin
              gen[60][18].run()  ;
            end
            begin
              drv[60][18].run()  ;
            end
            begin
              mem_check[60][18].run()  ;
            end
            begin
              rf_driver[60][18].run()  ;
            end

            begin
              gen[60][19].run()  ;
            end
            begin
              drv[60][19].run()  ;
            end
            begin
              mem_check[60][19].run()  ;
            end
            begin
              rf_driver[60][19].run()  ;
            end

            begin
              gen[60][20].run()  ;
            end
            begin
              drv[60][20].run()  ;
            end
            begin
              mem_check[60][20].run()  ;
            end
            begin
              rf_driver[60][20].run()  ;
            end

            begin
              gen[60][21].run()  ;
            end
            begin
              drv[60][21].run()  ;
            end
            begin
              mem_check[60][21].run()  ;
            end
            begin
              rf_driver[60][21].run()  ;
            end

            begin
              gen[60][22].run()  ;
            end
            begin
              drv[60][22].run()  ;
            end
            begin
              mem_check[60][22].run()  ;
            end
            begin
              rf_driver[60][22].run()  ;
            end

            begin
              gen[60][23].run()  ;
            end
            begin
              drv[60][23].run()  ;
            end
            begin
              mem_check[60][23].run()  ;
            end
            begin
              rf_driver[60][23].run()  ;
            end

            begin
              gen[60][24].run()  ;
            end
            begin
              drv[60][24].run()  ;
            end
            begin
              mem_check[60][24].run()  ;
            end
            begin
              rf_driver[60][24].run()  ;
            end

            begin
              gen[60][25].run()  ;
            end
            begin
              drv[60][25].run()  ;
            end
            begin
              mem_check[60][25].run()  ;
            end
            begin
              rf_driver[60][25].run()  ;
            end

            begin
              gen[60][26].run()  ;
            end
            begin
              drv[60][26].run()  ;
            end
            begin
              mem_check[60][26].run()  ;
            end
            begin
              rf_driver[60][26].run()  ;
            end

            begin
              gen[60][27].run()  ;
            end
            begin
              drv[60][27].run()  ;
            end
            begin
              mem_check[60][27].run()  ;
            end
            begin
              rf_driver[60][27].run()  ;
            end

            begin
              gen[60][28].run()  ;
            end
            begin
              drv[60][28].run()  ;
            end
            begin
              mem_check[60][28].run()  ;
            end
            begin
              rf_driver[60][28].run()  ;
            end

            begin
              gen[60][29].run()  ;
            end
            begin
              drv[60][29].run()  ;
            end
            begin
              mem_check[60][29].run()  ;
            end
            begin
              rf_driver[60][29].run()  ;
            end

            begin
              gen[60][30].run()  ;
            end
            begin
              drv[60][30].run()  ;
            end
            begin
              mem_check[60][30].run()  ;
            end
            begin
              rf_driver[60][30].run()  ;
            end

            begin
              gen[60][31].run()  ;
            end
            begin
              drv[60][31].run()  ;
            end
            begin
              mem_check[60][31].run()  ;
            end
            begin
              rf_driver[60][31].run()  ;
            end

            begin
              ldst_driver[61].run()  ;
            end
            begin
              mgr[61].run()  ;
            end
            begin
              oob_drv[61].run()  ;
            end
            begin
              up_check[61].run()  ;
            end
            begin
              gen[61][0].run()  ;
            end
            begin
              drv[61][0].run()  ;
            end
            begin
              mem_check[61][0].run()  ;
            end
            begin
              rf_driver[61][0].run()  ;
            end

            begin
              gen[61][1].run()  ;
            end
            begin
              drv[61][1].run()  ;
            end
            begin
              mem_check[61][1].run()  ;
            end
            begin
              rf_driver[61][1].run()  ;
            end

            begin
              gen[61][2].run()  ;
            end
            begin
              drv[61][2].run()  ;
            end
            begin
              mem_check[61][2].run()  ;
            end
            begin
              rf_driver[61][2].run()  ;
            end

            begin
              gen[61][3].run()  ;
            end
            begin
              drv[61][3].run()  ;
            end
            begin
              mem_check[61][3].run()  ;
            end
            begin
              rf_driver[61][3].run()  ;
            end

            begin
              gen[61][4].run()  ;
            end
            begin
              drv[61][4].run()  ;
            end
            begin
              mem_check[61][4].run()  ;
            end
            begin
              rf_driver[61][4].run()  ;
            end

            begin
              gen[61][5].run()  ;
            end
            begin
              drv[61][5].run()  ;
            end
            begin
              mem_check[61][5].run()  ;
            end
            begin
              rf_driver[61][5].run()  ;
            end

            begin
              gen[61][6].run()  ;
            end
            begin
              drv[61][6].run()  ;
            end
            begin
              mem_check[61][6].run()  ;
            end
            begin
              rf_driver[61][6].run()  ;
            end

            begin
              gen[61][7].run()  ;
            end
            begin
              drv[61][7].run()  ;
            end
            begin
              mem_check[61][7].run()  ;
            end
            begin
              rf_driver[61][7].run()  ;
            end

            begin
              gen[61][8].run()  ;
            end
            begin
              drv[61][8].run()  ;
            end
            begin
              mem_check[61][8].run()  ;
            end
            begin
              rf_driver[61][8].run()  ;
            end

            begin
              gen[61][9].run()  ;
            end
            begin
              drv[61][9].run()  ;
            end
            begin
              mem_check[61][9].run()  ;
            end
            begin
              rf_driver[61][9].run()  ;
            end

            begin
              gen[61][10].run()  ;
            end
            begin
              drv[61][10].run()  ;
            end
            begin
              mem_check[61][10].run()  ;
            end
            begin
              rf_driver[61][10].run()  ;
            end

            begin
              gen[61][11].run()  ;
            end
            begin
              drv[61][11].run()  ;
            end
            begin
              mem_check[61][11].run()  ;
            end
            begin
              rf_driver[61][11].run()  ;
            end

            begin
              gen[61][12].run()  ;
            end
            begin
              drv[61][12].run()  ;
            end
            begin
              mem_check[61][12].run()  ;
            end
            begin
              rf_driver[61][12].run()  ;
            end

            begin
              gen[61][13].run()  ;
            end
            begin
              drv[61][13].run()  ;
            end
            begin
              mem_check[61][13].run()  ;
            end
            begin
              rf_driver[61][13].run()  ;
            end

            begin
              gen[61][14].run()  ;
            end
            begin
              drv[61][14].run()  ;
            end
            begin
              mem_check[61][14].run()  ;
            end
            begin
              rf_driver[61][14].run()  ;
            end

            begin
              gen[61][15].run()  ;
            end
            begin
              drv[61][15].run()  ;
            end
            begin
              mem_check[61][15].run()  ;
            end
            begin
              rf_driver[61][15].run()  ;
            end

            begin
              gen[61][16].run()  ;
            end
            begin
              drv[61][16].run()  ;
            end
            begin
              mem_check[61][16].run()  ;
            end
            begin
              rf_driver[61][16].run()  ;
            end

            begin
              gen[61][17].run()  ;
            end
            begin
              drv[61][17].run()  ;
            end
            begin
              mem_check[61][17].run()  ;
            end
            begin
              rf_driver[61][17].run()  ;
            end

            begin
              gen[61][18].run()  ;
            end
            begin
              drv[61][18].run()  ;
            end
            begin
              mem_check[61][18].run()  ;
            end
            begin
              rf_driver[61][18].run()  ;
            end

            begin
              gen[61][19].run()  ;
            end
            begin
              drv[61][19].run()  ;
            end
            begin
              mem_check[61][19].run()  ;
            end
            begin
              rf_driver[61][19].run()  ;
            end

            begin
              gen[61][20].run()  ;
            end
            begin
              drv[61][20].run()  ;
            end
            begin
              mem_check[61][20].run()  ;
            end
            begin
              rf_driver[61][20].run()  ;
            end

            begin
              gen[61][21].run()  ;
            end
            begin
              drv[61][21].run()  ;
            end
            begin
              mem_check[61][21].run()  ;
            end
            begin
              rf_driver[61][21].run()  ;
            end

            begin
              gen[61][22].run()  ;
            end
            begin
              drv[61][22].run()  ;
            end
            begin
              mem_check[61][22].run()  ;
            end
            begin
              rf_driver[61][22].run()  ;
            end

            begin
              gen[61][23].run()  ;
            end
            begin
              drv[61][23].run()  ;
            end
            begin
              mem_check[61][23].run()  ;
            end
            begin
              rf_driver[61][23].run()  ;
            end

            begin
              gen[61][24].run()  ;
            end
            begin
              drv[61][24].run()  ;
            end
            begin
              mem_check[61][24].run()  ;
            end
            begin
              rf_driver[61][24].run()  ;
            end

            begin
              gen[61][25].run()  ;
            end
            begin
              drv[61][25].run()  ;
            end
            begin
              mem_check[61][25].run()  ;
            end
            begin
              rf_driver[61][25].run()  ;
            end

            begin
              gen[61][26].run()  ;
            end
            begin
              drv[61][26].run()  ;
            end
            begin
              mem_check[61][26].run()  ;
            end
            begin
              rf_driver[61][26].run()  ;
            end

            begin
              gen[61][27].run()  ;
            end
            begin
              drv[61][27].run()  ;
            end
            begin
              mem_check[61][27].run()  ;
            end
            begin
              rf_driver[61][27].run()  ;
            end

            begin
              gen[61][28].run()  ;
            end
            begin
              drv[61][28].run()  ;
            end
            begin
              mem_check[61][28].run()  ;
            end
            begin
              rf_driver[61][28].run()  ;
            end

            begin
              gen[61][29].run()  ;
            end
            begin
              drv[61][29].run()  ;
            end
            begin
              mem_check[61][29].run()  ;
            end
            begin
              rf_driver[61][29].run()  ;
            end

            begin
              gen[61][30].run()  ;
            end
            begin
              drv[61][30].run()  ;
            end
            begin
              mem_check[61][30].run()  ;
            end
            begin
              rf_driver[61][30].run()  ;
            end

            begin
              gen[61][31].run()  ;
            end
            begin
              drv[61][31].run()  ;
            end
            begin
              mem_check[61][31].run()  ;
            end
            begin
              rf_driver[61][31].run()  ;
            end

            begin
              ldst_driver[62].run()  ;
            end
            begin
              mgr[62].run()  ;
            end
            begin
              oob_drv[62].run()  ;
            end
            begin
              up_check[62].run()  ;
            end
            begin
              gen[62][0].run()  ;
            end
            begin
              drv[62][0].run()  ;
            end
            begin
              mem_check[62][0].run()  ;
            end
            begin
              rf_driver[62][0].run()  ;
            end

            begin
              gen[62][1].run()  ;
            end
            begin
              drv[62][1].run()  ;
            end
            begin
              mem_check[62][1].run()  ;
            end
            begin
              rf_driver[62][1].run()  ;
            end

            begin
              gen[62][2].run()  ;
            end
            begin
              drv[62][2].run()  ;
            end
            begin
              mem_check[62][2].run()  ;
            end
            begin
              rf_driver[62][2].run()  ;
            end

            begin
              gen[62][3].run()  ;
            end
            begin
              drv[62][3].run()  ;
            end
            begin
              mem_check[62][3].run()  ;
            end
            begin
              rf_driver[62][3].run()  ;
            end

            begin
              gen[62][4].run()  ;
            end
            begin
              drv[62][4].run()  ;
            end
            begin
              mem_check[62][4].run()  ;
            end
            begin
              rf_driver[62][4].run()  ;
            end

            begin
              gen[62][5].run()  ;
            end
            begin
              drv[62][5].run()  ;
            end
            begin
              mem_check[62][5].run()  ;
            end
            begin
              rf_driver[62][5].run()  ;
            end

            begin
              gen[62][6].run()  ;
            end
            begin
              drv[62][6].run()  ;
            end
            begin
              mem_check[62][6].run()  ;
            end
            begin
              rf_driver[62][6].run()  ;
            end

            begin
              gen[62][7].run()  ;
            end
            begin
              drv[62][7].run()  ;
            end
            begin
              mem_check[62][7].run()  ;
            end
            begin
              rf_driver[62][7].run()  ;
            end

            begin
              gen[62][8].run()  ;
            end
            begin
              drv[62][8].run()  ;
            end
            begin
              mem_check[62][8].run()  ;
            end
            begin
              rf_driver[62][8].run()  ;
            end

            begin
              gen[62][9].run()  ;
            end
            begin
              drv[62][9].run()  ;
            end
            begin
              mem_check[62][9].run()  ;
            end
            begin
              rf_driver[62][9].run()  ;
            end

            begin
              gen[62][10].run()  ;
            end
            begin
              drv[62][10].run()  ;
            end
            begin
              mem_check[62][10].run()  ;
            end
            begin
              rf_driver[62][10].run()  ;
            end

            begin
              gen[62][11].run()  ;
            end
            begin
              drv[62][11].run()  ;
            end
            begin
              mem_check[62][11].run()  ;
            end
            begin
              rf_driver[62][11].run()  ;
            end

            begin
              gen[62][12].run()  ;
            end
            begin
              drv[62][12].run()  ;
            end
            begin
              mem_check[62][12].run()  ;
            end
            begin
              rf_driver[62][12].run()  ;
            end

            begin
              gen[62][13].run()  ;
            end
            begin
              drv[62][13].run()  ;
            end
            begin
              mem_check[62][13].run()  ;
            end
            begin
              rf_driver[62][13].run()  ;
            end

            begin
              gen[62][14].run()  ;
            end
            begin
              drv[62][14].run()  ;
            end
            begin
              mem_check[62][14].run()  ;
            end
            begin
              rf_driver[62][14].run()  ;
            end

            begin
              gen[62][15].run()  ;
            end
            begin
              drv[62][15].run()  ;
            end
            begin
              mem_check[62][15].run()  ;
            end
            begin
              rf_driver[62][15].run()  ;
            end

            begin
              gen[62][16].run()  ;
            end
            begin
              drv[62][16].run()  ;
            end
            begin
              mem_check[62][16].run()  ;
            end
            begin
              rf_driver[62][16].run()  ;
            end

            begin
              gen[62][17].run()  ;
            end
            begin
              drv[62][17].run()  ;
            end
            begin
              mem_check[62][17].run()  ;
            end
            begin
              rf_driver[62][17].run()  ;
            end

            begin
              gen[62][18].run()  ;
            end
            begin
              drv[62][18].run()  ;
            end
            begin
              mem_check[62][18].run()  ;
            end
            begin
              rf_driver[62][18].run()  ;
            end

            begin
              gen[62][19].run()  ;
            end
            begin
              drv[62][19].run()  ;
            end
            begin
              mem_check[62][19].run()  ;
            end
            begin
              rf_driver[62][19].run()  ;
            end

            begin
              gen[62][20].run()  ;
            end
            begin
              drv[62][20].run()  ;
            end
            begin
              mem_check[62][20].run()  ;
            end
            begin
              rf_driver[62][20].run()  ;
            end

            begin
              gen[62][21].run()  ;
            end
            begin
              drv[62][21].run()  ;
            end
            begin
              mem_check[62][21].run()  ;
            end
            begin
              rf_driver[62][21].run()  ;
            end

            begin
              gen[62][22].run()  ;
            end
            begin
              drv[62][22].run()  ;
            end
            begin
              mem_check[62][22].run()  ;
            end
            begin
              rf_driver[62][22].run()  ;
            end

            begin
              gen[62][23].run()  ;
            end
            begin
              drv[62][23].run()  ;
            end
            begin
              mem_check[62][23].run()  ;
            end
            begin
              rf_driver[62][23].run()  ;
            end

            begin
              gen[62][24].run()  ;
            end
            begin
              drv[62][24].run()  ;
            end
            begin
              mem_check[62][24].run()  ;
            end
            begin
              rf_driver[62][24].run()  ;
            end

            begin
              gen[62][25].run()  ;
            end
            begin
              drv[62][25].run()  ;
            end
            begin
              mem_check[62][25].run()  ;
            end
            begin
              rf_driver[62][25].run()  ;
            end

            begin
              gen[62][26].run()  ;
            end
            begin
              drv[62][26].run()  ;
            end
            begin
              mem_check[62][26].run()  ;
            end
            begin
              rf_driver[62][26].run()  ;
            end

            begin
              gen[62][27].run()  ;
            end
            begin
              drv[62][27].run()  ;
            end
            begin
              mem_check[62][27].run()  ;
            end
            begin
              rf_driver[62][27].run()  ;
            end

            begin
              gen[62][28].run()  ;
            end
            begin
              drv[62][28].run()  ;
            end
            begin
              mem_check[62][28].run()  ;
            end
            begin
              rf_driver[62][28].run()  ;
            end

            begin
              gen[62][29].run()  ;
            end
            begin
              drv[62][29].run()  ;
            end
            begin
              mem_check[62][29].run()  ;
            end
            begin
              rf_driver[62][29].run()  ;
            end

            begin
              gen[62][30].run()  ;
            end
            begin
              drv[62][30].run()  ;
            end
            begin
              mem_check[62][30].run()  ;
            end
            begin
              rf_driver[62][30].run()  ;
            end

            begin
              gen[62][31].run()  ;
            end
            begin
              drv[62][31].run()  ;
            end
            begin
              mem_check[62][31].run()  ;
            end
            begin
              rf_driver[62][31].run()  ;
            end

            begin
              ldst_driver[63].run()  ;
            end
            begin
              mgr[63].run()  ;
            end
            begin
              oob_drv[63].run()  ;
            end
            begin
              up_check[63].run()  ;
            end
            begin
              gen[63][0].run()  ;
            end
            begin
              drv[63][0].run()  ;
            end
            begin
              mem_check[63][0].run()  ;
            end
            begin
              rf_driver[63][0].run()  ;
            end

            begin
              gen[63][1].run()  ;
            end
            begin
              drv[63][1].run()  ;
            end
            begin
              mem_check[63][1].run()  ;
            end
            begin
              rf_driver[63][1].run()  ;
            end

            begin
              gen[63][2].run()  ;
            end
            begin
              drv[63][2].run()  ;
            end
            begin
              mem_check[63][2].run()  ;
            end
            begin
              rf_driver[63][2].run()  ;
            end

            begin
              gen[63][3].run()  ;
            end
            begin
              drv[63][3].run()  ;
            end
            begin
              mem_check[63][3].run()  ;
            end
            begin
              rf_driver[63][3].run()  ;
            end

            begin
              gen[63][4].run()  ;
            end
            begin
              drv[63][4].run()  ;
            end
            begin
              mem_check[63][4].run()  ;
            end
            begin
              rf_driver[63][4].run()  ;
            end

            begin
              gen[63][5].run()  ;
            end
            begin
              drv[63][5].run()  ;
            end
            begin
              mem_check[63][5].run()  ;
            end
            begin
              rf_driver[63][5].run()  ;
            end

            begin
              gen[63][6].run()  ;
            end
            begin
              drv[63][6].run()  ;
            end
            begin
              mem_check[63][6].run()  ;
            end
            begin
              rf_driver[63][6].run()  ;
            end

            begin
              gen[63][7].run()  ;
            end
            begin
              drv[63][7].run()  ;
            end
            begin
              mem_check[63][7].run()  ;
            end
            begin
              rf_driver[63][7].run()  ;
            end

            begin
              gen[63][8].run()  ;
            end
            begin
              drv[63][8].run()  ;
            end
            begin
              mem_check[63][8].run()  ;
            end
            begin
              rf_driver[63][8].run()  ;
            end

            begin
              gen[63][9].run()  ;
            end
            begin
              drv[63][9].run()  ;
            end
            begin
              mem_check[63][9].run()  ;
            end
            begin
              rf_driver[63][9].run()  ;
            end

            begin
              gen[63][10].run()  ;
            end
            begin
              drv[63][10].run()  ;
            end
            begin
              mem_check[63][10].run()  ;
            end
            begin
              rf_driver[63][10].run()  ;
            end

            begin
              gen[63][11].run()  ;
            end
            begin
              drv[63][11].run()  ;
            end
            begin
              mem_check[63][11].run()  ;
            end
            begin
              rf_driver[63][11].run()  ;
            end

            begin
              gen[63][12].run()  ;
            end
            begin
              drv[63][12].run()  ;
            end
            begin
              mem_check[63][12].run()  ;
            end
            begin
              rf_driver[63][12].run()  ;
            end

            begin
              gen[63][13].run()  ;
            end
            begin
              drv[63][13].run()  ;
            end
            begin
              mem_check[63][13].run()  ;
            end
            begin
              rf_driver[63][13].run()  ;
            end

            begin
              gen[63][14].run()  ;
            end
            begin
              drv[63][14].run()  ;
            end
            begin
              mem_check[63][14].run()  ;
            end
            begin
              rf_driver[63][14].run()  ;
            end

            begin
              gen[63][15].run()  ;
            end
            begin
              drv[63][15].run()  ;
            end
            begin
              mem_check[63][15].run()  ;
            end
            begin
              rf_driver[63][15].run()  ;
            end

            begin
              gen[63][16].run()  ;
            end
            begin
              drv[63][16].run()  ;
            end
            begin
              mem_check[63][16].run()  ;
            end
            begin
              rf_driver[63][16].run()  ;
            end

            begin
              gen[63][17].run()  ;
            end
            begin
              drv[63][17].run()  ;
            end
            begin
              mem_check[63][17].run()  ;
            end
            begin
              rf_driver[63][17].run()  ;
            end

            begin
              gen[63][18].run()  ;
            end
            begin
              drv[63][18].run()  ;
            end
            begin
              mem_check[63][18].run()  ;
            end
            begin
              rf_driver[63][18].run()  ;
            end

            begin
              gen[63][19].run()  ;
            end
            begin
              drv[63][19].run()  ;
            end
            begin
              mem_check[63][19].run()  ;
            end
            begin
              rf_driver[63][19].run()  ;
            end

            begin
              gen[63][20].run()  ;
            end
            begin
              drv[63][20].run()  ;
            end
            begin
              mem_check[63][20].run()  ;
            end
            begin
              rf_driver[63][20].run()  ;
            end

            begin
              gen[63][21].run()  ;
            end
            begin
              drv[63][21].run()  ;
            end
            begin
              mem_check[63][21].run()  ;
            end
            begin
              rf_driver[63][21].run()  ;
            end

            begin
              gen[63][22].run()  ;
            end
            begin
              drv[63][22].run()  ;
            end
            begin
              mem_check[63][22].run()  ;
            end
            begin
              rf_driver[63][22].run()  ;
            end

            begin
              gen[63][23].run()  ;
            end
            begin
              drv[63][23].run()  ;
            end
            begin
              mem_check[63][23].run()  ;
            end
            begin
              rf_driver[63][23].run()  ;
            end

            begin
              gen[63][24].run()  ;
            end
            begin
              drv[63][24].run()  ;
            end
            begin
              mem_check[63][24].run()  ;
            end
            begin
              rf_driver[63][24].run()  ;
            end

            begin
              gen[63][25].run()  ;
            end
            begin
              drv[63][25].run()  ;
            end
            begin
              mem_check[63][25].run()  ;
            end
            begin
              rf_driver[63][25].run()  ;
            end

            begin
              gen[63][26].run()  ;
            end
            begin
              drv[63][26].run()  ;
            end
            begin
              mem_check[63][26].run()  ;
            end
            begin
              rf_driver[63][26].run()  ;
            end

            begin
              gen[63][27].run()  ;
            end
            begin
              drv[63][27].run()  ;
            end
            begin
              mem_check[63][27].run()  ;
            end
            begin
              rf_driver[63][27].run()  ;
            end

            begin
              gen[63][28].run()  ;
            end
            begin
              drv[63][28].run()  ;
            end
            begin
              mem_check[63][28].run()  ;
            end
            begin
              rf_driver[63][28].run()  ;
            end

            begin
              gen[63][29].run()  ;
            end
            begin
              drv[63][29].run()  ;
            end
            begin
              mem_check[63][29].run()  ;
            end
            begin
              rf_driver[63][29].run()  ;
            end

            begin
              gen[63][30].run()  ;
            end
            begin
              drv[63][30].run()  ;
            end
            begin
              mem_check[63][30].run()  ;
            end
            begin
              rf_driver[63][30].run()  ;
            end

            begin
              gen[63][31].run()  ;
            end
            begin
              drv[63][31].run()  ;
            end
            begin
              mem_check[63][31].run()  ;
            end
            begin
              rf_driver[63][31].run()  ;
            end
