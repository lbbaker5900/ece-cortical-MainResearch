
            pe0__stu__valid          ,
            pe0__stu__cntl           ,
            stu__pe0__ready          ,
            pe0__stu__type           ,
            pe0__stu__data           ,
            pe0__stu__oob_data       ,

            pe1__stu__valid          ,
            pe1__stu__cntl           ,
            stu__pe1__ready          ,
            pe1__stu__type           ,
            pe1__stu__data           ,
            pe1__stu__oob_data       ,

            pe2__stu__valid          ,
            pe2__stu__cntl           ,
            stu__pe2__ready          ,
            pe2__stu__type           ,
            pe2__stu__data           ,
            pe2__stu__oob_data       ,

            pe3__stu__valid          ,
            pe3__stu__cntl           ,
            stu__pe3__ready          ,
            pe3__stu__type           ,
            pe3__stu__data           ,
            pe3__stu__oob_data       ,

            pe4__stu__valid          ,
            pe4__stu__cntl           ,
            stu__pe4__ready          ,
            pe4__stu__type           ,
            pe4__stu__data           ,
            pe4__stu__oob_data       ,

            pe5__stu__valid          ,
            pe5__stu__cntl           ,
            stu__pe5__ready          ,
            pe5__stu__type           ,
            pe5__stu__data           ,
            pe5__stu__oob_data       ,

            pe6__stu__valid          ,
            pe6__stu__cntl           ,
            stu__pe6__ready          ,
            pe6__stu__type           ,
            pe6__stu__data           ,
            pe6__stu__oob_data       ,

            pe7__stu__valid          ,
            pe7__stu__cntl           ,
            stu__pe7__ready          ,
            pe7__stu__type           ,
            pe7__stu__data           ,
            pe7__stu__oob_data       ,

            pe8__stu__valid          ,
            pe8__stu__cntl           ,
            stu__pe8__ready          ,
            pe8__stu__type           ,
            pe8__stu__data           ,
            pe8__stu__oob_data       ,

            pe9__stu__valid          ,
            pe9__stu__cntl           ,
            stu__pe9__ready          ,
            pe9__stu__type           ,
            pe9__stu__data           ,
            pe9__stu__oob_data       ,

            pe10__stu__valid          ,
            pe10__stu__cntl           ,
            stu__pe10__ready          ,
            pe10__stu__type           ,
            pe10__stu__data           ,
            pe10__stu__oob_data       ,

            pe11__stu__valid          ,
            pe11__stu__cntl           ,
            stu__pe11__ready          ,
            pe11__stu__type           ,
            pe11__stu__data           ,
            pe11__stu__oob_data       ,

            pe12__stu__valid          ,
            pe12__stu__cntl           ,
            stu__pe12__ready          ,
            pe12__stu__type           ,
            pe12__stu__data           ,
            pe12__stu__oob_data       ,

            pe13__stu__valid          ,
            pe13__stu__cntl           ,
            stu__pe13__ready          ,
            pe13__stu__type           ,
            pe13__stu__data           ,
            pe13__stu__oob_data       ,

            pe14__stu__valid          ,
            pe14__stu__cntl           ,
            stu__pe14__ready          ,
            pe14__stu__type           ,
            pe14__stu__data           ,
            pe14__stu__oob_data       ,

            pe15__stu__valid          ,
            pe15__stu__cntl           ,
            stu__pe15__ready          ,
            pe15__stu__type           ,
            pe15__stu__data           ,
            pe15__stu__oob_data       ,

            pe16__stu__valid          ,
            pe16__stu__cntl           ,
            stu__pe16__ready          ,
            pe16__stu__type           ,
            pe16__stu__data           ,
            pe16__stu__oob_data       ,

            pe17__stu__valid          ,
            pe17__stu__cntl           ,
            stu__pe17__ready          ,
            pe17__stu__type           ,
            pe17__stu__data           ,
            pe17__stu__oob_data       ,

            pe18__stu__valid          ,
            pe18__stu__cntl           ,
            stu__pe18__ready          ,
            pe18__stu__type           ,
            pe18__stu__data           ,
            pe18__stu__oob_data       ,

            pe19__stu__valid          ,
            pe19__stu__cntl           ,
            stu__pe19__ready          ,
            pe19__stu__type           ,
            pe19__stu__data           ,
            pe19__stu__oob_data       ,

            pe20__stu__valid          ,
            pe20__stu__cntl           ,
            stu__pe20__ready          ,
            pe20__stu__type           ,
            pe20__stu__data           ,
            pe20__stu__oob_data       ,

            pe21__stu__valid          ,
            pe21__stu__cntl           ,
            stu__pe21__ready          ,
            pe21__stu__type           ,
            pe21__stu__data           ,
            pe21__stu__oob_data       ,

            pe22__stu__valid          ,
            pe22__stu__cntl           ,
            stu__pe22__ready          ,
            pe22__stu__type           ,
            pe22__stu__data           ,
            pe22__stu__oob_data       ,

            pe23__stu__valid          ,
            pe23__stu__cntl           ,
            stu__pe23__ready          ,
            pe23__stu__type           ,
            pe23__stu__data           ,
            pe23__stu__oob_data       ,

            pe24__stu__valid          ,
            pe24__stu__cntl           ,
            stu__pe24__ready          ,
            pe24__stu__type           ,
            pe24__stu__data           ,
            pe24__stu__oob_data       ,

            pe25__stu__valid          ,
            pe25__stu__cntl           ,
            stu__pe25__ready          ,
            pe25__stu__type           ,
            pe25__stu__data           ,
            pe25__stu__oob_data       ,

            pe26__stu__valid          ,
            pe26__stu__cntl           ,
            stu__pe26__ready          ,
            pe26__stu__type           ,
            pe26__stu__data           ,
            pe26__stu__oob_data       ,

            pe27__stu__valid          ,
            pe27__stu__cntl           ,
            stu__pe27__ready          ,
            pe27__stu__type           ,
            pe27__stu__data           ,
            pe27__stu__oob_data       ,

            pe28__stu__valid          ,
            pe28__stu__cntl           ,
            stu__pe28__ready          ,
            pe28__stu__type           ,
            pe28__stu__data           ,
            pe28__stu__oob_data       ,

            pe29__stu__valid          ,
            pe29__stu__cntl           ,
            stu__pe29__ready          ,
            pe29__stu__type           ,
            pe29__stu__data           ,
            pe29__stu__oob_data       ,

            pe30__stu__valid          ,
            pe30__stu__cntl           ,
            stu__pe30__ready          ,
            pe30__stu__type           ,
            pe30__stu__data           ,
            pe30__stu__oob_data       ,

            pe31__stu__valid          ,
            pe31__stu__cntl           ,
            stu__pe31__ready          ,
            pe31__stu__type           ,
            pe31__stu__data           ,
            pe31__stu__oob_data       ,

            pe32__stu__valid          ,
            pe32__stu__cntl           ,
            stu__pe32__ready          ,
            pe32__stu__type           ,
            pe32__stu__data           ,
            pe32__stu__oob_data       ,

            pe33__stu__valid          ,
            pe33__stu__cntl           ,
            stu__pe33__ready          ,
            pe33__stu__type           ,
            pe33__stu__data           ,
            pe33__stu__oob_data       ,

            pe34__stu__valid          ,
            pe34__stu__cntl           ,
            stu__pe34__ready          ,
            pe34__stu__type           ,
            pe34__stu__data           ,
            pe34__stu__oob_data       ,

            pe35__stu__valid          ,
            pe35__stu__cntl           ,
            stu__pe35__ready          ,
            pe35__stu__type           ,
            pe35__stu__data           ,
            pe35__stu__oob_data       ,

            pe36__stu__valid          ,
            pe36__stu__cntl           ,
            stu__pe36__ready          ,
            pe36__stu__type           ,
            pe36__stu__data           ,
            pe36__stu__oob_data       ,

            pe37__stu__valid          ,
            pe37__stu__cntl           ,
            stu__pe37__ready          ,
            pe37__stu__type           ,
            pe37__stu__data           ,
            pe37__stu__oob_data       ,

            pe38__stu__valid          ,
            pe38__stu__cntl           ,
            stu__pe38__ready          ,
            pe38__stu__type           ,
            pe38__stu__data           ,
            pe38__stu__oob_data       ,

            pe39__stu__valid          ,
            pe39__stu__cntl           ,
            stu__pe39__ready          ,
            pe39__stu__type           ,
            pe39__stu__data           ,
            pe39__stu__oob_data       ,

            pe40__stu__valid          ,
            pe40__stu__cntl           ,
            stu__pe40__ready          ,
            pe40__stu__type           ,
            pe40__stu__data           ,
            pe40__stu__oob_data       ,

            pe41__stu__valid          ,
            pe41__stu__cntl           ,
            stu__pe41__ready          ,
            pe41__stu__type           ,
            pe41__stu__data           ,
            pe41__stu__oob_data       ,

            pe42__stu__valid          ,
            pe42__stu__cntl           ,
            stu__pe42__ready          ,
            pe42__stu__type           ,
            pe42__stu__data           ,
            pe42__stu__oob_data       ,

            pe43__stu__valid          ,
            pe43__stu__cntl           ,
            stu__pe43__ready          ,
            pe43__stu__type           ,
            pe43__stu__data           ,
            pe43__stu__oob_data       ,

            pe44__stu__valid          ,
            pe44__stu__cntl           ,
            stu__pe44__ready          ,
            pe44__stu__type           ,
            pe44__stu__data           ,
            pe44__stu__oob_data       ,

            pe45__stu__valid          ,
            pe45__stu__cntl           ,
            stu__pe45__ready          ,
            pe45__stu__type           ,
            pe45__stu__data           ,
            pe45__stu__oob_data       ,

            pe46__stu__valid          ,
            pe46__stu__cntl           ,
            stu__pe46__ready          ,
            pe46__stu__type           ,
            pe46__stu__data           ,
            pe46__stu__oob_data       ,

            pe47__stu__valid          ,
            pe47__stu__cntl           ,
            stu__pe47__ready          ,
            pe47__stu__type           ,
            pe47__stu__data           ,
            pe47__stu__oob_data       ,

            pe48__stu__valid          ,
            pe48__stu__cntl           ,
            stu__pe48__ready          ,
            pe48__stu__type           ,
            pe48__stu__data           ,
            pe48__stu__oob_data       ,

            pe49__stu__valid          ,
            pe49__stu__cntl           ,
            stu__pe49__ready          ,
            pe49__stu__type           ,
            pe49__stu__data           ,
            pe49__stu__oob_data       ,

            pe50__stu__valid          ,
            pe50__stu__cntl           ,
            stu__pe50__ready          ,
            pe50__stu__type           ,
            pe50__stu__data           ,
            pe50__stu__oob_data       ,

            pe51__stu__valid          ,
            pe51__stu__cntl           ,
            stu__pe51__ready          ,
            pe51__stu__type           ,
            pe51__stu__data           ,
            pe51__stu__oob_data       ,

            pe52__stu__valid          ,
            pe52__stu__cntl           ,
            stu__pe52__ready          ,
            pe52__stu__type           ,
            pe52__stu__data           ,
            pe52__stu__oob_data       ,

            pe53__stu__valid          ,
            pe53__stu__cntl           ,
            stu__pe53__ready          ,
            pe53__stu__type           ,
            pe53__stu__data           ,
            pe53__stu__oob_data       ,

            pe54__stu__valid          ,
            pe54__stu__cntl           ,
            stu__pe54__ready          ,
            pe54__stu__type           ,
            pe54__stu__data           ,
            pe54__stu__oob_data       ,

            pe55__stu__valid          ,
            pe55__stu__cntl           ,
            stu__pe55__ready          ,
            pe55__stu__type           ,
            pe55__stu__data           ,
            pe55__stu__oob_data       ,

            pe56__stu__valid          ,
            pe56__stu__cntl           ,
            stu__pe56__ready          ,
            pe56__stu__type           ,
            pe56__stu__data           ,
            pe56__stu__oob_data       ,

            pe57__stu__valid          ,
            pe57__stu__cntl           ,
            stu__pe57__ready          ,
            pe57__stu__type           ,
            pe57__stu__data           ,
            pe57__stu__oob_data       ,

            pe58__stu__valid          ,
            pe58__stu__cntl           ,
            stu__pe58__ready          ,
            pe58__stu__type           ,
            pe58__stu__data           ,
            pe58__stu__oob_data       ,

            pe59__stu__valid          ,
            pe59__stu__cntl           ,
            stu__pe59__ready          ,
            pe59__stu__type           ,
            pe59__stu__data           ,
            pe59__stu__oob_data       ,

            pe60__stu__valid          ,
            pe60__stu__cntl           ,
            stu__pe60__ready          ,
            pe60__stu__type           ,
            pe60__stu__data           ,
            pe60__stu__oob_data       ,

            pe61__stu__valid          ,
            pe61__stu__cntl           ,
            stu__pe61__ready          ,
            pe61__stu__type           ,
            pe61__stu__data           ,
            pe61__stu__oob_data       ,

            pe62__stu__valid          ,
            pe62__stu__cntl           ,
            stu__pe62__ready          ,
            pe62__stu__type           ,
            pe62__stu__data           ,
            pe62__stu__oob_data       ,

            pe63__stu__valid          ,
            pe63__stu__cntl           ,
            stu__pe63__ready          ,
            pe63__stu__type           ,
            pe63__stu__data           ,
            pe63__stu__oob_data       ,

