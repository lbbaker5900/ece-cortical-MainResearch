
  assign reg__scntl__lane0_ready  = 1'b1          ;
  assign reg__scntl__lane1_ready  = 1'b1          ;
  assign reg__scntl__lane2_ready  = 1'b1          ;
  assign reg__scntl__lane3_ready  = 1'b1          ;
  assign reg__scntl__lane4_ready  = 1'b1          ;
  assign reg__scntl__lane5_ready  = 1'b1          ;
  assign reg__scntl__lane6_ready  = 1'b1          ;
  assign reg__scntl__lane7_ready  = 1'b1          ;
  assign reg__scntl__lane8_ready  = 1'b1          ;
  assign reg__scntl__lane9_ready  = 1'b1          ;
  assign reg__scntl__lane10_ready  = 1'b1          ;
  assign reg__scntl__lane11_ready  = 1'b1          ;
  assign reg__scntl__lane12_ready  = 1'b1          ;
  assign reg__scntl__lane13_ready  = 1'b1          ;
  assign reg__scntl__lane14_ready  = 1'b1          ;
  assign reg__scntl__lane15_ready  = 1'b1          ;
  assign reg__scntl__lane16_ready  = 1'b1          ;
  assign reg__scntl__lane17_ready  = 1'b1          ;
  assign reg__scntl__lane18_ready  = 1'b1          ;
  assign reg__scntl__lane19_ready  = 1'b1          ;
  assign reg__scntl__lane20_ready  = 1'b1          ;
  assign reg__scntl__lane21_ready  = 1'b1          ;
  assign reg__scntl__lane22_ready  = 1'b1          ;
  assign reg__scntl__lane23_ready  = 1'b1          ;
  assign reg__scntl__lane24_ready  = 1'b1          ;
  assign reg__scntl__lane25_ready  = 1'b1          ;
  assign reg__scntl__lane26_ready  = 1'b1          ;
  assign reg__scntl__lane27_ready  = 1'b1          ;
  assign reg__scntl__lane28_ready  = 1'b1          ;
  assign reg__scntl__lane29_ready  = 1'b1          ;
  assign reg__scntl__lane30_ready  = 1'b1          ;
  assign reg__scntl__lane31_ready  = 1'b1          ;
