
  wire                                    reg__scntl__lane0_ready    ;
  wire                                    scntl__reg__lane0_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane0_data     ;
  wire                                    reg__scntl__lane1_ready    ;
  wire                                    scntl__reg__lane1_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane1_data     ;
  wire                                    reg__scntl__lane2_ready    ;
  wire                                    scntl__reg__lane2_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane2_data     ;
  wire                                    reg__scntl__lane3_ready    ;
  wire                                    scntl__reg__lane3_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane3_data     ;
  wire                                    reg__scntl__lane4_ready    ;
  wire                                    scntl__reg__lane4_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane4_data     ;
  wire                                    reg__scntl__lane5_ready    ;
  wire                                    scntl__reg__lane5_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane5_data     ;
  wire                                    reg__scntl__lane6_ready    ;
  wire                                    scntl__reg__lane6_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane6_data     ;
  wire                                    reg__scntl__lane7_ready    ;
  wire                                    scntl__reg__lane7_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane7_data     ;
  wire                                    reg__scntl__lane8_ready    ;
  wire                                    scntl__reg__lane8_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane8_data     ;
  wire                                    reg__scntl__lane9_ready    ;
  wire                                    scntl__reg__lane9_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane9_data     ;
  wire                                    reg__scntl__lane10_ready    ;
  wire                                    scntl__reg__lane10_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane10_data     ;
  wire                                    reg__scntl__lane11_ready    ;
  wire                                    scntl__reg__lane11_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane11_data     ;
  wire                                    reg__scntl__lane12_ready    ;
  wire                                    scntl__reg__lane12_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane12_data     ;
  wire                                    reg__scntl__lane13_ready    ;
  wire                                    scntl__reg__lane13_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane13_data     ;
  wire                                    reg__scntl__lane14_ready    ;
  wire                                    scntl__reg__lane14_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane14_data     ;
  wire                                    reg__scntl__lane15_ready    ;
  wire                                    scntl__reg__lane15_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane15_data     ;
  wire                                    reg__scntl__lane16_ready    ;
  wire                                    scntl__reg__lane16_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane16_data     ;
  wire                                    reg__scntl__lane17_ready    ;
  wire                                    scntl__reg__lane17_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane17_data     ;
  wire                                    reg__scntl__lane18_ready    ;
  wire                                    scntl__reg__lane18_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane18_data     ;
  wire                                    reg__scntl__lane19_ready    ;
  wire                                    scntl__reg__lane19_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane19_data     ;
  wire                                    reg__scntl__lane20_ready    ;
  wire                                    scntl__reg__lane20_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane20_data     ;
  wire                                    reg__scntl__lane21_ready    ;
  wire                                    scntl__reg__lane21_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane21_data     ;
  wire                                    reg__scntl__lane22_ready    ;
  wire                                    scntl__reg__lane22_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane22_data     ;
  wire                                    reg__scntl__lane23_ready    ;
  wire                                    scntl__reg__lane23_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane23_data     ;
  wire                                    reg__scntl__lane24_ready    ;
  wire                                    scntl__reg__lane24_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane24_data     ;
  wire                                    reg__scntl__lane25_ready    ;
  wire                                    scntl__reg__lane25_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane25_data     ;
  wire                                    reg__scntl__lane26_ready    ;
  wire                                    scntl__reg__lane26_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane26_data     ;
  wire                                    reg__scntl__lane27_ready    ;
  wire                                    scntl__reg__lane27_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane27_data     ;
  wire                                    reg__scntl__lane28_ready    ;
  wire                                    scntl__reg__lane28_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane28_data     ;
  wire                                    reg__scntl__lane29_ready    ;
  wire                                    scntl__reg__lane29_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane29_data     ;
  wire                                    reg__scntl__lane30_ready    ;
  wire                                    scntl__reg__lane30_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane30_data     ;
  wire                                    reg__scntl__lane31_ready    ;
  wire                                    scntl__reg__lane31_valid    ;
  wire   [`STREAMING_OP_RESULT_RANGE   ]  scntl__reg__lane31_data     ;
