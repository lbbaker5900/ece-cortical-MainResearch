
            pe0__stu__valid          ,
            pe0__stu__cntl           ,
            stu__pe0__ready          ,
            pe0__stu__type           ,
            pe0__stu__data           ,
            pe0__stu__oob_data       ,

            pe1__stu__valid          ,
            pe1__stu__cntl           ,
            stu__pe1__ready          ,
            pe1__stu__type           ,
            pe1__stu__data           ,
            pe1__stu__oob_data       ,

            pe2__stu__valid          ,
            pe2__stu__cntl           ,
            stu__pe2__ready          ,
            pe2__stu__type           ,
            pe2__stu__data           ,
            pe2__stu__oob_data       ,

            pe3__stu__valid          ,
            pe3__stu__cntl           ,
            stu__pe3__ready          ,
            pe3__stu__type           ,
            pe3__stu__data           ,
            pe3__stu__oob_data       ,

