
               // PE 0, Lane 0                 
               .pe0__std__lane0_strm0_ready         ( pe0__std__lane0_strm0_ready      ),      
               .std__pe0__lane0_strm0_cntl          ( std__pe0__lane0_strm0_cntl       ),      
               .std__pe0__lane0_strm0_data          ( std__pe0__lane0_strm0_data       ),      
               .std__pe0__lane0_strm0_data_valid    ( std__pe0__lane0_strm0_data_valid ),      
               .std__pe0__lane0_strm0_data_mask     ( std__pe0__lane0_strm0_data_mask  ),      

               .pe0__std__lane0_strm1_ready         ( pe0__std__lane0_strm1_ready      ),      
               .std__pe0__lane0_strm1_cntl          ( std__pe0__lane0_strm1_cntl       ),      
               .std__pe0__lane0_strm1_data          ( std__pe0__lane0_strm1_data       ),      
               .std__pe0__lane0_strm1_data_valid    ( std__pe0__lane0_strm1_data_valid ),      
               .std__pe0__lane0_strm1_data_mask     ( std__pe0__lane0_strm1_data_mask  ),      

               // PE 0, Lane 1                 
               .pe0__std__lane1_strm0_ready         ( pe0__std__lane1_strm0_ready      ),      
               .std__pe0__lane1_strm0_cntl          ( std__pe0__lane1_strm0_cntl       ),      
               .std__pe0__lane1_strm0_data          ( std__pe0__lane1_strm0_data       ),      
               .std__pe0__lane1_strm0_data_valid    ( std__pe0__lane1_strm0_data_valid ),      
               .std__pe0__lane1_strm0_data_mask     ( std__pe0__lane1_strm0_data_mask  ),      

               .pe0__std__lane1_strm1_ready         ( pe0__std__lane1_strm1_ready      ),      
               .std__pe0__lane1_strm1_cntl          ( std__pe0__lane1_strm1_cntl       ),      
               .std__pe0__lane1_strm1_data          ( std__pe0__lane1_strm1_data       ),      
               .std__pe0__lane1_strm1_data_valid    ( std__pe0__lane1_strm1_data_valid ),      
               .std__pe0__lane1_strm1_data_mask     ( std__pe0__lane1_strm1_data_mask  ),      

               // PE 0, Lane 2                 
               .pe0__std__lane2_strm0_ready         ( pe0__std__lane2_strm0_ready      ),      
               .std__pe0__lane2_strm0_cntl          ( std__pe0__lane2_strm0_cntl       ),      
               .std__pe0__lane2_strm0_data          ( std__pe0__lane2_strm0_data       ),      
               .std__pe0__lane2_strm0_data_valid    ( std__pe0__lane2_strm0_data_valid ),      
               .std__pe0__lane2_strm0_data_mask     ( std__pe0__lane2_strm0_data_mask  ),      

               .pe0__std__lane2_strm1_ready         ( pe0__std__lane2_strm1_ready      ),      
               .std__pe0__lane2_strm1_cntl          ( std__pe0__lane2_strm1_cntl       ),      
               .std__pe0__lane2_strm1_data          ( std__pe0__lane2_strm1_data       ),      
               .std__pe0__lane2_strm1_data_valid    ( std__pe0__lane2_strm1_data_valid ),      
               .std__pe0__lane2_strm1_data_mask     ( std__pe0__lane2_strm1_data_mask  ),      

               // PE 0, Lane 3                 
               .pe0__std__lane3_strm0_ready         ( pe0__std__lane3_strm0_ready      ),      
               .std__pe0__lane3_strm0_cntl          ( std__pe0__lane3_strm0_cntl       ),      
               .std__pe0__lane3_strm0_data          ( std__pe0__lane3_strm0_data       ),      
               .std__pe0__lane3_strm0_data_valid    ( std__pe0__lane3_strm0_data_valid ),      
               .std__pe0__lane3_strm0_data_mask     ( std__pe0__lane3_strm0_data_mask  ),      

               .pe0__std__lane3_strm1_ready         ( pe0__std__lane3_strm1_ready      ),      
               .std__pe0__lane3_strm1_cntl          ( std__pe0__lane3_strm1_cntl       ),      
               .std__pe0__lane3_strm1_data          ( std__pe0__lane3_strm1_data       ),      
               .std__pe0__lane3_strm1_data_valid    ( std__pe0__lane3_strm1_data_valid ),      
               .std__pe0__lane3_strm1_data_mask     ( std__pe0__lane3_strm1_data_mask  ),      

               // PE 0, Lane 4                 
               .pe0__std__lane4_strm0_ready         ( pe0__std__lane4_strm0_ready      ),      
               .std__pe0__lane4_strm0_cntl          ( std__pe0__lane4_strm0_cntl       ),      
               .std__pe0__lane4_strm0_data          ( std__pe0__lane4_strm0_data       ),      
               .std__pe0__lane4_strm0_data_valid    ( std__pe0__lane4_strm0_data_valid ),      
               .std__pe0__lane4_strm0_data_mask     ( std__pe0__lane4_strm0_data_mask  ),      

               .pe0__std__lane4_strm1_ready         ( pe0__std__lane4_strm1_ready      ),      
               .std__pe0__lane4_strm1_cntl          ( std__pe0__lane4_strm1_cntl       ),      
               .std__pe0__lane4_strm1_data          ( std__pe0__lane4_strm1_data       ),      
               .std__pe0__lane4_strm1_data_valid    ( std__pe0__lane4_strm1_data_valid ),      
               .std__pe0__lane4_strm1_data_mask     ( std__pe0__lane4_strm1_data_mask  ),      

               // PE 0, Lane 5                 
               .pe0__std__lane5_strm0_ready         ( pe0__std__lane5_strm0_ready      ),      
               .std__pe0__lane5_strm0_cntl          ( std__pe0__lane5_strm0_cntl       ),      
               .std__pe0__lane5_strm0_data          ( std__pe0__lane5_strm0_data       ),      
               .std__pe0__lane5_strm0_data_valid    ( std__pe0__lane5_strm0_data_valid ),      
               .std__pe0__lane5_strm0_data_mask     ( std__pe0__lane5_strm0_data_mask  ),      

               .pe0__std__lane5_strm1_ready         ( pe0__std__lane5_strm1_ready      ),      
               .std__pe0__lane5_strm1_cntl          ( std__pe0__lane5_strm1_cntl       ),      
               .std__pe0__lane5_strm1_data          ( std__pe0__lane5_strm1_data       ),      
               .std__pe0__lane5_strm1_data_valid    ( std__pe0__lane5_strm1_data_valid ),      
               .std__pe0__lane5_strm1_data_mask     ( std__pe0__lane5_strm1_data_mask  ),      

               // PE 0, Lane 6                 
               .pe0__std__lane6_strm0_ready         ( pe0__std__lane6_strm0_ready      ),      
               .std__pe0__lane6_strm0_cntl          ( std__pe0__lane6_strm0_cntl       ),      
               .std__pe0__lane6_strm0_data          ( std__pe0__lane6_strm0_data       ),      
               .std__pe0__lane6_strm0_data_valid    ( std__pe0__lane6_strm0_data_valid ),      
               .std__pe0__lane6_strm0_data_mask     ( std__pe0__lane6_strm0_data_mask  ),      

               .pe0__std__lane6_strm1_ready         ( pe0__std__lane6_strm1_ready      ),      
               .std__pe0__lane6_strm1_cntl          ( std__pe0__lane6_strm1_cntl       ),      
               .std__pe0__lane6_strm1_data          ( std__pe0__lane6_strm1_data       ),      
               .std__pe0__lane6_strm1_data_valid    ( std__pe0__lane6_strm1_data_valid ),      
               .std__pe0__lane6_strm1_data_mask     ( std__pe0__lane6_strm1_data_mask  ),      

               // PE 0, Lane 7                 
               .pe0__std__lane7_strm0_ready         ( pe0__std__lane7_strm0_ready      ),      
               .std__pe0__lane7_strm0_cntl          ( std__pe0__lane7_strm0_cntl       ),      
               .std__pe0__lane7_strm0_data          ( std__pe0__lane7_strm0_data       ),      
               .std__pe0__lane7_strm0_data_valid    ( std__pe0__lane7_strm0_data_valid ),      
               .std__pe0__lane7_strm0_data_mask     ( std__pe0__lane7_strm0_data_mask  ),      

               .pe0__std__lane7_strm1_ready         ( pe0__std__lane7_strm1_ready      ),      
               .std__pe0__lane7_strm1_cntl          ( std__pe0__lane7_strm1_cntl       ),      
               .std__pe0__lane7_strm1_data          ( std__pe0__lane7_strm1_data       ),      
               .std__pe0__lane7_strm1_data_valid    ( std__pe0__lane7_strm1_data_valid ),      
               .std__pe0__lane7_strm1_data_mask     ( std__pe0__lane7_strm1_data_mask  ),      

               // PE 0, Lane 8                 
               .pe0__std__lane8_strm0_ready         ( pe0__std__lane8_strm0_ready      ),      
               .std__pe0__lane8_strm0_cntl          ( std__pe0__lane8_strm0_cntl       ),      
               .std__pe0__lane8_strm0_data          ( std__pe0__lane8_strm0_data       ),      
               .std__pe0__lane8_strm0_data_valid    ( std__pe0__lane8_strm0_data_valid ),      
               .std__pe0__lane8_strm0_data_mask     ( std__pe0__lane8_strm0_data_mask  ),      

               .pe0__std__lane8_strm1_ready         ( pe0__std__lane8_strm1_ready      ),      
               .std__pe0__lane8_strm1_cntl          ( std__pe0__lane8_strm1_cntl       ),      
               .std__pe0__lane8_strm1_data          ( std__pe0__lane8_strm1_data       ),      
               .std__pe0__lane8_strm1_data_valid    ( std__pe0__lane8_strm1_data_valid ),      
               .std__pe0__lane8_strm1_data_mask     ( std__pe0__lane8_strm1_data_mask  ),      

               // PE 0, Lane 9                 
               .pe0__std__lane9_strm0_ready         ( pe0__std__lane9_strm0_ready      ),      
               .std__pe0__lane9_strm0_cntl          ( std__pe0__lane9_strm0_cntl       ),      
               .std__pe0__lane9_strm0_data          ( std__pe0__lane9_strm0_data       ),      
               .std__pe0__lane9_strm0_data_valid    ( std__pe0__lane9_strm0_data_valid ),      
               .std__pe0__lane9_strm0_data_mask     ( std__pe0__lane9_strm0_data_mask  ),      

               .pe0__std__lane9_strm1_ready         ( pe0__std__lane9_strm1_ready      ),      
               .std__pe0__lane9_strm1_cntl          ( std__pe0__lane9_strm1_cntl       ),      
               .std__pe0__lane9_strm1_data          ( std__pe0__lane9_strm1_data       ),      
               .std__pe0__lane9_strm1_data_valid    ( std__pe0__lane9_strm1_data_valid ),      
               .std__pe0__lane9_strm1_data_mask     ( std__pe0__lane9_strm1_data_mask  ),      

               // PE 0, Lane 10                 
               .pe0__std__lane10_strm0_ready         ( pe0__std__lane10_strm0_ready      ),      
               .std__pe0__lane10_strm0_cntl          ( std__pe0__lane10_strm0_cntl       ),      
               .std__pe0__lane10_strm0_data          ( std__pe0__lane10_strm0_data       ),      
               .std__pe0__lane10_strm0_data_valid    ( std__pe0__lane10_strm0_data_valid ),      
               .std__pe0__lane10_strm0_data_mask     ( std__pe0__lane10_strm0_data_mask  ),      

               .pe0__std__lane10_strm1_ready         ( pe0__std__lane10_strm1_ready      ),      
               .std__pe0__lane10_strm1_cntl          ( std__pe0__lane10_strm1_cntl       ),      
               .std__pe0__lane10_strm1_data          ( std__pe0__lane10_strm1_data       ),      
               .std__pe0__lane10_strm1_data_valid    ( std__pe0__lane10_strm1_data_valid ),      
               .std__pe0__lane10_strm1_data_mask     ( std__pe0__lane10_strm1_data_mask  ),      

               // PE 0, Lane 11                 
               .pe0__std__lane11_strm0_ready         ( pe0__std__lane11_strm0_ready      ),      
               .std__pe0__lane11_strm0_cntl          ( std__pe0__lane11_strm0_cntl       ),      
               .std__pe0__lane11_strm0_data          ( std__pe0__lane11_strm0_data       ),      
               .std__pe0__lane11_strm0_data_valid    ( std__pe0__lane11_strm0_data_valid ),      
               .std__pe0__lane11_strm0_data_mask     ( std__pe0__lane11_strm0_data_mask  ),      

               .pe0__std__lane11_strm1_ready         ( pe0__std__lane11_strm1_ready      ),      
               .std__pe0__lane11_strm1_cntl          ( std__pe0__lane11_strm1_cntl       ),      
               .std__pe0__lane11_strm1_data          ( std__pe0__lane11_strm1_data       ),      
               .std__pe0__lane11_strm1_data_valid    ( std__pe0__lane11_strm1_data_valid ),      
               .std__pe0__lane11_strm1_data_mask     ( std__pe0__lane11_strm1_data_mask  ),      

               // PE 0, Lane 12                 
               .pe0__std__lane12_strm0_ready         ( pe0__std__lane12_strm0_ready      ),      
               .std__pe0__lane12_strm0_cntl          ( std__pe0__lane12_strm0_cntl       ),      
               .std__pe0__lane12_strm0_data          ( std__pe0__lane12_strm0_data       ),      
               .std__pe0__lane12_strm0_data_valid    ( std__pe0__lane12_strm0_data_valid ),      
               .std__pe0__lane12_strm0_data_mask     ( std__pe0__lane12_strm0_data_mask  ),      

               .pe0__std__lane12_strm1_ready         ( pe0__std__lane12_strm1_ready      ),      
               .std__pe0__lane12_strm1_cntl          ( std__pe0__lane12_strm1_cntl       ),      
               .std__pe0__lane12_strm1_data          ( std__pe0__lane12_strm1_data       ),      
               .std__pe0__lane12_strm1_data_valid    ( std__pe0__lane12_strm1_data_valid ),      
               .std__pe0__lane12_strm1_data_mask     ( std__pe0__lane12_strm1_data_mask  ),      

               // PE 0, Lane 13                 
               .pe0__std__lane13_strm0_ready         ( pe0__std__lane13_strm0_ready      ),      
               .std__pe0__lane13_strm0_cntl          ( std__pe0__lane13_strm0_cntl       ),      
               .std__pe0__lane13_strm0_data          ( std__pe0__lane13_strm0_data       ),      
               .std__pe0__lane13_strm0_data_valid    ( std__pe0__lane13_strm0_data_valid ),      
               .std__pe0__lane13_strm0_data_mask     ( std__pe0__lane13_strm0_data_mask  ),      

               .pe0__std__lane13_strm1_ready         ( pe0__std__lane13_strm1_ready      ),      
               .std__pe0__lane13_strm1_cntl          ( std__pe0__lane13_strm1_cntl       ),      
               .std__pe0__lane13_strm1_data          ( std__pe0__lane13_strm1_data       ),      
               .std__pe0__lane13_strm1_data_valid    ( std__pe0__lane13_strm1_data_valid ),      
               .std__pe0__lane13_strm1_data_mask     ( std__pe0__lane13_strm1_data_mask  ),      

               // PE 0, Lane 14                 
               .pe0__std__lane14_strm0_ready         ( pe0__std__lane14_strm0_ready      ),      
               .std__pe0__lane14_strm0_cntl          ( std__pe0__lane14_strm0_cntl       ),      
               .std__pe0__lane14_strm0_data          ( std__pe0__lane14_strm0_data       ),      
               .std__pe0__lane14_strm0_data_valid    ( std__pe0__lane14_strm0_data_valid ),      
               .std__pe0__lane14_strm0_data_mask     ( std__pe0__lane14_strm0_data_mask  ),      

               .pe0__std__lane14_strm1_ready         ( pe0__std__lane14_strm1_ready      ),      
               .std__pe0__lane14_strm1_cntl          ( std__pe0__lane14_strm1_cntl       ),      
               .std__pe0__lane14_strm1_data          ( std__pe0__lane14_strm1_data       ),      
               .std__pe0__lane14_strm1_data_valid    ( std__pe0__lane14_strm1_data_valid ),      
               .std__pe0__lane14_strm1_data_mask     ( std__pe0__lane14_strm1_data_mask  ),      

               // PE 0, Lane 15                 
               .pe0__std__lane15_strm0_ready         ( pe0__std__lane15_strm0_ready      ),      
               .std__pe0__lane15_strm0_cntl          ( std__pe0__lane15_strm0_cntl       ),      
               .std__pe0__lane15_strm0_data          ( std__pe0__lane15_strm0_data       ),      
               .std__pe0__lane15_strm0_data_valid    ( std__pe0__lane15_strm0_data_valid ),      
               .std__pe0__lane15_strm0_data_mask     ( std__pe0__lane15_strm0_data_mask  ),      

               .pe0__std__lane15_strm1_ready         ( pe0__std__lane15_strm1_ready      ),      
               .std__pe0__lane15_strm1_cntl          ( std__pe0__lane15_strm1_cntl       ),      
               .std__pe0__lane15_strm1_data          ( std__pe0__lane15_strm1_data       ),      
               .std__pe0__lane15_strm1_data_valid    ( std__pe0__lane15_strm1_data_valid ),      
               .std__pe0__lane15_strm1_data_mask     ( std__pe0__lane15_strm1_data_mask  ),      

               // PE 0, Lane 16                 
               .pe0__std__lane16_strm0_ready         ( pe0__std__lane16_strm0_ready      ),      
               .std__pe0__lane16_strm0_cntl          ( std__pe0__lane16_strm0_cntl       ),      
               .std__pe0__lane16_strm0_data          ( std__pe0__lane16_strm0_data       ),      
               .std__pe0__lane16_strm0_data_valid    ( std__pe0__lane16_strm0_data_valid ),      
               .std__pe0__lane16_strm0_data_mask     ( std__pe0__lane16_strm0_data_mask  ),      

               .pe0__std__lane16_strm1_ready         ( pe0__std__lane16_strm1_ready      ),      
               .std__pe0__lane16_strm1_cntl          ( std__pe0__lane16_strm1_cntl       ),      
               .std__pe0__lane16_strm1_data          ( std__pe0__lane16_strm1_data       ),      
               .std__pe0__lane16_strm1_data_valid    ( std__pe0__lane16_strm1_data_valid ),      
               .std__pe0__lane16_strm1_data_mask     ( std__pe0__lane16_strm1_data_mask  ),      

               // PE 0, Lane 17                 
               .pe0__std__lane17_strm0_ready         ( pe0__std__lane17_strm0_ready      ),      
               .std__pe0__lane17_strm0_cntl          ( std__pe0__lane17_strm0_cntl       ),      
               .std__pe0__lane17_strm0_data          ( std__pe0__lane17_strm0_data       ),      
               .std__pe0__lane17_strm0_data_valid    ( std__pe0__lane17_strm0_data_valid ),      
               .std__pe0__lane17_strm0_data_mask     ( std__pe0__lane17_strm0_data_mask  ),      

               .pe0__std__lane17_strm1_ready         ( pe0__std__lane17_strm1_ready      ),      
               .std__pe0__lane17_strm1_cntl          ( std__pe0__lane17_strm1_cntl       ),      
               .std__pe0__lane17_strm1_data          ( std__pe0__lane17_strm1_data       ),      
               .std__pe0__lane17_strm1_data_valid    ( std__pe0__lane17_strm1_data_valid ),      
               .std__pe0__lane17_strm1_data_mask     ( std__pe0__lane17_strm1_data_mask  ),      

               // PE 0, Lane 18                 
               .pe0__std__lane18_strm0_ready         ( pe0__std__lane18_strm0_ready      ),      
               .std__pe0__lane18_strm0_cntl          ( std__pe0__lane18_strm0_cntl       ),      
               .std__pe0__lane18_strm0_data          ( std__pe0__lane18_strm0_data       ),      
               .std__pe0__lane18_strm0_data_valid    ( std__pe0__lane18_strm0_data_valid ),      
               .std__pe0__lane18_strm0_data_mask     ( std__pe0__lane18_strm0_data_mask  ),      

               .pe0__std__lane18_strm1_ready         ( pe0__std__lane18_strm1_ready      ),      
               .std__pe0__lane18_strm1_cntl          ( std__pe0__lane18_strm1_cntl       ),      
               .std__pe0__lane18_strm1_data          ( std__pe0__lane18_strm1_data       ),      
               .std__pe0__lane18_strm1_data_valid    ( std__pe0__lane18_strm1_data_valid ),      
               .std__pe0__lane18_strm1_data_mask     ( std__pe0__lane18_strm1_data_mask  ),      

               // PE 0, Lane 19                 
               .pe0__std__lane19_strm0_ready         ( pe0__std__lane19_strm0_ready      ),      
               .std__pe0__lane19_strm0_cntl          ( std__pe0__lane19_strm0_cntl       ),      
               .std__pe0__lane19_strm0_data          ( std__pe0__lane19_strm0_data       ),      
               .std__pe0__lane19_strm0_data_valid    ( std__pe0__lane19_strm0_data_valid ),      
               .std__pe0__lane19_strm0_data_mask     ( std__pe0__lane19_strm0_data_mask  ),      

               .pe0__std__lane19_strm1_ready         ( pe0__std__lane19_strm1_ready      ),      
               .std__pe0__lane19_strm1_cntl          ( std__pe0__lane19_strm1_cntl       ),      
               .std__pe0__lane19_strm1_data          ( std__pe0__lane19_strm1_data       ),      
               .std__pe0__lane19_strm1_data_valid    ( std__pe0__lane19_strm1_data_valid ),      
               .std__pe0__lane19_strm1_data_mask     ( std__pe0__lane19_strm1_data_mask  ),      

               // PE 0, Lane 20                 
               .pe0__std__lane20_strm0_ready         ( pe0__std__lane20_strm0_ready      ),      
               .std__pe0__lane20_strm0_cntl          ( std__pe0__lane20_strm0_cntl       ),      
               .std__pe0__lane20_strm0_data          ( std__pe0__lane20_strm0_data       ),      
               .std__pe0__lane20_strm0_data_valid    ( std__pe0__lane20_strm0_data_valid ),      
               .std__pe0__lane20_strm0_data_mask     ( std__pe0__lane20_strm0_data_mask  ),      

               .pe0__std__lane20_strm1_ready         ( pe0__std__lane20_strm1_ready      ),      
               .std__pe0__lane20_strm1_cntl          ( std__pe0__lane20_strm1_cntl       ),      
               .std__pe0__lane20_strm1_data          ( std__pe0__lane20_strm1_data       ),      
               .std__pe0__lane20_strm1_data_valid    ( std__pe0__lane20_strm1_data_valid ),      
               .std__pe0__lane20_strm1_data_mask     ( std__pe0__lane20_strm1_data_mask  ),      

               // PE 0, Lane 21                 
               .pe0__std__lane21_strm0_ready         ( pe0__std__lane21_strm0_ready      ),      
               .std__pe0__lane21_strm0_cntl          ( std__pe0__lane21_strm0_cntl       ),      
               .std__pe0__lane21_strm0_data          ( std__pe0__lane21_strm0_data       ),      
               .std__pe0__lane21_strm0_data_valid    ( std__pe0__lane21_strm0_data_valid ),      
               .std__pe0__lane21_strm0_data_mask     ( std__pe0__lane21_strm0_data_mask  ),      

               .pe0__std__lane21_strm1_ready         ( pe0__std__lane21_strm1_ready      ),      
               .std__pe0__lane21_strm1_cntl          ( std__pe0__lane21_strm1_cntl       ),      
               .std__pe0__lane21_strm1_data          ( std__pe0__lane21_strm1_data       ),      
               .std__pe0__lane21_strm1_data_valid    ( std__pe0__lane21_strm1_data_valid ),      
               .std__pe0__lane21_strm1_data_mask     ( std__pe0__lane21_strm1_data_mask  ),      

               // PE 0, Lane 22                 
               .pe0__std__lane22_strm0_ready         ( pe0__std__lane22_strm0_ready      ),      
               .std__pe0__lane22_strm0_cntl          ( std__pe0__lane22_strm0_cntl       ),      
               .std__pe0__lane22_strm0_data          ( std__pe0__lane22_strm0_data       ),      
               .std__pe0__lane22_strm0_data_valid    ( std__pe0__lane22_strm0_data_valid ),      
               .std__pe0__lane22_strm0_data_mask     ( std__pe0__lane22_strm0_data_mask  ),      

               .pe0__std__lane22_strm1_ready         ( pe0__std__lane22_strm1_ready      ),      
               .std__pe0__lane22_strm1_cntl          ( std__pe0__lane22_strm1_cntl       ),      
               .std__pe0__lane22_strm1_data          ( std__pe0__lane22_strm1_data       ),      
               .std__pe0__lane22_strm1_data_valid    ( std__pe0__lane22_strm1_data_valid ),      
               .std__pe0__lane22_strm1_data_mask     ( std__pe0__lane22_strm1_data_mask  ),      

               // PE 0, Lane 23                 
               .pe0__std__lane23_strm0_ready         ( pe0__std__lane23_strm0_ready      ),      
               .std__pe0__lane23_strm0_cntl          ( std__pe0__lane23_strm0_cntl       ),      
               .std__pe0__lane23_strm0_data          ( std__pe0__lane23_strm0_data       ),      
               .std__pe0__lane23_strm0_data_valid    ( std__pe0__lane23_strm0_data_valid ),      
               .std__pe0__lane23_strm0_data_mask     ( std__pe0__lane23_strm0_data_mask  ),      

               .pe0__std__lane23_strm1_ready         ( pe0__std__lane23_strm1_ready      ),      
               .std__pe0__lane23_strm1_cntl          ( std__pe0__lane23_strm1_cntl       ),      
               .std__pe0__lane23_strm1_data          ( std__pe0__lane23_strm1_data       ),      
               .std__pe0__lane23_strm1_data_valid    ( std__pe0__lane23_strm1_data_valid ),      
               .std__pe0__lane23_strm1_data_mask     ( std__pe0__lane23_strm1_data_mask  ),      

               // PE 0, Lane 24                 
               .pe0__std__lane24_strm0_ready         ( pe0__std__lane24_strm0_ready      ),      
               .std__pe0__lane24_strm0_cntl          ( std__pe0__lane24_strm0_cntl       ),      
               .std__pe0__lane24_strm0_data          ( std__pe0__lane24_strm0_data       ),      
               .std__pe0__lane24_strm0_data_valid    ( std__pe0__lane24_strm0_data_valid ),      
               .std__pe0__lane24_strm0_data_mask     ( std__pe0__lane24_strm0_data_mask  ),      

               .pe0__std__lane24_strm1_ready         ( pe0__std__lane24_strm1_ready      ),      
               .std__pe0__lane24_strm1_cntl          ( std__pe0__lane24_strm1_cntl       ),      
               .std__pe0__lane24_strm1_data          ( std__pe0__lane24_strm1_data       ),      
               .std__pe0__lane24_strm1_data_valid    ( std__pe0__lane24_strm1_data_valid ),      
               .std__pe0__lane24_strm1_data_mask     ( std__pe0__lane24_strm1_data_mask  ),      

               // PE 0, Lane 25                 
               .pe0__std__lane25_strm0_ready         ( pe0__std__lane25_strm0_ready      ),      
               .std__pe0__lane25_strm0_cntl          ( std__pe0__lane25_strm0_cntl       ),      
               .std__pe0__lane25_strm0_data          ( std__pe0__lane25_strm0_data       ),      
               .std__pe0__lane25_strm0_data_valid    ( std__pe0__lane25_strm0_data_valid ),      
               .std__pe0__lane25_strm0_data_mask     ( std__pe0__lane25_strm0_data_mask  ),      

               .pe0__std__lane25_strm1_ready         ( pe0__std__lane25_strm1_ready      ),      
               .std__pe0__lane25_strm1_cntl          ( std__pe0__lane25_strm1_cntl       ),      
               .std__pe0__lane25_strm1_data          ( std__pe0__lane25_strm1_data       ),      
               .std__pe0__lane25_strm1_data_valid    ( std__pe0__lane25_strm1_data_valid ),      
               .std__pe0__lane25_strm1_data_mask     ( std__pe0__lane25_strm1_data_mask  ),      

               // PE 0, Lane 26                 
               .pe0__std__lane26_strm0_ready         ( pe0__std__lane26_strm0_ready      ),      
               .std__pe0__lane26_strm0_cntl          ( std__pe0__lane26_strm0_cntl       ),      
               .std__pe0__lane26_strm0_data          ( std__pe0__lane26_strm0_data       ),      
               .std__pe0__lane26_strm0_data_valid    ( std__pe0__lane26_strm0_data_valid ),      
               .std__pe0__lane26_strm0_data_mask     ( std__pe0__lane26_strm0_data_mask  ),      

               .pe0__std__lane26_strm1_ready         ( pe0__std__lane26_strm1_ready      ),      
               .std__pe0__lane26_strm1_cntl          ( std__pe0__lane26_strm1_cntl       ),      
               .std__pe0__lane26_strm1_data          ( std__pe0__lane26_strm1_data       ),      
               .std__pe0__lane26_strm1_data_valid    ( std__pe0__lane26_strm1_data_valid ),      
               .std__pe0__lane26_strm1_data_mask     ( std__pe0__lane26_strm1_data_mask  ),      

               // PE 0, Lane 27                 
               .pe0__std__lane27_strm0_ready         ( pe0__std__lane27_strm0_ready      ),      
               .std__pe0__lane27_strm0_cntl          ( std__pe0__lane27_strm0_cntl       ),      
               .std__pe0__lane27_strm0_data          ( std__pe0__lane27_strm0_data       ),      
               .std__pe0__lane27_strm0_data_valid    ( std__pe0__lane27_strm0_data_valid ),      
               .std__pe0__lane27_strm0_data_mask     ( std__pe0__lane27_strm0_data_mask  ),      

               .pe0__std__lane27_strm1_ready         ( pe0__std__lane27_strm1_ready      ),      
               .std__pe0__lane27_strm1_cntl          ( std__pe0__lane27_strm1_cntl       ),      
               .std__pe0__lane27_strm1_data          ( std__pe0__lane27_strm1_data       ),      
               .std__pe0__lane27_strm1_data_valid    ( std__pe0__lane27_strm1_data_valid ),      
               .std__pe0__lane27_strm1_data_mask     ( std__pe0__lane27_strm1_data_mask  ),      

               // PE 0, Lane 28                 
               .pe0__std__lane28_strm0_ready         ( pe0__std__lane28_strm0_ready      ),      
               .std__pe0__lane28_strm0_cntl          ( std__pe0__lane28_strm0_cntl       ),      
               .std__pe0__lane28_strm0_data          ( std__pe0__lane28_strm0_data       ),      
               .std__pe0__lane28_strm0_data_valid    ( std__pe0__lane28_strm0_data_valid ),      
               .std__pe0__lane28_strm0_data_mask     ( std__pe0__lane28_strm0_data_mask  ),      

               .pe0__std__lane28_strm1_ready         ( pe0__std__lane28_strm1_ready      ),      
               .std__pe0__lane28_strm1_cntl          ( std__pe0__lane28_strm1_cntl       ),      
               .std__pe0__lane28_strm1_data          ( std__pe0__lane28_strm1_data       ),      
               .std__pe0__lane28_strm1_data_valid    ( std__pe0__lane28_strm1_data_valid ),      
               .std__pe0__lane28_strm1_data_mask     ( std__pe0__lane28_strm1_data_mask  ),      

               // PE 0, Lane 29                 
               .pe0__std__lane29_strm0_ready         ( pe0__std__lane29_strm0_ready      ),      
               .std__pe0__lane29_strm0_cntl          ( std__pe0__lane29_strm0_cntl       ),      
               .std__pe0__lane29_strm0_data          ( std__pe0__lane29_strm0_data       ),      
               .std__pe0__lane29_strm0_data_valid    ( std__pe0__lane29_strm0_data_valid ),      
               .std__pe0__lane29_strm0_data_mask     ( std__pe0__lane29_strm0_data_mask  ),      

               .pe0__std__lane29_strm1_ready         ( pe0__std__lane29_strm1_ready      ),      
               .std__pe0__lane29_strm1_cntl          ( std__pe0__lane29_strm1_cntl       ),      
               .std__pe0__lane29_strm1_data          ( std__pe0__lane29_strm1_data       ),      
               .std__pe0__lane29_strm1_data_valid    ( std__pe0__lane29_strm1_data_valid ),      
               .std__pe0__lane29_strm1_data_mask     ( std__pe0__lane29_strm1_data_mask  ),      

               // PE 0, Lane 30                 
               .pe0__std__lane30_strm0_ready         ( pe0__std__lane30_strm0_ready      ),      
               .std__pe0__lane30_strm0_cntl          ( std__pe0__lane30_strm0_cntl       ),      
               .std__pe0__lane30_strm0_data          ( std__pe0__lane30_strm0_data       ),      
               .std__pe0__lane30_strm0_data_valid    ( std__pe0__lane30_strm0_data_valid ),      
               .std__pe0__lane30_strm0_data_mask     ( std__pe0__lane30_strm0_data_mask  ),      

               .pe0__std__lane30_strm1_ready         ( pe0__std__lane30_strm1_ready      ),      
               .std__pe0__lane30_strm1_cntl          ( std__pe0__lane30_strm1_cntl       ),      
               .std__pe0__lane30_strm1_data          ( std__pe0__lane30_strm1_data       ),      
               .std__pe0__lane30_strm1_data_valid    ( std__pe0__lane30_strm1_data_valid ),      
               .std__pe0__lane30_strm1_data_mask     ( std__pe0__lane30_strm1_data_mask  ),      

               // PE 0, Lane 31                 
               .pe0__std__lane31_strm0_ready         ( pe0__std__lane31_strm0_ready      ),      
               .std__pe0__lane31_strm0_cntl          ( std__pe0__lane31_strm0_cntl       ),      
               .std__pe0__lane31_strm0_data          ( std__pe0__lane31_strm0_data       ),      
               .std__pe0__lane31_strm0_data_valid    ( std__pe0__lane31_strm0_data_valid ),      
               .std__pe0__lane31_strm0_data_mask     ( std__pe0__lane31_strm0_data_mask  ),      

               .pe0__std__lane31_strm1_ready         ( pe0__std__lane31_strm1_ready      ),      
               .std__pe0__lane31_strm1_cntl          ( std__pe0__lane31_strm1_cntl       ),      
               .std__pe0__lane31_strm1_data          ( std__pe0__lane31_strm1_data       ),      
               .std__pe0__lane31_strm1_data_valid    ( std__pe0__lane31_strm1_data_valid ),      
               .std__pe0__lane31_strm1_data_mask     ( std__pe0__lane31_strm1_data_mask  ),      

               // PE 1, Lane 0                 
               .pe1__std__lane0_strm0_ready         ( pe1__std__lane0_strm0_ready      ),      
               .std__pe1__lane0_strm0_cntl          ( std__pe1__lane0_strm0_cntl       ),      
               .std__pe1__lane0_strm0_data          ( std__pe1__lane0_strm0_data       ),      
               .std__pe1__lane0_strm0_data_valid    ( std__pe1__lane0_strm0_data_valid ),      
               .std__pe1__lane0_strm0_data_mask     ( std__pe1__lane0_strm0_data_mask  ),      

               .pe1__std__lane0_strm1_ready         ( pe1__std__lane0_strm1_ready      ),      
               .std__pe1__lane0_strm1_cntl          ( std__pe1__lane0_strm1_cntl       ),      
               .std__pe1__lane0_strm1_data          ( std__pe1__lane0_strm1_data       ),      
               .std__pe1__lane0_strm1_data_valid    ( std__pe1__lane0_strm1_data_valid ),      
               .std__pe1__lane0_strm1_data_mask     ( std__pe1__lane0_strm1_data_mask  ),      

               // PE 1, Lane 1                 
               .pe1__std__lane1_strm0_ready         ( pe1__std__lane1_strm0_ready      ),      
               .std__pe1__lane1_strm0_cntl          ( std__pe1__lane1_strm0_cntl       ),      
               .std__pe1__lane1_strm0_data          ( std__pe1__lane1_strm0_data       ),      
               .std__pe1__lane1_strm0_data_valid    ( std__pe1__lane1_strm0_data_valid ),      
               .std__pe1__lane1_strm0_data_mask     ( std__pe1__lane1_strm0_data_mask  ),      

               .pe1__std__lane1_strm1_ready         ( pe1__std__lane1_strm1_ready      ),      
               .std__pe1__lane1_strm1_cntl          ( std__pe1__lane1_strm1_cntl       ),      
               .std__pe1__lane1_strm1_data          ( std__pe1__lane1_strm1_data       ),      
               .std__pe1__lane1_strm1_data_valid    ( std__pe1__lane1_strm1_data_valid ),      
               .std__pe1__lane1_strm1_data_mask     ( std__pe1__lane1_strm1_data_mask  ),      

               // PE 1, Lane 2                 
               .pe1__std__lane2_strm0_ready         ( pe1__std__lane2_strm0_ready      ),      
               .std__pe1__lane2_strm0_cntl          ( std__pe1__lane2_strm0_cntl       ),      
               .std__pe1__lane2_strm0_data          ( std__pe1__lane2_strm0_data       ),      
               .std__pe1__lane2_strm0_data_valid    ( std__pe1__lane2_strm0_data_valid ),      
               .std__pe1__lane2_strm0_data_mask     ( std__pe1__lane2_strm0_data_mask  ),      

               .pe1__std__lane2_strm1_ready         ( pe1__std__lane2_strm1_ready      ),      
               .std__pe1__lane2_strm1_cntl          ( std__pe1__lane2_strm1_cntl       ),      
               .std__pe1__lane2_strm1_data          ( std__pe1__lane2_strm1_data       ),      
               .std__pe1__lane2_strm1_data_valid    ( std__pe1__lane2_strm1_data_valid ),      
               .std__pe1__lane2_strm1_data_mask     ( std__pe1__lane2_strm1_data_mask  ),      

               // PE 1, Lane 3                 
               .pe1__std__lane3_strm0_ready         ( pe1__std__lane3_strm0_ready      ),      
               .std__pe1__lane3_strm0_cntl          ( std__pe1__lane3_strm0_cntl       ),      
               .std__pe1__lane3_strm0_data          ( std__pe1__lane3_strm0_data       ),      
               .std__pe1__lane3_strm0_data_valid    ( std__pe1__lane3_strm0_data_valid ),      
               .std__pe1__lane3_strm0_data_mask     ( std__pe1__lane3_strm0_data_mask  ),      

               .pe1__std__lane3_strm1_ready         ( pe1__std__lane3_strm1_ready      ),      
               .std__pe1__lane3_strm1_cntl          ( std__pe1__lane3_strm1_cntl       ),      
               .std__pe1__lane3_strm1_data          ( std__pe1__lane3_strm1_data       ),      
               .std__pe1__lane3_strm1_data_valid    ( std__pe1__lane3_strm1_data_valid ),      
               .std__pe1__lane3_strm1_data_mask     ( std__pe1__lane3_strm1_data_mask  ),      

               // PE 1, Lane 4                 
               .pe1__std__lane4_strm0_ready         ( pe1__std__lane4_strm0_ready      ),      
               .std__pe1__lane4_strm0_cntl          ( std__pe1__lane4_strm0_cntl       ),      
               .std__pe1__lane4_strm0_data          ( std__pe1__lane4_strm0_data       ),      
               .std__pe1__lane4_strm0_data_valid    ( std__pe1__lane4_strm0_data_valid ),      
               .std__pe1__lane4_strm0_data_mask     ( std__pe1__lane4_strm0_data_mask  ),      

               .pe1__std__lane4_strm1_ready         ( pe1__std__lane4_strm1_ready      ),      
               .std__pe1__lane4_strm1_cntl          ( std__pe1__lane4_strm1_cntl       ),      
               .std__pe1__lane4_strm1_data          ( std__pe1__lane4_strm1_data       ),      
               .std__pe1__lane4_strm1_data_valid    ( std__pe1__lane4_strm1_data_valid ),      
               .std__pe1__lane4_strm1_data_mask     ( std__pe1__lane4_strm1_data_mask  ),      

               // PE 1, Lane 5                 
               .pe1__std__lane5_strm0_ready         ( pe1__std__lane5_strm0_ready      ),      
               .std__pe1__lane5_strm0_cntl          ( std__pe1__lane5_strm0_cntl       ),      
               .std__pe1__lane5_strm0_data          ( std__pe1__lane5_strm0_data       ),      
               .std__pe1__lane5_strm0_data_valid    ( std__pe1__lane5_strm0_data_valid ),      
               .std__pe1__lane5_strm0_data_mask     ( std__pe1__lane5_strm0_data_mask  ),      

               .pe1__std__lane5_strm1_ready         ( pe1__std__lane5_strm1_ready      ),      
               .std__pe1__lane5_strm1_cntl          ( std__pe1__lane5_strm1_cntl       ),      
               .std__pe1__lane5_strm1_data          ( std__pe1__lane5_strm1_data       ),      
               .std__pe1__lane5_strm1_data_valid    ( std__pe1__lane5_strm1_data_valid ),      
               .std__pe1__lane5_strm1_data_mask     ( std__pe1__lane5_strm1_data_mask  ),      

               // PE 1, Lane 6                 
               .pe1__std__lane6_strm0_ready         ( pe1__std__lane6_strm0_ready      ),      
               .std__pe1__lane6_strm0_cntl          ( std__pe1__lane6_strm0_cntl       ),      
               .std__pe1__lane6_strm0_data          ( std__pe1__lane6_strm0_data       ),      
               .std__pe1__lane6_strm0_data_valid    ( std__pe1__lane6_strm0_data_valid ),      
               .std__pe1__lane6_strm0_data_mask     ( std__pe1__lane6_strm0_data_mask  ),      

               .pe1__std__lane6_strm1_ready         ( pe1__std__lane6_strm1_ready      ),      
               .std__pe1__lane6_strm1_cntl          ( std__pe1__lane6_strm1_cntl       ),      
               .std__pe1__lane6_strm1_data          ( std__pe1__lane6_strm1_data       ),      
               .std__pe1__lane6_strm1_data_valid    ( std__pe1__lane6_strm1_data_valid ),      
               .std__pe1__lane6_strm1_data_mask     ( std__pe1__lane6_strm1_data_mask  ),      

               // PE 1, Lane 7                 
               .pe1__std__lane7_strm0_ready         ( pe1__std__lane7_strm0_ready      ),      
               .std__pe1__lane7_strm0_cntl          ( std__pe1__lane7_strm0_cntl       ),      
               .std__pe1__lane7_strm0_data          ( std__pe1__lane7_strm0_data       ),      
               .std__pe1__lane7_strm0_data_valid    ( std__pe1__lane7_strm0_data_valid ),      
               .std__pe1__lane7_strm0_data_mask     ( std__pe1__lane7_strm0_data_mask  ),      

               .pe1__std__lane7_strm1_ready         ( pe1__std__lane7_strm1_ready      ),      
               .std__pe1__lane7_strm1_cntl          ( std__pe1__lane7_strm1_cntl       ),      
               .std__pe1__lane7_strm1_data          ( std__pe1__lane7_strm1_data       ),      
               .std__pe1__lane7_strm1_data_valid    ( std__pe1__lane7_strm1_data_valid ),      
               .std__pe1__lane7_strm1_data_mask     ( std__pe1__lane7_strm1_data_mask  ),      

               // PE 1, Lane 8                 
               .pe1__std__lane8_strm0_ready         ( pe1__std__lane8_strm0_ready      ),      
               .std__pe1__lane8_strm0_cntl          ( std__pe1__lane8_strm0_cntl       ),      
               .std__pe1__lane8_strm0_data          ( std__pe1__lane8_strm0_data       ),      
               .std__pe1__lane8_strm0_data_valid    ( std__pe1__lane8_strm0_data_valid ),      
               .std__pe1__lane8_strm0_data_mask     ( std__pe1__lane8_strm0_data_mask  ),      

               .pe1__std__lane8_strm1_ready         ( pe1__std__lane8_strm1_ready      ),      
               .std__pe1__lane8_strm1_cntl          ( std__pe1__lane8_strm1_cntl       ),      
               .std__pe1__lane8_strm1_data          ( std__pe1__lane8_strm1_data       ),      
               .std__pe1__lane8_strm1_data_valid    ( std__pe1__lane8_strm1_data_valid ),      
               .std__pe1__lane8_strm1_data_mask     ( std__pe1__lane8_strm1_data_mask  ),      

               // PE 1, Lane 9                 
               .pe1__std__lane9_strm0_ready         ( pe1__std__lane9_strm0_ready      ),      
               .std__pe1__lane9_strm0_cntl          ( std__pe1__lane9_strm0_cntl       ),      
               .std__pe1__lane9_strm0_data          ( std__pe1__lane9_strm0_data       ),      
               .std__pe1__lane9_strm0_data_valid    ( std__pe1__lane9_strm0_data_valid ),      
               .std__pe1__lane9_strm0_data_mask     ( std__pe1__lane9_strm0_data_mask  ),      

               .pe1__std__lane9_strm1_ready         ( pe1__std__lane9_strm1_ready      ),      
               .std__pe1__lane9_strm1_cntl          ( std__pe1__lane9_strm1_cntl       ),      
               .std__pe1__lane9_strm1_data          ( std__pe1__lane9_strm1_data       ),      
               .std__pe1__lane9_strm1_data_valid    ( std__pe1__lane9_strm1_data_valid ),      
               .std__pe1__lane9_strm1_data_mask     ( std__pe1__lane9_strm1_data_mask  ),      

               // PE 1, Lane 10                 
               .pe1__std__lane10_strm0_ready         ( pe1__std__lane10_strm0_ready      ),      
               .std__pe1__lane10_strm0_cntl          ( std__pe1__lane10_strm0_cntl       ),      
               .std__pe1__lane10_strm0_data          ( std__pe1__lane10_strm0_data       ),      
               .std__pe1__lane10_strm0_data_valid    ( std__pe1__lane10_strm0_data_valid ),      
               .std__pe1__lane10_strm0_data_mask     ( std__pe1__lane10_strm0_data_mask  ),      

               .pe1__std__lane10_strm1_ready         ( pe1__std__lane10_strm1_ready      ),      
               .std__pe1__lane10_strm1_cntl          ( std__pe1__lane10_strm1_cntl       ),      
               .std__pe1__lane10_strm1_data          ( std__pe1__lane10_strm1_data       ),      
               .std__pe1__lane10_strm1_data_valid    ( std__pe1__lane10_strm1_data_valid ),      
               .std__pe1__lane10_strm1_data_mask     ( std__pe1__lane10_strm1_data_mask  ),      

               // PE 1, Lane 11                 
               .pe1__std__lane11_strm0_ready         ( pe1__std__lane11_strm0_ready      ),      
               .std__pe1__lane11_strm0_cntl          ( std__pe1__lane11_strm0_cntl       ),      
               .std__pe1__lane11_strm0_data          ( std__pe1__lane11_strm0_data       ),      
               .std__pe1__lane11_strm0_data_valid    ( std__pe1__lane11_strm0_data_valid ),      
               .std__pe1__lane11_strm0_data_mask     ( std__pe1__lane11_strm0_data_mask  ),      

               .pe1__std__lane11_strm1_ready         ( pe1__std__lane11_strm1_ready      ),      
               .std__pe1__lane11_strm1_cntl          ( std__pe1__lane11_strm1_cntl       ),      
               .std__pe1__lane11_strm1_data          ( std__pe1__lane11_strm1_data       ),      
               .std__pe1__lane11_strm1_data_valid    ( std__pe1__lane11_strm1_data_valid ),      
               .std__pe1__lane11_strm1_data_mask     ( std__pe1__lane11_strm1_data_mask  ),      

               // PE 1, Lane 12                 
               .pe1__std__lane12_strm0_ready         ( pe1__std__lane12_strm0_ready      ),      
               .std__pe1__lane12_strm0_cntl          ( std__pe1__lane12_strm0_cntl       ),      
               .std__pe1__lane12_strm0_data          ( std__pe1__lane12_strm0_data       ),      
               .std__pe1__lane12_strm0_data_valid    ( std__pe1__lane12_strm0_data_valid ),      
               .std__pe1__lane12_strm0_data_mask     ( std__pe1__lane12_strm0_data_mask  ),      

               .pe1__std__lane12_strm1_ready         ( pe1__std__lane12_strm1_ready      ),      
               .std__pe1__lane12_strm1_cntl          ( std__pe1__lane12_strm1_cntl       ),      
               .std__pe1__lane12_strm1_data          ( std__pe1__lane12_strm1_data       ),      
               .std__pe1__lane12_strm1_data_valid    ( std__pe1__lane12_strm1_data_valid ),      
               .std__pe1__lane12_strm1_data_mask     ( std__pe1__lane12_strm1_data_mask  ),      

               // PE 1, Lane 13                 
               .pe1__std__lane13_strm0_ready         ( pe1__std__lane13_strm0_ready      ),      
               .std__pe1__lane13_strm0_cntl          ( std__pe1__lane13_strm0_cntl       ),      
               .std__pe1__lane13_strm0_data          ( std__pe1__lane13_strm0_data       ),      
               .std__pe1__lane13_strm0_data_valid    ( std__pe1__lane13_strm0_data_valid ),      
               .std__pe1__lane13_strm0_data_mask     ( std__pe1__lane13_strm0_data_mask  ),      

               .pe1__std__lane13_strm1_ready         ( pe1__std__lane13_strm1_ready      ),      
               .std__pe1__lane13_strm1_cntl          ( std__pe1__lane13_strm1_cntl       ),      
               .std__pe1__lane13_strm1_data          ( std__pe1__lane13_strm1_data       ),      
               .std__pe1__lane13_strm1_data_valid    ( std__pe1__lane13_strm1_data_valid ),      
               .std__pe1__lane13_strm1_data_mask     ( std__pe1__lane13_strm1_data_mask  ),      

               // PE 1, Lane 14                 
               .pe1__std__lane14_strm0_ready         ( pe1__std__lane14_strm0_ready      ),      
               .std__pe1__lane14_strm0_cntl          ( std__pe1__lane14_strm0_cntl       ),      
               .std__pe1__lane14_strm0_data          ( std__pe1__lane14_strm0_data       ),      
               .std__pe1__lane14_strm0_data_valid    ( std__pe1__lane14_strm0_data_valid ),      
               .std__pe1__lane14_strm0_data_mask     ( std__pe1__lane14_strm0_data_mask  ),      

               .pe1__std__lane14_strm1_ready         ( pe1__std__lane14_strm1_ready      ),      
               .std__pe1__lane14_strm1_cntl          ( std__pe1__lane14_strm1_cntl       ),      
               .std__pe1__lane14_strm1_data          ( std__pe1__lane14_strm1_data       ),      
               .std__pe1__lane14_strm1_data_valid    ( std__pe1__lane14_strm1_data_valid ),      
               .std__pe1__lane14_strm1_data_mask     ( std__pe1__lane14_strm1_data_mask  ),      

               // PE 1, Lane 15                 
               .pe1__std__lane15_strm0_ready         ( pe1__std__lane15_strm0_ready      ),      
               .std__pe1__lane15_strm0_cntl          ( std__pe1__lane15_strm0_cntl       ),      
               .std__pe1__lane15_strm0_data          ( std__pe1__lane15_strm0_data       ),      
               .std__pe1__lane15_strm0_data_valid    ( std__pe1__lane15_strm0_data_valid ),      
               .std__pe1__lane15_strm0_data_mask     ( std__pe1__lane15_strm0_data_mask  ),      

               .pe1__std__lane15_strm1_ready         ( pe1__std__lane15_strm1_ready      ),      
               .std__pe1__lane15_strm1_cntl          ( std__pe1__lane15_strm1_cntl       ),      
               .std__pe1__lane15_strm1_data          ( std__pe1__lane15_strm1_data       ),      
               .std__pe1__lane15_strm1_data_valid    ( std__pe1__lane15_strm1_data_valid ),      
               .std__pe1__lane15_strm1_data_mask     ( std__pe1__lane15_strm1_data_mask  ),      

               // PE 1, Lane 16                 
               .pe1__std__lane16_strm0_ready         ( pe1__std__lane16_strm0_ready      ),      
               .std__pe1__lane16_strm0_cntl          ( std__pe1__lane16_strm0_cntl       ),      
               .std__pe1__lane16_strm0_data          ( std__pe1__lane16_strm0_data       ),      
               .std__pe1__lane16_strm0_data_valid    ( std__pe1__lane16_strm0_data_valid ),      
               .std__pe1__lane16_strm0_data_mask     ( std__pe1__lane16_strm0_data_mask  ),      

               .pe1__std__lane16_strm1_ready         ( pe1__std__lane16_strm1_ready      ),      
               .std__pe1__lane16_strm1_cntl          ( std__pe1__lane16_strm1_cntl       ),      
               .std__pe1__lane16_strm1_data          ( std__pe1__lane16_strm1_data       ),      
               .std__pe1__lane16_strm1_data_valid    ( std__pe1__lane16_strm1_data_valid ),      
               .std__pe1__lane16_strm1_data_mask     ( std__pe1__lane16_strm1_data_mask  ),      

               // PE 1, Lane 17                 
               .pe1__std__lane17_strm0_ready         ( pe1__std__lane17_strm0_ready      ),      
               .std__pe1__lane17_strm0_cntl          ( std__pe1__lane17_strm0_cntl       ),      
               .std__pe1__lane17_strm0_data          ( std__pe1__lane17_strm0_data       ),      
               .std__pe1__lane17_strm0_data_valid    ( std__pe1__lane17_strm0_data_valid ),      
               .std__pe1__lane17_strm0_data_mask     ( std__pe1__lane17_strm0_data_mask  ),      

               .pe1__std__lane17_strm1_ready         ( pe1__std__lane17_strm1_ready      ),      
               .std__pe1__lane17_strm1_cntl          ( std__pe1__lane17_strm1_cntl       ),      
               .std__pe1__lane17_strm1_data          ( std__pe1__lane17_strm1_data       ),      
               .std__pe1__lane17_strm1_data_valid    ( std__pe1__lane17_strm1_data_valid ),      
               .std__pe1__lane17_strm1_data_mask     ( std__pe1__lane17_strm1_data_mask  ),      

               // PE 1, Lane 18                 
               .pe1__std__lane18_strm0_ready         ( pe1__std__lane18_strm0_ready      ),      
               .std__pe1__lane18_strm0_cntl          ( std__pe1__lane18_strm0_cntl       ),      
               .std__pe1__lane18_strm0_data          ( std__pe1__lane18_strm0_data       ),      
               .std__pe1__lane18_strm0_data_valid    ( std__pe1__lane18_strm0_data_valid ),      
               .std__pe1__lane18_strm0_data_mask     ( std__pe1__lane18_strm0_data_mask  ),      

               .pe1__std__lane18_strm1_ready         ( pe1__std__lane18_strm1_ready      ),      
               .std__pe1__lane18_strm1_cntl          ( std__pe1__lane18_strm1_cntl       ),      
               .std__pe1__lane18_strm1_data          ( std__pe1__lane18_strm1_data       ),      
               .std__pe1__lane18_strm1_data_valid    ( std__pe1__lane18_strm1_data_valid ),      
               .std__pe1__lane18_strm1_data_mask     ( std__pe1__lane18_strm1_data_mask  ),      

               // PE 1, Lane 19                 
               .pe1__std__lane19_strm0_ready         ( pe1__std__lane19_strm0_ready      ),      
               .std__pe1__lane19_strm0_cntl          ( std__pe1__lane19_strm0_cntl       ),      
               .std__pe1__lane19_strm0_data          ( std__pe1__lane19_strm0_data       ),      
               .std__pe1__lane19_strm0_data_valid    ( std__pe1__lane19_strm0_data_valid ),      
               .std__pe1__lane19_strm0_data_mask     ( std__pe1__lane19_strm0_data_mask  ),      

               .pe1__std__lane19_strm1_ready         ( pe1__std__lane19_strm1_ready      ),      
               .std__pe1__lane19_strm1_cntl          ( std__pe1__lane19_strm1_cntl       ),      
               .std__pe1__lane19_strm1_data          ( std__pe1__lane19_strm1_data       ),      
               .std__pe1__lane19_strm1_data_valid    ( std__pe1__lane19_strm1_data_valid ),      
               .std__pe1__lane19_strm1_data_mask     ( std__pe1__lane19_strm1_data_mask  ),      

               // PE 1, Lane 20                 
               .pe1__std__lane20_strm0_ready         ( pe1__std__lane20_strm0_ready      ),      
               .std__pe1__lane20_strm0_cntl          ( std__pe1__lane20_strm0_cntl       ),      
               .std__pe1__lane20_strm0_data          ( std__pe1__lane20_strm0_data       ),      
               .std__pe1__lane20_strm0_data_valid    ( std__pe1__lane20_strm0_data_valid ),      
               .std__pe1__lane20_strm0_data_mask     ( std__pe1__lane20_strm0_data_mask  ),      

               .pe1__std__lane20_strm1_ready         ( pe1__std__lane20_strm1_ready      ),      
               .std__pe1__lane20_strm1_cntl          ( std__pe1__lane20_strm1_cntl       ),      
               .std__pe1__lane20_strm1_data          ( std__pe1__lane20_strm1_data       ),      
               .std__pe1__lane20_strm1_data_valid    ( std__pe1__lane20_strm1_data_valid ),      
               .std__pe1__lane20_strm1_data_mask     ( std__pe1__lane20_strm1_data_mask  ),      

               // PE 1, Lane 21                 
               .pe1__std__lane21_strm0_ready         ( pe1__std__lane21_strm0_ready      ),      
               .std__pe1__lane21_strm0_cntl          ( std__pe1__lane21_strm0_cntl       ),      
               .std__pe1__lane21_strm0_data          ( std__pe1__lane21_strm0_data       ),      
               .std__pe1__lane21_strm0_data_valid    ( std__pe1__lane21_strm0_data_valid ),      
               .std__pe1__lane21_strm0_data_mask     ( std__pe1__lane21_strm0_data_mask  ),      

               .pe1__std__lane21_strm1_ready         ( pe1__std__lane21_strm1_ready      ),      
               .std__pe1__lane21_strm1_cntl          ( std__pe1__lane21_strm1_cntl       ),      
               .std__pe1__lane21_strm1_data          ( std__pe1__lane21_strm1_data       ),      
               .std__pe1__lane21_strm1_data_valid    ( std__pe1__lane21_strm1_data_valid ),      
               .std__pe1__lane21_strm1_data_mask     ( std__pe1__lane21_strm1_data_mask  ),      

               // PE 1, Lane 22                 
               .pe1__std__lane22_strm0_ready         ( pe1__std__lane22_strm0_ready      ),      
               .std__pe1__lane22_strm0_cntl          ( std__pe1__lane22_strm0_cntl       ),      
               .std__pe1__lane22_strm0_data          ( std__pe1__lane22_strm0_data       ),      
               .std__pe1__lane22_strm0_data_valid    ( std__pe1__lane22_strm0_data_valid ),      
               .std__pe1__lane22_strm0_data_mask     ( std__pe1__lane22_strm0_data_mask  ),      

               .pe1__std__lane22_strm1_ready         ( pe1__std__lane22_strm1_ready      ),      
               .std__pe1__lane22_strm1_cntl          ( std__pe1__lane22_strm1_cntl       ),      
               .std__pe1__lane22_strm1_data          ( std__pe1__lane22_strm1_data       ),      
               .std__pe1__lane22_strm1_data_valid    ( std__pe1__lane22_strm1_data_valid ),      
               .std__pe1__lane22_strm1_data_mask     ( std__pe1__lane22_strm1_data_mask  ),      

               // PE 1, Lane 23                 
               .pe1__std__lane23_strm0_ready         ( pe1__std__lane23_strm0_ready      ),      
               .std__pe1__lane23_strm0_cntl          ( std__pe1__lane23_strm0_cntl       ),      
               .std__pe1__lane23_strm0_data          ( std__pe1__lane23_strm0_data       ),      
               .std__pe1__lane23_strm0_data_valid    ( std__pe1__lane23_strm0_data_valid ),      
               .std__pe1__lane23_strm0_data_mask     ( std__pe1__lane23_strm0_data_mask  ),      

               .pe1__std__lane23_strm1_ready         ( pe1__std__lane23_strm1_ready      ),      
               .std__pe1__lane23_strm1_cntl          ( std__pe1__lane23_strm1_cntl       ),      
               .std__pe1__lane23_strm1_data          ( std__pe1__lane23_strm1_data       ),      
               .std__pe1__lane23_strm1_data_valid    ( std__pe1__lane23_strm1_data_valid ),      
               .std__pe1__lane23_strm1_data_mask     ( std__pe1__lane23_strm1_data_mask  ),      

               // PE 1, Lane 24                 
               .pe1__std__lane24_strm0_ready         ( pe1__std__lane24_strm0_ready      ),      
               .std__pe1__lane24_strm0_cntl          ( std__pe1__lane24_strm0_cntl       ),      
               .std__pe1__lane24_strm0_data          ( std__pe1__lane24_strm0_data       ),      
               .std__pe1__lane24_strm0_data_valid    ( std__pe1__lane24_strm0_data_valid ),      
               .std__pe1__lane24_strm0_data_mask     ( std__pe1__lane24_strm0_data_mask  ),      

               .pe1__std__lane24_strm1_ready         ( pe1__std__lane24_strm1_ready      ),      
               .std__pe1__lane24_strm1_cntl          ( std__pe1__lane24_strm1_cntl       ),      
               .std__pe1__lane24_strm1_data          ( std__pe1__lane24_strm1_data       ),      
               .std__pe1__lane24_strm1_data_valid    ( std__pe1__lane24_strm1_data_valid ),      
               .std__pe1__lane24_strm1_data_mask     ( std__pe1__lane24_strm1_data_mask  ),      

               // PE 1, Lane 25                 
               .pe1__std__lane25_strm0_ready         ( pe1__std__lane25_strm0_ready      ),      
               .std__pe1__lane25_strm0_cntl          ( std__pe1__lane25_strm0_cntl       ),      
               .std__pe1__lane25_strm0_data          ( std__pe1__lane25_strm0_data       ),      
               .std__pe1__lane25_strm0_data_valid    ( std__pe1__lane25_strm0_data_valid ),      
               .std__pe1__lane25_strm0_data_mask     ( std__pe1__lane25_strm0_data_mask  ),      

               .pe1__std__lane25_strm1_ready         ( pe1__std__lane25_strm1_ready      ),      
               .std__pe1__lane25_strm1_cntl          ( std__pe1__lane25_strm1_cntl       ),      
               .std__pe1__lane25_strm1_data          ( std__pe1__lane25_strm1_data       ),      
               .std__pe1__lane25_strm1_data_valid    ( std__pe1__lane25_strm1_data_valid ),      
               .std__pe1__lane25_strm1_data_mask     ( std__pe1__lane25_strm1_data_mask  ),      

               // PE 1, Lane 26                 
               .pe1__std__lane26_strm0_ready         ( pe1__std__lane26_strm0_ready      ),      
               .std__pe1__lane26_strm0_cntl          ( std__pe1__lane26_strm0_cntl       ),      
               .std__pe1__lane26_strm0_data          ( std__pe1__lane26_strm0_data       ),      
               .std__pe1__lane26_strm0_data_valid    ( std__pe1__lane26_strm0_data_valid ),      
               .std__pe1__lane26_strm0_data_mask     ( std__pe1__lane26_strm0_data_mask  ),      

               .pe1__std__lane26_strm1_ready         ( pe1__std__lane26_strm1_ready      ),      
               .std__pe1__lane26_strm1_cntl          ( std__pe1__lane26_strm1_cntl       ),      
               .std__pe1__lane26_strm1_data          ( std__pe1__lane26_strm1_data       ),      
               .std__pe1__lane26_strm1_data_valid    ( std__pe1__lane26_strm1_data_valid ),      
               .std__pe1__lane26_strm1_data_mask     ( std__pe1__lane26_strm1_data_mask  ),      

               // PE 1, Lane 27                 
               .pe1__std__lane27_strm0_ready         ( pe1__std__lane27_strm0_ready      ),      
               .std__pe1__lane27_strm0_cntl          ( std__pe1__lane27_strm0_cntl       ),      
               .std__pe1__lane27_strm0_data          ( std__pe1__lane27_strm0_data       ),      
               .std__pe1__lane27_strm0_data_valid    ( std__pe1__lane27_strm0_data_valid ),      
               .std__pe1__lane27_strm0_data_mask     ( std__pe1__lane27_strm0_data_mask  ),      

               .pe1__std__lane27_strm1_ready         ( pe1__std__lane27_strm1_ready      ),      
               .std__pe1__lane27_strm1_cntl          ( std__pe1__lane27_strm1_cntl       ),      
               .std__pe1__lane27_strm1_data          ( std__pe1__lane27_strm1_data       ),      
               .std__pe1__lane27_strm1_data_valid    ( std__pe1__lane27_strm1_data_valid ),      
               .std__pe1__lane27_strm1_data_mask     ( std__pe1__lane27_strm1_data_mask  ),      

               // PE 1, Lane 28                 
               .pe1__std__lane28_strm0_ready         ( pe1__std__lane28_strm0_ready      ),      
               .std__pe1__lane28_strm0_cntl          ( std__pe1__lane28_strm0_cntl       ),      
               .std__pe1__lane28_strm0_data          ( std__pe1__lane28_strm0_data       ),      
               .std__pe1__lane28_strm0_data_valid    ( std__pe1__lane28_strm0_data_valid ),      
               .std__pe1__lane28_strm0_data_mask     ( std__pe1__lane28_strm0_data_mask  ),      

               .pe1__std__lane28_strm1_ready         ( pe1__std__lane28_strm1_ready      ),      
               .std__pe1__lane28_strm1_cntl          ( std__pe1__lane28_strm1_cntl       ),      
               .std__pe1__lane28_strm1_data          ( std__pe1__lane28_strm1_data       ),      
               .std__pe1__lane28_strm1_data_valid    ( std__pe1__lane28_strm1_data_valid ),      
               .std__pe1__lane28_strm1_data_mask     ( std__pe1__lane28_strm1_data_mask  ),      

               // PE 1, Lane 29                 
               .pe1__std__lane29_strm0_ready         ( pe1__std__lane29_strm0_ready      ),      
               .std__pe1__lane29_strm0_cntl          ( std__pe1__lane29_strm0_cntl       ),      
               .std__pe1__lane29_strm0_data          ( std__pe1__lane29_strm0_data       ),      
               .std__pe1__lane29_strm0_data_valid    ( std__pe1__lane29_strm0_data_valid ),      
               .std__pe1__lane29_strm0_data_mask     ( std__pe1__lane29_strm0_data_mask  ),      

               .pe1__std__lane29_strm1_ready         ( pe1__std__lane29_strm1_ready      ),      
               .std__pe1__lane29_strm1_cntl          ( std__pe1__lane29_strm1_cntl       ),      
               .std__pe1__lane29_strm1_data          ( std__pe1__lane29_strm1_data       ),      
               .std__pe1__lane29_strm1_data_valid    ( std__pe1__lane29_strm1_data_valid ),      
               .std__pe1__lane29_strm1_data_mask     ( std__pe1__lane29_strm1_data_mask  ),      

               // PE 1, Lane 30                 
               .pe1__std__lane30_strm0_ready         ( pe1__std__lane30_strm0_ready      ),      
               .std__pe1__lane30_strm0_cntl          ( std__pe1__lane30_strm0_cntl       ),      
               .std__pe1__lane30_strm0_data          ( std__pe1__lane30_strm0_data       ),      
               .std__pe1__lane30_strm0_data_valid    ( std__pe1__lane30_strm0_data_valid ),      
               .std__pe1__lane30_strm0_data_mask     ( std__pe1__lane30_strm0_data_mask  ),      

               .pe1__std__lane30_strm1_ready         ( pe1__std__lane30_strm1_ready      ),      
               .std__pe1__lane30_strm1_cntl          ( std__pe1__lane30_strm1_cntl       ),      
               .std__pe1__lane30_strm1_data          ( std__pe1__lane30_strm1_data       ),      
               .std__pe1__lane30_strm1_data_valid    ( std__pe1__lane30_strm1_data_valid ),      
               .std__pe1__lane30_strm1_data_mask     ( std__pe1__lane30_strm1_data_mask  ),      

               // PE 1, Lane 31                 
               .pe1__std__lane31_strm0_ready         ( pe1__std__lane31_strm0_ready      ),      
               .std__pe1__lane31_strm0_cntl          ( std__pe1__lane31_strm0_cntl       ),      
               .std__pe1__lane31_strm0_data          ( std__pe1__lane31_strm0_data       ),      
               .std__pe1__lane31_strm0_data_valid    ( std__pe1__lane31_strm0_data_valid ),      
               .std__pe1__lane31_strm0_data_mask     ( std__pe1__lane31_strm0_data_mask  ),      

               .pe1__std__lane31_strm1_ready         ( pe1__std__lane31_strm1_ready      ),      
               .std__pe1__lane31_strm1_cntl          ( std__pe1__lane31_strm1_cntl       ),      
               .std__pe1__lane31_strm1_data          ( std__pe1__lane31_strm1_data       ),      
               .std__pe1__lane31_strm1_data_valid    ( std__pe1__lane31_strm1_data_valid ),      
               .std__pe1__lane31_strm1_data_mask     ( std__pe1__lane31_strm1_data_mask  ),      

               // PE 2, Lane 0                 
               .pe2__std__lane0_strm0_ready         ( pe2__std__lane0_strm0_ready      ),      
               .std__pe2__lane0_strm0_cntl          ( std__pe2__lane0_strm0_cntl       ),      
               .std__pe2__lane0_strm0_data          ( std__pe2__lane0_strm0_data       ),      
               .std__pe2__lane0_strm0_data_valid    ( std__pe2__lane0_strm0_data_valid ),      
               .std__pe2__lane0_strm0_data_mask     ( std__pe2__lane0_strm0_data_mask  ),      

               .pe2__std__lane0_strm1_ready         ( pe2__std__lane0_strm1_ready      ),      
               .std__pe2__lane0_strm1_cntl          ( std__pe2__lane0_strm1_cntl       ),      
               .std__pe2__lane0_strm1_data          ( std__pe2__lane0_strm1_data       ),      
               .std__pe2__lane0_strm1_data_valid    ( std__pe2__lane0_strm1_data_valid ),      
               .std__pe2__lane0_strm1_data_mask     ( std__pe2__lane0_strm1_data_mask  ),      

               // PE 2, Lane 1                 
               .pe2__std__lane1_strm0_ready         ( pe2__std__lane1_strm0_ready      ),      
               .std__pe2__lane1_strm0_cntl          ( std__pe2__lane1_strm0_cntl       ),      
               .std__pe2__lane1_strm0_data          ( std__pe2__lane1_strm0_data       ),      
               .std__pe2__lane1_strm0_data_valid    ( std__pe2__lane1_strm0_data_valid ),      
               .std__pe2__lane1_strm0_data_mask     ( std__pe2__lane1_strm0_data_mask  ),      

               .pe2__std__lane1_strm1_ready         ( pe2__std__lane1_strm1_ready      ),      
               .std__pe2__lane1_strm1_cntl          ( std__pe2__lane1_strm1_cntl       ),      
               .std__pe2__lane1_strm1_data          ( std__pe2__lane1_strm1_data       ),      
               .std__pe2__lane1_strm1_data_valid    ( std__pe2__lane1_strm1_data_valid ),      
               .std__pe2__lane1_strm1_data_mask     ( std__pe2__lane1_strm1_data_mask  ),      

               // PE 2, Lane 2                 
               .pe2__std__lane2_strm0_ready         ( pe2__std__lane2_strm0_ready      ),      
               .std__pe2__lane2_strm0_cntl          ( std__pe2__lane2_strm0_cntl       ),      
               .std__pe2__lane2_strm0_data          ( std__pe2__lane2_strm0_data       ),      
               .std__pe2__lane2_strm0_data_valid    ( std__pe2__lane2_strm0_data_valid ),      
               .std__pe2__lane2_strm0_data_mask     ( std__pe2__lane2_strm0_data_mask  ),      

               .pe2__std__lane2_strm1_ready         ( pe2__std__lane2_strm1_ready      ),      
               .std__pe2__lane2_strm1_cntl          ( std__pe2__lane2_strm1_cntl       ),      
               .std__pe2__lane2_strm1_data          ( std__pe2__lane2_strm1_data       ),      
               .std__pe2__lane2_strm1_data_valid    ( std__pe2__lane2_strm1_data_valid ),      
               .std__pe2__lane2_strm1_data_mask     ( std__pe2__lane2_strm1_data_mask  ),      

               // PE 2, Lane 3                 
               .pe2__std__lane3_strm0_ready         ( pe2__std__lane3_strm0_ready      ),      
               .std__pe2__lane3_strm0_cntl          ( std__pe2__lane3_strm0_cntl       ),      
               .std__pe2__lane3_strm0_data          ( std__pe2__lane3_strm0_data       ),      
               .std__pe2__lane3_strm0_data_valid    ( std__pe2__lane3_strm0_data_valid ),      
               .std__pe2__lane3_strm0_data_mask     ( std__pe2__lane3_strm0_data_mask  ),      

               .pe2__std__lane3_strm1_ready         ( pe2__std__lane3_strm1_ready      ),      
               .std__pe2__lane3_strm1_cntl          ( std__pe2__lane3_strm1_cntl       ),      
               .std__pe2__lane3_strm1_data          ( std__pe2__lane3_strm1_data       ),      
               .std__pe2__lane3_strm1_data_valid    ( std__pe2__lane3_strm1_data_valid ),      
               .std__pe2__lane3_strm1_data_mask     ( std__pe2__lane3_strm1_data_mask  ),      

               // PE 2, Lane 4                 
               .pe2__std__lane4_strm0_ready         ( pe2__std__lane4_strm0_ready      ),      
               .std__pe2__lane4_strm0_cntl          ( std__pe2__lane4_strm0_cntl       ),      
               .std__pe2__lane4_strm0_data          ( std__pe2__lane4_strm0_data       ),      
               .std__pe2__lane4_strm0_data_valid    ( std__pe2__lane4_strm0_data_valid ),      
               .std__pe2__lane4_strm0_data_mask     ( std__pe2__lane4_strm0_data_mask  ),      

               .pe2__std__lane4_strm1_ready         ( pe2__std__lane4_strm1_ready      ),      
               .std__pe2__lane4_strm1_cntl          ( std__pe2__lane4_strm1_cntl       ),      
               .std__pe2__lane4_strm1_data          ( std__pe2__lane4_strm1_data       ),      
               .std__pe2__lane4_strm1_data_valid    ( std__pe2__lane4_strm1_data_valid ),      
               .std__pe2__lane4_strm1_data_mask     ( std__pe2__lane4_strm1_data_mask  ),      

               // PE 2, Lane 5                 
               .pe2__std__lane5_strm0_ready         ( pe2__std__lane5_strm0_ready      ),      
               .std__pe2__lane5_strm0_cntl          ( std__pe2__lane5_strm0_cntl       ),      
               .std__pe2__lane5_strm0_data          ( std__pe2__lane5_strm0_data       ),      
               .std__pe2__lane5_strm0_data_valid    ( std__pe2__lane5_strm0_data_valid ),      
               .std__pe2__lane5_strm0_data_mask     ( std__pe2__lane5_strm0_data_mask  ),      

               .pe2__std__lane5_strm1_ready         ( pe2__std__lane5_strm1_ready      ),      
               .std__pe2__lane5_strm1_cntl          ( std__pe2__lane5_strm1_cntl       ),      
               .std__pe2__lane5_strm1_data          ( std__pe2__lane5_strm1_data       ),      
               .std__pe2__lane5_strm1_data_valid    ( std__pe2__lane5_strm1_data_valid ),      
               .std__pe2__lane5_strm1_data_mask     ( std__pe2__lane5_strm1_data_mask  ),      

               // PE 2, Lane 6                 
               .pe2__std__lane6_strm0_ready         ( pe2__std__lane6_strm0_ready      ),      
               .std__pe2__lane6_strm0_cntl          ( std__pe2__lane6_strm0_cntl       ),      
               .std__pe2__lane6_strm0_data          ( std__pe2__lane6_strm0_data       ),      
               .std__pe2__lane6_strm0_data_valid    ( std__pe2__lane6_strm0_data_valid ),      
               .std__pe2__lane6_strm0_data_mask     ( std__pe2__lane6_strm0_data_mask  ),      

               .pe2__std__lane6_strm1_ready         ( pe2__std__lane6_strm1_ready      ),      
               .std__pe2__lane6_strm1_cntl          ( std__pe2__lane6_strm1_cntl       ),      
               .std__pe2__lane6_strm1_data          ( std__pe2__lane6_strm1_data       ),      
               .std__pe2__lane6_strm1_data_valid    ( std__pe2__lane6_strm1_data_valid ),      
               .std__pe2__lane6_strm1_data_mask     ( std__pe2__lane6_strm1_data_mask  ),      

               // PE 2, Lane 7                 
               .pe2__std__lane7_strm0_ready         ( pe2__std__lane7_strm0_ready      ),      
               .std__pe2__lane7_strm0_cntl          ( std__pe2__lane7_strm0_cntl       ),      
               .std__pe2__lane7_strm0_data          ( std__pe2__lane7_strm0_data       ),      
               .std__pe2__lane7_strm0_data_valid    ( std__pe2__lane7_strm0_data_valid ),      
               .std__pe2__lane7_strm0_data_mask     ( std__pe2__lane7_strm0_data_mask  ),      

               .pe2__std__lane7_strm1_ready         ( pe2__std__lane7_strm1_ready      ),      
               .std__pe2__lane7_strm1_cntl          ( std__pe2__lane7_strm1_cntl       ),      
               .std__pe2__lane7_strm1_data          ( std__pe2__lane7_strm1_data       ),      
               .std__pe2__lane7_strm1_data_valid    ( std__pe2__lane7_strm1_data_valid ),      
               .std__pe2__lane7_strm1_data_mask     ( std__pe2__lane7_strm1_data_mask  ),      

               // PE 2, Lane 8                 
               .pe2__std__lane8_strm0_ready         ( pe2__std__lane8_strm0_ready      ),      
               .std__pe2__lane8_strm0_cntl          ( std__pe2__lane8_strm0_cntl       ),      
               .std__pe2__lane8_strm0_data          ( std__pe2__lane8_strm0_data       ),      
               .std__pe2__lane8_strm0_data_valid    ( std__pe2__lane8_strm0_data_valid ),      
               .std__pe2__lane8_strm0_data_mask     ( std__pe2__lane8_strm0_data_mask  ),      

               .pe2__std__lane8_strm1_ready         ( pe2__std__lane8_strm1_ready      ),      
               .std__pe2__lane8_strm1_cntl          ( std__pe2__lane8_strm1_cntl       ),      
               .std__pe2__lane8_strm1_data          ( std__pe2__lane8_strm1_data       ),      
               .std__pe2__lane8_strm1_data_valid    ( std__pe2__lane8_strm1_data_valid ),      
               .std__pe2__lane8_strm1_data_mask     ( std__pe2__lane8_strm1_data_mask  ),      

               // PE 2, Lane 9                 
               .pe2__std__lane9_strm0_ready         ( pe2__std__lane9_strm0_ready      ),      
               .std__pe2__lane9_strm0_cntl          ( std__pe2__lane9_strm0_cntl       ),      
               .std__pe2__lane9_strm0_data          ( std__pe2__lane9_strm0_data       ),      
               .std__pe2__lane9_strm0_data_valid    ( std__pe2__lane9_strm0_data_valid ),      
               .std__pe2__lane9_strm0_data_mask     ( std__pe2__lane9_strm0_data_mask  ),      

               .pe2__std__lane9_strm1_ready         ( pe2__std__lane9_strm1_ready      ),      
               .std__pe2__lane9_strm1_cntl          ( std__pe2__lane9_strm1_cntl       ),      
               .std__pe2__lane9_strm1_data          ( std__pe2__lane9_strm1_data       ),      
               .std__pe2__lane9_strm1_data_valid    ( std__pe2__lane9_strm1_data_valid ),      
               .std__pe2__lane9_strm1_data_mask     ( std__pe2__lane9_strm1_data_mask  ),      

               // PE 2, Lane 10                 
               .pe2__std__lane10_strm0_ready         ( pe2__std__lane10_strm0_ready      ),      
               .std__pe2__lane10_strm0_cntl          ( std__pe2__lane10_strm0_cntl       ),      
               .std__pe2__lane10_strm0_data          ( std__pe2__lane10_strm0_data       ),      
               .std__pe2__lane10_strm0_data_valid    ( std__pe2__lane10_strm0_data_valid ),      
               .std__pe2__lane10_strm0_data_mask     ( std__pe2__lane10_strm0_data_mask  ),      

               .pe2__std__lane10_strm1_ready         ( pe2__std__lane10_strm1_ready      ),      
               .std__pe2__lane10_strm1_cntl          ( std__pe2__lane10_strm1_cntl       ),      
               .std__pe2__lane10_strm1_data          ( std__pe2__lane10_strm1_data       ),      
               .std__pe2__lane10_strm1_data_valid    ( std__pe2__lane10_strm1_data_valid ),      
               .std__pe2__lane10_strm1_data_mask     ( std__pe2__lane10_strm1_data_mask  ),      

               // PE 2, Lane 11                 
               .pe2__std__lane11_strm0_ready         ( pe2__std__lane11_strm0_ready      ),      
               .std__pe2__lane11_strm0_cntl          ( std__pe2__lane11_strm0_cntl       ),      
               .std__pe2__lane11_strm0_data          ( std__pe2__lane11_strm0_data       ),      
               .std__pe2__lane11_strm0_data_valid    ( std__pe2__lane11_strm0_data_valid ),      
               .std__pe2__lane11_strm0_data_mask     ( std__pe2__lane11_strm0_data_mask  ),      

               .pe2__std__lane11_strm1_ready         ( pe2__std__lane11_strm1_ready      ),      
               .std__pe2__lane11_strm1_cntl          ( std__pe2__lane11_strm1_cntl       ),      
               .std__pe2__lane11_strm1_data          ( std__pe2__lane11_strm1_data       ),      
               .std__pe2__lane11_strm1_data_valid    ( std__pe2__lane11_strm1_data_valid ),      
               .std__pe2__lane11_strm1_data_mask     ( std__pe2__lane11_strm1_data_mask  ),      

               // PE 2, Lane 12                 
               .pe2__std__lane12_strm0_ready         ( pe2__std__lane12_strm0_ready      ),      
               .std__pe2__lane12_strm0_cntl          ( std__pe2__lane12_strm0_cntl       ),      
               .std__pe2__lane12_strm0_data          ( std__pe2__lane12_strm0_data       ),      
               .std__pe2__lane12_strm0_data_valid    ( std__pe2__lane12_strm0_data_valid ),      
               .std__pe2__lane12_strm0_data_mask     ( std__pe2__lane12_strm0_data_mask  ),      

               .pe2__std__lane12_strm1_ready         ( pe2__std__lane12_strm1_ready      ),      
               .std__pe2__lane12_strm1_cntl          ( std__pe2__lane12_strm1_cntl       ),      
               .std__pe2__lane12_strm1_data          ( std__pe2__lane12_strm1_data       ),      
               .std__pe2__lane12_strm1_data_valid    ( std__pe2__lane12_strm1_data_valid ),      
               .std__pe2__lane12_strm1_data_mask     ( std__pe2__lane12_strm1_data_mask  ),      

               // PE 2, Lane 13                 
               .pe2__std__lane13_strm0_ready         ( pe2__std__lane13_strm0_ready      ),      
               .std__pe2__lane13_strm0_cntl          ( std__pe2__lane13_strm0_cntl       ),      
               .std__pe2__lane13_strm0_data          ( std__pe2__lane13_strm0_data       ),      
               .std__pe2__lane13_strm0_data_valid    ( std__pe2__lane13_strm0_data_valid ),      
               .std__pe2__lane13_strm0_data_mask     ( std__pe2__lane13_strm0_data_mask  ),      

               .pe2__std__lane13_strm1_ready         ( pe2__std__lane13_strm1_ready      ),      
               .std__pe2__lane13_strm1_cntl          ( std__pe2__lane13_strm1_cntl       ),      
               .std__pe2__lane13_strm1_data          ( std__pe2__lane13_strm1_data       ),      
               .std__pe2__lane13_strm1_data_valid    ( std__pe2__lane13_strm1_data_valid ),      
               .std__pe2__lane13_strm1_data_mask     ( std__pe2__lane13_strm1_data_mask  ),      

               // PE 2, Lane 14                 
               .pe2__std__lane14_strm0_ready         ( pe2__std__lane14_strm0_ready      ),      
               .std__pe2__lane14_strm0_cntl          ( std__pe2__lane14_strm0_cntl       ),      
               .std__pe2__lane14_strm0_data          ( std__pe2__lane14_strm0_data       ),      
               .std__pe2__lane14_strm0_data_valid    ( std__pe2__lane14_strm0_data_valid ),      
               .std__pe2__lane14_strm0_data_mask     ( std__pe2__lane14_strm0_data_mask  ),      

               .pe2__std__lane14_strm1_ready         ( pe2__std__lane14_strm1_ready      ),      
               .std__pe2__lane14_strm1_cntl          ( std__pe2__lane14_strm1_cntl       ),      
               .std__pe2__lane14_strm1_data          ( std__pe2__lane14_strm1_data       ),      
               .std__pe2__lane14_strm1_data_valid    ( std__pe2__lane14_strm1_data_valid ),      
               .std__pe2__lane14_strm1_data_mask     ( std__pe2__lane14_strm1_data_mask  ),      

               // PE 2, Lane 15                 
               .pe2__std__lane15_strm0_ready         ( pe2__std__lane15_strm0_ready      ),      
               .std__pe2__lane15_strm0_cntl          ( std__pe2__lane15_strm0_cntl       ),      
               .std__pe2__lane15_strm0_data          ( std__pe2__lane15_strm0_data       ),      
               .std__pe2__lane15_strm0_data_valid    ( std__pe2__lane15_strm0_data_valid ),      
               .std__pe2__lane15_strm0_data_mask     ( std__pe2__lane15_strm0_data_mask  ),      

               .pe2__std__lane15_strm1_ready         ( pe2__std__lane15_strm1_ready      ),      
               .std__pe2__lane15_strm1_cntl          ( std__pe2__lane15_strm1_cntl       ),      
               .std__pe2__lane15_strm1_data          ( std__pe2__lane15_strm1_data       ),      
               .std__pe2__lane15_strm1_data_valid    ( std__pe2__lane15_strm1_data_valid ),      
               .std__pe2__lane15_strm1_data_mask     ( std__pe2__lane15_strm1_data_mask  ),      

               // PE 2, Lane 16                 
               .pe2__std__lane16_strm0_ready         ( pe2__std__lane16_strm0_ready      ),      
               .std__pe2__lane16_strm0_cntl          ( std__pe2__lane16_strm0_cntl       ),      
               .std__pe2__lane16_strm0_data          ( std__pe2__lane16_strm0_data       ),      
               .std__pe2__lane16_strm0_data_valid    ( std__pe2__lane16_strm0_data_valid ),      
               .std__pe2__lane16_strm0_data_mask     ( std__pe2__lane16_strm0_data_mask  ),      

               .pe2__std__lane16_strm1_ready         ( pe2__std__lane16_strm1_ready      ),      
               .std__pe2__lane16_strm1_cntl          ( std__pe2__lane16_strm1_cntl       ),      
               .std__pe2__lane16_strm1_data          ( std__pe2__lane16_strm1_data       ),      
               .std__pe2__lane16_strm1_data_valid    ( std__pe2__lane16_strm1_data_valid ),      
               .std__pe2__lane16_strm1_data_mask     ( std__pe2__lane16_strm1_data_mask  ),      

               // PE 2, Lane 17                 
               .pe2__std__lane17_strm0_ready         ( pe2__std__lane17_strm0_ready      ),      
               .std__pe2__lane17_strm0_cntl          ( std__pe2__lane17_strm0_cntl       ),      
               .std__pe2__lane17_strm0_data          ( std__pe2__lane17_strm0_data       ),      
               .std__pe2__lane17_strm0_data_valid    ( std__pe2__lane17_strm0_data_valid ),      
               .std__pe2__lane17_strm0_data_mask     ( std__pe2__lane17_strm0_data_mask  ),      

               .pe2__std__lane17_strm1_ready         ( pe2__std__lane17_strm1_ready      ),      
               .std__pe2__lane17_strm1_cntl          ( std__pe2__lane17_strm1_cntl       ),      
               .std__pe2__lane17_strm1_data          ( std__pe2__lane17_strm1_data       ),      
               .std__pe2__lane17_strm1_data_valid    ( std__pe2__lane17_strm1_data_valid ),      
               .std__pe2__lane17_strm1_data_mask     ( std__pe2__lane17_strm1_data_mask  ),      

               // PE 2, Lane 18                 
               .pe2__std__lane18_strm0_ready         ( pe2__std__lane18_strm0_ready      ),      
               .std__pe2__lane18_strm0_cntl          ( std__pe2__lane18_strm0_cntl       ),      
               .std__pe2__lane18_strm0_data          ( std__pe2__lane18_strm0_data       ),      
               .std__pe2__lane18_strm0_data_valid    ( std__pe2__lane18_strm0_data_valid ),      
               .std__pe2__lane18_strm0_data_mask     ( std__pe2__lane18_strm0_data_mask  ),      

               .pe2__std__lane18_strm1_ready         ( pe2__std__lane18_strm1_ready      ),      
               .std__pe2__lane18_strm1_cntl          ( std__pe2__lane18_strm1_cntl       ),      
               .std__pe2__lane18_strm1_data          ( std__pe2__lane18_strm1_data       ),      
               .std__pe2__lane18_strm1_data_valid    ( std__pe2__lane18_strm1_data_valid ),      
               .std__pe2__lane18_strm1_data_mask     ( std__pe2__lane18_strm1_data_mask  ),      

               // PE 2, Lane 19                 
               .pe2__std__lane19_strm0_ready         ( pe2__std__lane19_strm0_ready      ),      
               .std__pe2__lane19_strm0_cntl          ( std__pe2__lane19_strm0_cntl       ),      
               .std__pe2__lane19_strm0_data          ( std__pe2__lane19_strm0_data       ),      
               .std__pe2__lane19_strm0_data_valid    ( std__pe2__lane19_strm0_data_valid ),      
               .std__pe2__lane19_strm0_data_mask     ( std__pe2__lane19_strm0_data_mask  ),      

               .pe2__std__lane19_strm1_ready         ( pe2__std__lane19_strm1_ready      ),      
               .std__pe2__lane19_strm1_cntl          ( std__pe2__lane19_strm1_cntl       ),      
               .std__pe2__lane19_strm1_data          ( std__pe2__lane19_strm1_data       ),      
               .std__pe2__lane19_strm1_data_valid    ( std__pe2__lane19_strm1_data_valid ),      
               .std__pe2__lane19_strm1_data_mask     ( std__pe2__lane19_strm1_data_mask  ),      

               // PE 2, Lane 20                 
               .pe2__std__lane20_strm0_ready         ( pe2__std__lane20_strm0_ready      ),      
               .std__pe2__lane20_strm0_cntl          ( std__pe2__lane20_strm0_cntl       ),      
               .std__pe2__lane20_strm0_data          ( std__pe2__lane20_strm0_data       ),      
               .std__pe2__lane20_strm0_data_valid    ( std__pe2__lane20_strm0_data_valid ),      
               .std__pe2__lane20_strm0_data_mask     ( std__pe2__lane20_strm0_data_mask  ),      

               .pe2__std__lane20_strm1_ready         ( pe2__std__lane20_strm1_ready      ),      
               .std__pe2__lane20_strm1_cntl          ( std__pe2__lane20_strm1_cntl       ),      
               .std__pe2__lane20_strm1_data          ( std__pe2__lane20_strm1_data       ),      
               .std__pe2__lane20_strm1_data_valid    ( std__pe2__lane20_strm1_data_valid ),      
               .std__pe2__lane20_strm1_data_mask     ( std__pe2__lane20_strm1_data_mask  ),      

               // PE 2, Lane 21                 
               .pe2__std__lane21_strm0_ready         ( pe2__std__lane21_strm0_ready      ),      
               .std__pe2__lane21_strm0_cntl          ( std__pe2__lane21_strm0_cntl       ),      
               .std__pe2__lane21_strm0_data          ( std__pe2__lane21_strm0_data       ),      
               .std__pe2__lane21_strm0_data_valid    ( std__pe2__lane21_strm0_data_valid ),      
               .std__pe2__lane21_strm0_data_mask     ( std__pe2__lane21_strm0_data_mask  ),      

               .pe2__std__lane21_strm1_ready         ( pe2__std__lane21_strm1_ready      ),      
               .std__pe2__lane21_strm1_cntl          ( std__pe2__lane21_strm1_cntl       ),      
               .std__pe2__lane21_strm1_data          ( std__pe2__lane21_strm1_data       ),      
               .std__pe2__lane21_strm1_data_valid    ( std__pe2__lane21_strm1_data_valid ),      
               .std__pe2__lane21_strm1_data_mask     ( std__pe2__lane21_strm1_data_mask  ),      

               // PE 2, Lane 22                 
               .pe2__std__lane22_strm0_ready         ( pe2__std__lane22_strm0_ready      ),      
               .std__pe2__lane22_strm0_cntl          ( std__pe2__lane22_strm0_cntl       ),      
               .std__pe2__lane22_strm0_data          ( std__pe2__lane22_strm0_data       ),      
               .std__pe2__lane22_strm0_data_valid    ( std__pe2__lane22_strm0_data_valid ),      
               .std__pe2__lane22_strm0_data_mask     ( std__pe2__lane22_strm0_data_mask  ),      

               .pe2__std__lane22_strm1_ready         ( pe2__std__lane22_strm1_ready      ),      
               .std__pe2__lane22_strm1_cntl          ( std__pe2__lane22_strm1_cntl       ),      
               .std__pe2__lane22_strm1_data          ( std__pe2__lane22_strm1_data       ),      
               .std__pe2__lane22_strm1_data_valid    ( std__pe2__lane22_strm1_data_valid ),      
               .std__pe2__lane22_strm1_data_mask     ( std__pe2__lane22_strm1_data_mask  ),      

               // PE 2, Lane 23                 
               .pe2__std__lane23_strm0_ready         ( pe2__std__lane23_strm0_ready      ),      
               .std__pe2__lane23_strm0_cntl          ( std__pe2__lane23_strm0_cntl       ),      
               .std__pe2__lane23_strm0_data          ( std__pe2__lane23_strm0_data       ),      
               .std__pe2__lane23_strm0_data_valid    ( std__pe2__lane23_strm0_data_valid ),      
               .std__pe2__lane23_strm0_data_mask     ( std__pe2__lane23_strm0_data_mask  ),      

               .pe2__std__lane23_strm1_ready         ( pe2__std__lane23_strm1_ready      ),      
               .std__pe2__lane23_strm1_cntl          ( std__pe2__lane23_strm1_cntl       ),      
               .std__pe2__lane23_strm1_data          ( std__pe2__lane23_strm1_data       ),      
               .std__pe2__lane23_strm1_data_valid    ( std__pe2__lane23_strm1_data_valid ),      
               .std__pe2__lane23_strm1_data_mask     ( std__pe2__lane23_strm1_data_mask  ),      

               // PE 2, Lane 24                 
               .pe2__std__lane24_strm0_ready         ( pe2__std__lane24_strm0_ready      ),      
               .std__pe2__lane24_strm0_cntl          ( std__pe2__lane24_strm0_cntl       ),      
               .std__pe2__lane24_strm0_data          ( std__pe2__lane24_strm0_data       ),      
               .std__pe2__lane24_strm0_data_valid    ( std__pe2__lane24_strm0_data_valid ),      
               .std__pe2__lane24_strm0_data_mask     ( std__pe2__lane24_strm0_data_mask  ),      

               .pe2__std__lane24_strm1_ready         ( pe2__std__lane24_strm1_ready      ),      
               .std__pe2__lane24_strm1_cntl          ( std__pe2__lane24_strm1_cntl       ),      
               .std__pe2__lane24_strm1_data          ( std__pe2__lane24_strm1_data       ),      
               .std__pe2__lane24_strm1_data_valid    ( std__pe2__lane24_strm1_data_valid ),      
               .std__pe2__lane24_strm1_data_mask     ( std__pe2__lane24_strm1_data_mask  ),      

               // PE 2, Lane 25                 
               .pe2__std__lane25_strm0_ready         ( pe2__std__lane25_strm0_ready      ),      
               .std__pe2__lane25_strm0_cntl          ( std__pe2__lane25_strm0_cntl       ),      
               .std__pe2__lane25_strm0_data          ( std__pe2__lane25_strm0_data       ),      
               .std__pe2__lane25_strm0_data_valid    ( std__pe2__lane25_strm0_data_valid ),      
               .std__pe2__lane25_strm0_data_mask     ( std__pe2__lane25_strm0_data_mask  ),      

               .pe2__std__lane25_strm1_ready         ( pe2__std__lane25_strm1_ready      ),      
               .std__pe2__lane25_strm1_cntl          ( std__pe2__lane25_strm1_cntl       ),      
               .std__pe2__lane25_strm1_data          ( std__pe2__lane25_strm1_data       ),      
               .std__pe2__lane25_strm1_data_valid    ( std__pe2__lane25_strm1_data_valid ),      
               .std__pe2__lane25_strm1_data_mask     ( std__pe2__lane25_strm1_data_mask  ),      

               // PE 2, Lane 26                 
               .pe2__std__lane26_strm0_ready         ( pe2__std__lane26_strm0_ready      ),      
               .std__pe2__lane26_strm0_cntl          ( std__pe2__lane26_strm0_cntl       ),      
               .std__pe2__lane26_strm0_data          ( std__pe2__lane26_strm0_data       ),      
               .std__pe2__lane26_strm0_data_valid    ( std__pe2__lane26_strm0_data_valid ),      
               .std__pe2__lane26_strm0_data_mask     ( std__pe2__lane26_strm0_data_mask  ),      

               .pe2__std__lane26_strm1_ready         ( pe2__std__lane26_strm1_ready      ),      
               .std__pe2__lane26_strm1_cntl          ( std__pe2__lane26_strm1_cntl       ),      
               .std__pe2__lane26_strm1_data          ( std__pe2__lane26_strm1_data       ),      
               .std__pe2__lane26_strm1_data_valid    ( std__pe2__lane26_strm1_data_valid ),      
               .std__pe2__lane26_strm1_data_mask     ( std__pe2__lane26_strm1_data_mask  ),      

               // PE 2, Lane 27                 
               .pe2__std__lane27_strm0_ready         ( pe2__std__lane27_strm0_ready      ),      
               .std__pe2__lane27_strm0_cntl          ( std__pe2__lane27_strm0_cntl       ),      
               .std__pe2__lane27_strm0_data          ( std__pe2__lane27_strm0_data       ),      
               .std__pe2__lane27_strm0_data_valid    ( std__pe2__lane27_strm0_data_valid ),      
               .std__pe2__lane27_strm0_data_mask     ( std__pe2__lane27_strm0_data_mask  ),      

               .pe2__std__lane27_strm1_ready         ( pe2__std__lane27_strm1_ready      ),      
               .std__pe2__lane27_strm1_cntl          ( std__pe2__lane27_strm1_cntl       ),      
               .std__pe2__lane27_strm1_data          ( std__pe2__lane27_strm1_data       ),      
               .std__pe2__lane27_strm1_data_valid    ( std__pe2__lane27_strm1_data_valid ),      
               .std__pe2__lane27_strm1_data_mask     ( std__pe2__lane27_strm1_data_mask  ),      

               // PE 2, Lane 28                 
               .pe2__std__lane28_strm0_ready         ( pe2__std__lane28_strm0_ready      ),      
               .std__pe2__lane28_strm0_cntl          ( std__pe2__lane28_strm0_cntl       ),      
               .std__pe2__lane28_strm0_data          ( std__pe2__lane28_strm0_data       ),      
               .std__pe2__lane28_strm0_data_valid    ( std__pe2__lane28_strm0_data_valid ),      
               .std__pe2__lane28_strm0_data_mask     ( std__pe2__lane28_strm0_data_mask  ),      

               .pe2__std__lane28_strm1_ready         ( pe2__std__lane28_strm1_ready      ),      
               .std__pe2__lane28_strm1_cntl          ( std__pe2__lane28_strm1_cntl       ),      
               .std__pe2__lane28_strm1_data          ( std__pe2__lane28_strm1_data       ),      
               .std__pe2__lane28_strm1_data_valid    ( std__pe2__lane28_strm1_data_valid ),      
               .std__pe2__lane28_strm1_data_mask     ( std__pe2__lane28_strm1_data_mask  ),      

               // PE 2, Lane 29                 
               .pe2__std__lane29_strm0_ready         ( pe2__std__lane29_strm0_ready      ),      
               .std__pe2__lane29_strm0_cntl          ( std__pe2__lane29_strm0_cntl       ),      
               .std__pe2__lane29_strm0_data          ( std__pe2__lane29_strm0_data       ),      
               .std__pe2__lane29_strm0_data_valid    ( std__pe2__lane29_strm0_data_valid ),      
               .std__pe2__lane29_strm0_data_mask     ( std__pe2__lane29_strm0_data_mask  ),      

               .pe2__std__lane29_strm1_ready         ( pe2__std__lane29_strm1_ready      ),      
               .std__pe2__lane29_strm1_cntl          ( std__pe2__lane29_strm1_cntl       ),      
               .std__pe2__lane29_strm1_data          ( std__pe2__lane29_strm1_data       ),      
               .std__pe2__lane29_strm1_data_valid    ( std__pe2__lane29_strm1_data_valid ),      
               .std__pe2__lane29_strm1_data_mask     ( std__pe2__lane29_strm1_data_mask  ),      

               // PE 2, Lane 30                 
               .pe2__std__lane30_strm0_ready         ( pe2__std__lane30_strm0_ready      ),      
               .std__pe2__lane30_strm0_cntl          ( std__pe2__lane30_strm0_cntl       ),      
               .std__pe2__lane30_strm0_data          ( std__pe2__lane30_strm0_data       ),      
               .std__pe2__lane30_strm0_data_valid    ( std__pe2__lane30_strm0_data_valid ),      
               .std__pe2__lane30_strm0_data_mask     ( std__pe2__lane30_strm0_data_mask  ),      

               .pe2__std__lane30_strm1_ready         ( pe2__std__lane30_strm1_ready      ),      
               .std__pe2__lane30_strm1_cntl          ( std__pe2__lane30_strm1_cntl       ),      
               .std__pe2__lane30_strm1_data          ( std__pe2__lane30_strm1_data       ),      
               .std__pe2__lane30_strm1_data_valid    ( std__pe2__lane30_strm1_data_valid ),      
               .std__pe2__lane30_strm1_data_mask     ( std__pe2__lane30_strm1_data_mask  ),      

               // PE 2, Lane 31                 
               .pe2__std__lane31_strm0_ready         ( pe2__std__lane31_strm0_ready      ),      
               .std__pe2__lane31_strm0_cntl          ( std__pe2__lane31_strm0_cntl       ),      
               .std__pe2__lane31_strm0_data          ( std__pe2__lane31_strm0_data       ),      
               .std__pe2__lane31_strm0_data_valid    ( std__pe2__lane31_strm0_data_valid ),      
               .std__pe2__lane31_strm0_data_mask     ( std__pe2__lane31_strm0_data_mask  ),      

               .pe2__std__lane31_strm1_ready         ( pe2__std__lane31_strm1_ready      ),      
               .std__pe2__lane31_strm1_cntl          ( std__pe2__lane31_strm1_cntl       ),      
               .std__pe2__lane31_strm1_data          ( std__pe2__lane31_strm1_data       ),      
               .std__pe2__lane31_strm1_data_valid    ( std__pe2__lane31_strm1_data_valid ),      
               .std__pe2__lane31_strm1_data_mask     ( std__pe2__lane31_strm1_data_mask  ),      

               // PE 3, Lane 0                 
               .pe3__std__lane0_strm0_ready         ( pe3__std__lane0_strm0_ready      ),      
               .std__pe3__lane0_strm0_cntl          ( std__pe3__lane0_strm0_cntl       ),      
               .std__pe3__lane0_strm0_data          ( std__pe3__lane0_strm0_data       ),      
               .std__pe3__lane0_strm0_data_valid    ( std__pe3__lane0_strm0_data_valid ),      
               .std__pe3__lane0_strm0_data_mask     ( std__pe3__lane0_strm0_data_mask  ),      

               .pe3__std__lane0_strm1_ready         ( pe3__std__lane0_strm1_ready      ),      
               .std__pe3__lane0_strm1_cntl          ( std__pe3__lane0_strm1_cntl       ),      
               .std__pe3__lane0_strm1_data          ( std__pe3__lane0_strm1_data       ),      
               .std__pe3__lane0_strm1_data_valid    ( std__pe3__lane0_strm1_data_valid ),      
               .std__pe3__lane0_strm1_data_mask     ( std__pe3__lane0_strm1_data_mask  ),      

               // PE 3, Lane 1                 
               .pe3__std__lane1_strm0_ready         ( pe3__std__lane1_strm0_ready      ),      
               .std__pe3__lane1_strm0_cntl          ( std__pe3__lane1_strm0_cntl       ),      
               .std__pe3__lane1_strm0_data          ( std__pe3__lane1_strm0_data       ),      
               .std__pe3__lane1_strm0_data_valid    ( std__pe3__lane1_strm0_data_valid ),      
               .std__pe3__lane1_strm0_data_mask     ( std__pe3__lane1_strm0_data_mask  ),      

               .pe3__std__lane1_strm1_ready         ( pe3__std__lane1_strm1_ready      ),      
               .std__pe3__lane1_strm1_cntl          ( std__pe3__lane1_strm1_cntl       ),      
               .std__pe3__lane1_strm1_data          ( std__pe3__lane1_strm1_data       ),      
               .std__pe3__lane1_strm1_data_valid    ( std__pe3__lane1_strm1_data_valid ),      
               .std__pe3__lane1_strm1_data_mask     ( std__pe3__lane1_strm1_data_mask  ),      

               // PE 3, Lane 2                 
               .pe3__std__lane2_strm0_ready         ( pe3__std__lane2_strm0_ready      ),      
               .std__pe3__lane2_strm0_cntl          ( std__pe3__lane2_strm0_cntl       ),      
               .std__pe3__lane2_strm0_data          ( std__pe3__lane2_strm0_data       ),      
               .std__pe3__lane2_strm0_data_valid    ( std__pe3__lane2_strm0_data_valid ),      
               .std__pe3__lane2_strm0_data_mask     ( std__pe3__lane2_strm0_data_mask  ),      

               .pe3__std__lane2_strm1_ready         ( pe3__std__lane2_strm1_ready      ),      
               .std__pe3__lane2_strm1_cntl          ( std__pe3__lane2_strm1_cntl       ),      
               .std__pe3__lane2_strm1_data          ( std__pe3__lane2_strm1_data       ),      
               .std__pe3__lane2_strm1_data_valid    ( std__pe3__lane2_strm1_data_valid ),      
               .std__pe3__lane2_strm1_data_mask     ( std__pe3__lane2_strm1_data_mask  ),      

               // PE 3, Lane 3                 
               .pe3__std__lane3_strm0_ready         ( pe3__std__lane3_strm0_ready      ),      
               .std__pe3__lane3_strm0_cntl          ( std__pe3__lane3_strm0_cntl       ),      
               .std__pe3__lane3_strm0_data          ( std__pe3__lane3_strm0_data       ),      
               .std__pe3__lane3_strm0_data_valid    ( std__pe3__lane3_strm0_data_valid ),      
               .std__pe3__lane3_strm0_data_mask     ( std__pe3__lane3_strm0_data_mask  ),      

               .pe3__std__lane3_strm1_ready         ( pe3__std__lane3_strm1_ready      ),      
               .std__pe3__lane3_strm1_cntl          ( std__pe3__lane3_strm1_cntl       ),      
               .std__pe3__lane3_strm1_data          ( std__pe3__lane3_strm1_data       ),      
               .std__pe3__lane3_strm1_data_valid    ( std__pe3__lane3_strm1_data_valid ),      
               .std__pe3__lane3_strm1_data_mask     ( std__pe3__lane3_strm1_data_mask  ),      

               // PE 3, Lane 4                 
               .pe3__std__lane4_strm0_ready         ( pe3__std__lane4_strm0_ready      ),      
               .std__pe3__lane4_strm0_cntl          ( std__pe3__lane4_strm0_cntl       ),      
               .std__pe3__lane4_strm0_data          ( std__pe3__lane4_strm0_data       ),      
               .std__pe3__lane4_strm0_data_valid    ( std__pe3__lane4_strm0_data_valid ),      
               .std__pe3__lane4_strm0_data_mask     ( std__pe3__lane4_strm0_data_mask  ),      

               .pe3__std__lane4_strm1_ready         ( pe3__std__lane4_strm1_ready      ),      
               .std__pe3__lane4_strm1_cntl          ( std__pe3__lane4_strm1_cntl       ),      
               .std__pe3__lane4_strm1_data          ( std__pe3__lane4_strm1_data       ),      
               .std__pe3__lane4_strm1_data_valid    ( std__pe3__lane4_strm1_data_valid ),      
               .std__pe3__lane4_strm1_data_mask     ( std__pe3__lane4_strm1_data_mask  ),      

               // PE 3, Lane 5                 
               .pe3__std__lane5_strm0_ready         ( pe3__std__lane5_strm0_ready      ),      
               .std__pe3__lane5_strm0_cntl          ( std__pe3__lane5_strm0_cntl       ),      
               .std__pe3__lane5_strm0_data          ( std__pe3__lane5_strm0_data       ),      
               .std__pe3__lane5_strm0_data_valid    ( std__pe3__lane5_strm0_data_valid ),      
               .std__pe3__lane5_strm0_data_mask     ( std__pe3__lane5_strm0_data_mask  ),      

               .pe3__std__lane5_strm1_ready         ( pe3__std__lane5_strm1_ready      ),      
               .std__pe3__lane5_strm1_cntl          ( std__pe3__lane5_strm1_cntl       ),      
               .std__pe3__lane5_strm1_data          ( std__pe3__lane5_strm1_data       ),      
               .std__pe3__lane5_strm1_data_valid    ( std__pe3__lane5_strm1_data_valid ),      
               .std__pe3__lane5_strm1_data_mask     ( std__pe3__lane5_strm1_data_mask  ),      

               // PE 3, Lane 6                 
               .pe3__std__lane6_strm0_ready         ( pe3__std__lane6_strm0_ready      ),      
               .std__pe3__lane6_strm0_cntl          ( std__pe3__lane6_strm0_cntl       ),      
               .std__pe3__lane6_strm0_data          ( std__pe3__lane6_strm0_data       ),      
               .std__pe3__lane6_strm0_data_valid    ( std__pe3__lane6_strm0_data_valid ),      
               .std__pe3__lane6_strm0_data_mask     ( std__pe3__lane6_strm0_data_mask  ),      

               .pe3__std__lane6_strm1_ready         ( pe3__std__lane6_strm1_ready      ),      
               .std__pe3__lane6_strm1_cntl          ( std__pe3__lane6_strm1_cntl       ),      
               .std__pe3__lane6_strm1_data          ( std__pe3__lane6_strm1_data       ),      
               .std__pe3__lane6_strm1_data_valid    ( std__pe3__lane6_strm1_data_valid ),      
               .std__pe3__lane6_strm1_data_mask     ( std__pe3__lane6_strm1_data_mask  ),      

               // PE 3, Lane 7                 
               .pe3__std__lane7_strm0_ready         ( pe3__std__lane7_strm0_ready      ),      
               .std__pe3__lane7_strm0_cntl          ( std__pe3__lane7_strm0_cntl       ),      
               .std__pe3__lane7_strm0_data          ( std__pe3__lane7_strm0_data       ),      
               .std__pe3__lane7_strm0_data_valid    ( std__pe3__lane7_strm0_data_valid ),      
               .std__pe3__lane7_strm0_data_mask     ( std__pe3__lane7_strm0_data_mask  ),      

               .pe3__std__lane7_strm1_ready         ( pe3__std__lane7_strm1_ready      ),      
               .std__pe3__lane7_strm1_cntl          ( std__pe3__lane7_strm1_cntl       ),      
               .std__pe3__lane7_strm1_data          ( std__pe3__lane7_strm1_data       ),      
               .std__pe3__lane7_strm1_data_valid    ( std__pe3__lane7_strm1_data_valid ),      
               .std__pe3__lane7_strm1_data_mask     ( std__pe3__lane7_strm1_data_mask  ),      

               // PE 3, Lane 8                 
               .pe3__std__lane8_strm0_ready         ( pe3__std__lane8_strm0_ready      ),      
               .std__pe3__lane8_strm0_cntl          ( std__pe3__lane8_strm0_cntl       ),      
               .std__pe3__lane8_strm0_data          ( std__pe3__lane8_strm0_data       ),      
               .std__pe3__lane8_strm0_data_valid    ( std__pe3__lane8_strm0_data_valid ),      
               .std__pe3__lane8_strm0_data_mask     ( std__pe3__lane8_strm0_data_mask  ),      

               .pe3__std__lane8_strm1_ready         ( pe3__std__lane8_strm1_ready      ),      
               .std__pe3__lane8_strm1_cntl          ( std__pe3__lane8_strm1_cntl       ),      
               .std__pe3__lane8_strm1_data          ( std__pe3__lane8_strm1_data       ),      
               .std__pe3__lane8_strm1_data_valid    ( std__pe3__lane8_strm1_data_valid ),      
               .std__pe3__lane8_strm1_data_mask     ( std__pe3__lane8_strm1_data_mask  ),      

               // PE 3, Lane 9                 
               .pe3__std__lane9_strm0_ready         ( pe3__std__lane9_strm0_ready      ),      
               .std__pe3__lane9_strm0_cntl          ( std__pe3__lane9_strm0_cntl       ),      
               .std__pe3__lane9_strm0_data          ( std__pe3__lane9_strm0_data       ),      
               .std__pe3__lane9_strm0_data_valid    ( std__pe3__lane9_strm0_data_valid ),      
               .std__pe3__lane9_strm0_data_mask     ( std__pe3__lane9_strm0_data_mask  ),      

               .pe3__std__lane9_strm1_ready         ( pe3__std__lane9_strm1_ready      ),      
               .std__pe3__lane9_strm1_cntl          ( std__pe3__lane9_strm1_cntl       ),      
               .std__pe3__lane9_strm1_data          ( std__pe3__lane9_strm1_data       ),      
               .std__pe3__lane9_strm1_data_valid    ( std__pe3__lane9_strm1_data_valid ),      
               .std__pe3__lane9_strm1_data_mask     ( std__pe3__lane9_strm1_data_mask  ),      

               // PE 3, Lane 10                 
               .pe3__std__lane10_strm0_ready         ( pe3__std__lane10_strm0_ready      ),      
               .std__pe3__lane10_strm0_cntl          ( std__pe3__lane10_strm0_cntl       ),      
               .std__pe3__lane10_strm0_data          ( std__pe3__lane10_strm0_data       ),      
               .std__pe3__lane10_strm0_data_valid    ( std__pe3__lane10_strm0_data_valid ),      
               .std__pe3__lane10_strm0_data_mask     ( std__pe3__lane10_strm0_data_mask  ),      

               .pe3__std__lane10_strm1_ready         ( pe3__std__lane10_strm1_ready      ),      
               .std__pe3__lane10_strm1_cntl          ( std__pe3__lane10_strm1_cntl       ),      
               .std__pe3__lane10_strm1_data          ( std__pe3__lane10_strm1_data       ),      
               .std__pe3__lane10_strm1_data_valid    ( std__pe3__lane10_strm1_data_valid ),      
               .std__pe3__lane10_strm1_data_mask     ( std__pe3__lane10_strm1_data_mask  ),      

               // PE 3, Lane 11                 
               .pe3__std__lane11_strm0_ready         ( pe3__std__lane11_strm0_ready      ),      
               .std__pe3__lane11_strm0_cntl          ( std__pe3__lane11_strm0_cntl       ),      
               .std__pe3__lane11_strm0_data          ( std__pe3__lane11_strm0_data       ),      
               .std__pe3__lane11_strm0_data_valid    ( std__pe3__lane11_strm0_data_valid ),      
               .std__pe3__lane11_strm0_data_mask     ( std__pe3__lane11_strm0_data_mask  ),      

               .pe3__std__lane11_strm1_ready         ( pe3__std__lane11_strm1_ready      ),      
               .std__pe3__lane11_strm1_cntl          ( std__pe3__lane11_strm1_cntl       ),      
               .std__pe3__lane11_strm1_data          ( std__pe3__lane11_strm1_data       ),      
               .std__pe3__lane11_strm1_data_valid    ( std__pe3__lane11_strm1_data_valid ),      
               .std__pe3__lane11_strm1_data_mask     ( std__pe3__lane11_strm1_data_mask  ),      

               // PE 3, Lane 12                 
               .pe3__std__lane12_strm0_ready         ( pe3__std__lane12_strm0_ready      ),      
               .std__pe3__lane12_strm0_cntl          ( std__pe3__lane12_strm0_cntl       ),      
               .std__pe3__lane12_strm0_data          ( std__pe3__lane12_strm0_data       ),      
               .std__pe3__lane12_strm0_data_valid    ( std__pe3__lane12_strm0_data_valid ),      
               .std__pe3__lane12_strm0_data_mask     ( std__pe3__lane12_strm0_data_mask  ),      

               .pe3__std__lane12_strm1_ready         ( pe3__std__lane12_strm1_ready      ),      
               .std__pe3__lane12_strm1_cntl          ( std__pe3__lane12_strm1_cntl       ),      
               .std__pe3__lane12_strm1_data          ( std__pe3__lane12_strm1_data       ),      
               .std__pe3__lane12_strm1_data_valid    ( std__pe3__lane12_strm1_data_valid ),      
               .std__pe3__lane12_strm1_data_mask     ( std__pe3__lane12_strm1_data_mask  ),      

               // PE 3, Lane 13                 
               .pe3__std__lane13_strm0_ready         ( pe3__std__lane13_strm0_ready      ),      
               .std__pe3__lane13_strm0_cntl          ( std__pe3__lane13_strm0_cntl       ),      
               .std__pe3__lane13_strm0_data          ( std__pe3__lane13_strm0_data       ),      
               .std__pe3__lane13_strm0_data_valid    ( std__pe3__lane13_strm0_data_valid ),      
               .std__pe3__lane13_strm0_data_mask     ( std__pe3__lane13_strm0_data_mask  ),      

               .pe3__std__lane13_strm1_ready         ( pe3__std__lane13_strm1_ready      ),      
               .std__pe3__lane13_strm1_cntl          ( std__pe3__lane13_strm1_cntl       ),      
               .std__pe3__lane13_strm1_data          ( std__pe3__lane13_strm1_data       ),      
               .std__pe3__lane13_strm1_data_valid    ( std__pe3__lane13_strm1_data_valid ),      
               .std__pe3__lane13_strm1_data_mask     ( std__pe3__lane13_strm1_data_mask  ),      

               // PE 3, Lane 14                 
               .pe3__std__lane14_strm0_ready         ( pe3__std__lane14_strm0_ready      ),      
               .std__pe3__lane14_strm0_cntl          ( std__pe3__lane14_strm0_cntl       ),      
               .std__pe3__lane14_strm0_data          ( std__pe3__lane14_strm0_data       ),      
               .std__pe3__lane14_strm0_data_valid    ( std__pe3__lane14_strm0_data_valid ),      
               .std__pe3__lane14_strm0_data_mask     ( std__pe3__lane14_strm0_data_mask  ),      

               .pe3__std__lane14_strm1_ready         ( pe3__std__lane14_strm1_ready      ),      
               .std__pe3__lane14_strm1_cntl          ( std__pe3__lane14_strm1_cntl       ),      
               .std__pe3__lane14_strm1_data          ( std__pe3__lane14_strm1_data       ),      
               .std__pe3__lane14_strm1_data_valid    ( std__pe3__lane14_strm1_data_valid ),      
               .std__pe3__lane14_strm1_data_mask     ( std__pe3__lane14_strm1_data_mask  ),      

               // PE 3, Lane 15                 
               .pe3__std__lane15_strm0_ready         ( pe3__std__lane15_strm0_ready      ),      
               .std__pe3__lane15_strm0_cntl          ( std__pe3__lane15_strm0_cntl       ),      
               .std__pe3__lane15_strm0_data          ( std__pe3__lane15_strm0_data       ),      
               .std__pe3__lane15_strm0_data_valid    ( std__pe3__lane15_strm0_data_valid ),      
               .std__pe3__lane15_strm0_data_mask     ( std__pe3__lane15_strm0_data_mask  ),      

               .pe3__std__lane15_strm1_ready         ( pe3__std__lane15_strm1_ready      ),      
               .std__pe3__lane15_strm1_cntl          ( std__pe3__lane15_strm1_cntl       ),      
               .std__pe3__lane15_strm1_data          ( std__pe3__lane15_strm1_data       ),      
               .std__pe3__lane15_strm1_data_valid    ( std__pe3__lane15_strm1_data_valid ),      
               .std__pe3__lane15_strm1_data_mask     ( std__pe3__lane15_strm1_data_mask  ),      

               // PE 3, Lane 16                 
               .pe3__std__lane16_strm0_ready         ( pe3__std__lane16_strm0_ready      ),      
               .std__pe3__lane16_strm0_cntl          ( std__pe3__lane16_strm0_cntl       ),      
               .std__pe3__lane16_strm0_data          ( std__pe3__lane16_strm0_data       ),      
               .std__pe3__lane16_strm0_data_valid    ( std__pe3__lane16_strm0_data_valid ),      
               .std__pe3__lane16_strm0_data_mask     ( std__pe3__lane16_strm0_data_mask  ),      

               .pe3__std__lane16_strm1_ready         ( pe3__std__lane16_strm1_ready      ),      
               .std__pe3__lane16_strm1_cntl          ( std__pe3__lane16_strm1_cntl       ),      
               .std__pe3__lane16_strm1_data          ( std__pe3__lane16_strm1_data       ),      
               .std__pe3__lane16_strm1_data_valid    ( std__pe3__lane16_strm1_data_valid ),      
               .std__pe3__lane16_strm1_data_mask     ( std__pe3__lane16_strm1_data_mask  ),      

               // PE 3, Lane 17                 
               .pe3__std__lane17_strm0_ready         ( pe3__std__lane17_strm0_ready      ),      
               .std__pe3__lane17_strm0_cntl          ( std__pe3__lane17_strm0_cntl       ),      
               .std__pe3__lane17_strm0_data          ( std__pe3__lane17_strm0_data       ),      
               .std__pe3__lane17_strm0_data_valid    ( std__pe3__lane17_strm0_data_valid ),      
               .std__pe3__lane17_strm0_data_mask     ( std__pe3__lane17_strm0_data_mask  ),      

               .pe3__std__lane17_strm1_ready         ( pe3__std__lane17_strm1_ready      ),      
               .std__pe3__lane17_strm1_cntl          ( std__pe3__lane17_strm1_cntl       ),      
               .std__pe3__lane17_strm1_data          ( std__pe3__lane17_strm1_data       ),      
               .std__pe3__lane17_strm1_data_valid    ( std__pe3__lane17_strm1_data_valid ),      
               .std__pe3__lane17_strm1_data_mask     ( std__pe3__lane17_strm1_data_mask  ),      

               // PE 3, Lane 18                 
               .pe3__std__lane18_strm0_ready         ( pe3__std__lane18_strm0_ready      ),      
               .std__pe3__lane18_strm0_cntl          ( std__pe3__lane18_strm0_cntl       ),      
               .std__pe3__lane18_strm0_data          ( std__pe3__lane18_strm0_data       ),      
               .std__pe3__lane18_strm0_data_valid    ( std__pe3__lane18_strm0_data_valid ),      
               .std__pe3__lane18_strm0_data_mask     ( std__pe3__lane18_strm0_data_mask  ),      

               .pe3__std__lane18_strm1_ready         ( pe3__std__lane18_strm1_ready      ),      
               .std__pe3__lane18_strm1_cntl          ( std__pe3__lane18_strm1_cntl       ),      
               .std__pe3__lane18_strm1_data          ( std__pe3__lane18_strm1_data       ),      
               .std__pe3__lane18_strm1_data_valid    ( std__pe3__lane18_strm1_data_valid ),      
               .std__pe3__lane18_strm1_data_mask     ( std__pe3__lane18_strm1_data_mask  ),      

               // PE 3, Lane 19                 
               .pe3__std__lane19_strm0_ready         ( pe3__std__lane19_strm0_ready      ),      
               .std__pe3__lane19_strm0_cntl          ( std__pe3__lane19_strm0_cntl       ),      
               .std__pe3__lane19_strm0_data          ( std__pe3__lane19_strm0_data       ),      
               .std__pe3__lane19_strm0_data_valid    ( std__pe3__lane19_strm0_data_valid ),      
               .std__pe3__lane19_strm0_data_mask     ( std__pe3__lane19_strm0_data_mask  ),      

               .pe3__std__lane19_strm1_ready         ( pe3__std__lane19_strm1_ready      ),      
               .std__pe3__lane19_strm1_cntl          ( std__pe3__lane19_strm1_cntl       ),      
               .std__pe3__lane19_strm1_data          ( std__pe3__lane19_strm1_data       ),      
               .std__pe3__lane19_strm1_data_valid    ( std__pe3__lane19_strm1_data_valid ),      
               .std__pe3__lane19_strm1_data_mask     ( std__pe3__lane19_strm1_data_mask  ),      

               // PE 3, Lane 20                 
               .pe3__std__lane20_strm0_ready         ( pe3__std__lane20_strm0_ready      ),      
               .std__pe3__lane20_strm0_cntl          ( std__pe3__lane20_strm0_cntl       ),      
               .std__pe3__lane20_strm0_data          ( std__pe3__lane20_strm0_data       ),      
               .std__pe3__lane20_strm0_data_valid    ( std__pe3__lane20_strm0_data_valid ),      
               .std__pe3__lane20_strm0_data_mask     ( std__pe3__lane20_strm0_data_mask  ),      

               .pe3__std__lane20_strm1_ready         ( pe3__std__lane20_strm1_ready      ),      
               .std__pe3__lane20_strm1_cntl          ( std__pe3__lane20_strm1_cntl       ),      
               .std__pe3__lane20_strm1_data          ( std__pe3__lane20_strm1_data       ),      
               .std__pe3__lane20_strm1_data_valid    ( std__pe3__lane20_strm1_data_valid ),      
               .std__pe3__lane20_strm1_data_mask     ( std__pe3__lane20_strm1_data_mask  ),      

               // PE 3, Lane 21                 
               .pe3__std__lane21_strm0_ready         ( pe3__std__lane21_strm0_ready      ),      
               .std__pe3__lane21_strm0_cntl          ( std__pe3__lane21_strm0_cntl       ),      
               .std__pe3__lane21_strm0_data          ( std__pe3__lane21_strm0_data       ),      
               .std__pe3__lane21_strm0_data_valid    ( std__pe3__lane21_strm0_data_valid ),      
               .std__pe3__lane21_strm0_data_mask     ( std__pe3__lane21_strm0_data_mask  ),      

               .pe3__std__lane21_strm1_ready         ( pe3__std__lane21_strm1_ready      ),      
               .std__pe3__lane21_strm1_cntl          ( std__pe3__lane21_strm1_cntl       ),      
               .std__pe3__lane21_strm1_data          ( std__pe3__lane21_strm1_data       ),      
               .std__pe3__lane21_strm1_data_valid    ( std__pe3__lane21_strm1_data_valid ),      
               .std__pe3__lane21_strm1_data_mask     ( std__pe3__lane21_strm1_data_mask  ),      

               // PE 3, Lane 22                 
               .pe3__std__lane22_strm0_ready         ( pe3__std__lane22_strm0_ready      ),      
               .std__pe3__lane22_strm0_cntl          ( std__pe3__lane22_strm0_cntl       ),      
               .std__pe3__lane22_strm0_data          ( std__pe3__lane22_strm0_data       ),      
               .std__pe3__lane22_strm0_data_valid    ( std__pe3__lane22_strm0_data_valid ),      
               .std__pe3__lane22_strm0_data_mask     ( std__pe3__lane22_strm0_data_mask  ),      

               .pe3__std__lane22_strm1_ready         ( pe3__std__lane22_strm1_ready      ),      
               .std__pe3__lane22_strm1_cntl          ( std__pe3__lane22_strm1_cntl       ),      
               .std__pe3__lane22_strm1_data          ( std__pe3__lane22_strm1_data       ),      
               .std__pe3__lane22_strm1_data_valid    ( std__pe3__lane22_strm1_data_valid ),      
               .std__pe3__lane22_strm1_data_mask     ( std__pe3__lane22_strm1_data_mask  ),      

               // PE 3, Lane 23                 
               .pe3__std__lane23_strm0_ready         ( pe3__std__lane23_strm0_ready      ),      
               .std__pe3__lane23_strm0_cntl          ( std__pe3__lane23_strm0_cntl       ),      
               .std__pe3__lane23_strm0_data          ( std__pe3__lane23_strm0_data       ),      
               .std__pe3__lane23_strm0_data_valid    ( std__pe3__lane23_strm0_data_valid ),      
               .std__pe3__lane23_strm0_data_mask     ( std__pe3__lane23_strm0_data_mask  ),      

               .pe3__std__lane23_strm1_ready         ( pe3__std__lane23_strm1_ready      ),      
               .std__pe3__lane23_strm1_cntl          ( std__pe3__lane23_strm1_cntl       ),      
               .std__pe3__lane23_strm1_data          ( std__pe3__lane23_strm1_data       ),      
               .std__pe3__lane23_strm1_data_valid    ( std__pe3__lane23_strm1_data_valid ),      
               .std__pe3__lane23_strm1_data_mask     ( std__pe3__lane23_strm1_data_mask  ),      

               // PE 3, Lane 24                 
               .pe3__std__lane24_strm0_ready         ( pe3__std__lane24_strm0_ready      ),      
               .std__pe3__lane24_strm0_cntl          ( std__pe3__lane24_strm0_cntl       ),      
               .std__pe3__lane24_strm0_data          ( std__pe3__lane24_strm0_data       ),      
               .std__pe3__lane24_strm0_data_valid    ( std__pe3__lane24_strm0_data_valid ),      
               .std__pe3__lane24_strm0_data_mask     ( std__pe3__lane24_strm0_data_mask  ),      

               .pe3__std__lane24_strm1_ready         ( pe3__std__lane24_strm1_ready      ),      
               .std__pe3__lane24_strm1_cntl          ( std__pe3__lane24_strm1_cntl       ),      
               .std__pe3__lane24_strm1_data          ( std__pe3__lane24_strm1_data       ),      
               .std__pe3__lane24_strm1_data_valid    ( std__pe3__lane24_strm1_data_valid ),      
               .std__pe3__lane24_strm1_data_mask     ( std__pe3__lane24_strm1_data_mask  ),      

               // PE 3, Lane 25                 
               .pe3__std__lane25_strm0_ready         ( pe3__std__lane25_strm0_ready      ),      
               .std__pe3__lane25_strm0_cntl          ( std__pe3__lane25_strm0_cntl       ),      
               .std__pe3__lane25_strm0_data          ( std__pe3__lane25_strm0_data       ),      
               .std__pe3__lane25_strm0_data_valid    ( std__pe3__lane25_strm0_data_valid ),      
               .std__pe3__lane25_strm0_data_mask     ( std__pe3__lane25_strm0_data_mask  ),      

               .pe3__std__lane25_strm1_ready         ( pe3__std__lane25_strm1_ready      ),      
               .std__pe3__lane25_strm1_cntl          ( std__pe3__lane25_strm1_cntl       ),      
               .std__pe3__lane25_strm1_data          ( std__pe3__lane25_strm1_data       ),      
               .std__pe3__lane25_strm1_data_valid    ( std__pe3__lane25_strm1_data_valid ),      
               .std__pe3__lane25_strm1_data_mask     ( std__pe3__lane25_strm1_data_mask  ),      

               // PE 3, Lane 26                 
               .pe3__std__lane26_strm0_ready         ( pe3__std__lane26_strm0_ready      ),      
               .std__pe3__lane26_strm0_cntl          ( std__pe3__lane26_strm0_cntl       ),      
               .std__pe3__lane26_strm0_data          ( std__pe3__lane26_strm0_data       ),      
               .std__pe3__lane26_strm0_data_valid    ( std__pe3__lane26_strm0_data_valid ),      
               .std__pe3__lane26_strm0_data_mask     ( std__pe3__lane26_strm0_data_mask  ),      

               .pe3__std__lane26_strm1_ready         ( pe3__std__lane26_strm1_ready      ),      
               .std__pe3__lane26_strm1_cntl          ( std__pe3__lane26_strm1_cntl       ),      
               .std__pe3__lane26_strm1_data          ( std__pe3__lane26_strm1_data       ),      
               .std__pe3__lane26_strm1_data_valid    ( std__pe3__lane26_strm1_data_valid ),      
               .std__pe3__lane26_strm1_data_mask     ( std__pe3__lane26_strm1_data_mask  ),      

               // PE 3, Lane 27                 
               .pe3__std__lane27_strm0_ready         ( pe3__std__lane27_strm0_ready      ),      
               .std__pe3__lane27_strm0_cntl          ( std__pe3__lane27_strm0_cntl       ),      
               .std__pe3__lane27_strm0_data          ( std__pe3__lane27_strm0_data       ),      
               .std__pe3__lane27_strm0_data_valid    ( std__pe3__lane27_strm0_data_valid ),      
               .std__pe3__lane27_strm0_data_mask     ( std__pe3__lane27_strm0_data_mask  ),      

               .pe3__std__lane27_strm1_ready         ( pe3__std__lane27_strm1_ready      ),      
               .std__pe3__lane27_strm1_cntl          ( std__pe3__lane27_strm1_cntl       ),      
               .std__pe3__lane27_strm1_data          ( std__pe3__lane27_strm1_data       ),      
               .std__pe3__lane27_strm1_data_valid    ( std__pe3__lane27_strm1_data_valid ),      
               .std__pe3__lane27_strm1_data_mask     ( std__pe3__lane27_strm1_data_mask  ),      

               // PE 3, Lane 28                 
               .pe3__std__lane28_strm0_ready         ( pe3__std__lane28_strm0_ready      ),      
               .std__pe3__lane28_strm0_cntl          ( std__pe3__lane28_strm0_cntl       ),      
               .std__pe3__lane28_strm0_data          ( std__pe3__lane28_strm0_data       ),      
               .std__pe3__lane28_strm0_data_valid    ( std__pe3__lane28_strm0_data_valid ),      
               .std__pe3__lane28_strm0_data_mask     ( std__pe3__lane28_strm0_data_mask  ),      

               .pe3__std__lane28_strm1_ready         ( pe3__std__lane28_strm1_ready      ),      
               .std__pe3__lane28_strm1_cntl          ( std__pe3__lane28_strm1_cntl       ),      
               .std__pe3__lane28_strm1_data          ( std__pe3__lane28_strm1_data       ),      
               .std__pe3__lane28_strm1_data_valid    ( std__pe3__lane28_strm1_data_valid ),      
               .std__pe3__lane28_strm1_data_mask     ( std__pe3__lane28_strm1_data_mask  ),      

               // PE 3, Lane 29                 
               .pe3__std__lane29_strm0_ready         ( pe3__std__lane29_strm0_ready      ),      
               .std__pe3__lane29_strm0_cntl          ( std__pe3__lane29_strm0_cntl       ),      
               .std__pe3__lane29_strm0_data          ( std__pe3__lane29_strm0_data       ),      
               .std__pe3__lane29_strm0_data_valid    ( std__pe3__lane29_strm0_data_valid ),      
               .std__pe3__lane29_strm0_data_mask     ( std__pe3__lane29_strm0_data_mask  ),      

               .pe3__std__lane29_strm1_ready         ( pe3__std__lane29_strm1_ready      ),      
               .std__pe3__lane29_strm1_cntl          ( std__pe3__lane29_strm1_cntl       ),      
               .std__pe3__lane29_strm1_data          ( std__pe3__lane29_strm1_data       ),      
               .std__pe3__lane29_strm1_data_valid    ( std__pe3__lane29_strm1_data_valid ),      
               .std__pe3__lane29_strm1_data_mask     ( std__pe3__lane29_strm1_data_mask  ),      

               // PE 3, Lane 30                 
               .pe3__std__lane30_strm0_ready         ( pe3__std__lane30_strm0_ready      ),      
               .std__pe3__lane30_strm0_cntl          ( std__pe3__lane30_strm0_cntl       ),      
               .std__pe3__lane30_strm0_data          ( std__pe3__lane30_strm0_data       ),      
               .std__pe3__lane30_strm0_data_valid    ( std__pe3__lane30_strm0_data_valid ),      
               .std__pe3__lane30_strm0_data_mask     ( std__pe3__lane30_strm0_data_mask  ),      

               .pe3__std__lane30_strm1_ready         ( pe3__std__lane30_strm1_ready      ),      
               .std__pe3__lane30_strm1_cntl          ( std__pe3__lane30_strm1_cntl       ),      
               .std__pe3__lane30_strm1_data          ( std__pe3__lane30_strm1_data       ),      
               .std__pe3__lane30_strm1_data_valid    ( std__pe3__lane30_strm1_data_valid ),      
               .std__pe3__lane30_strm1_data_mask     ( std__pe3__lane30_strm1_data_mask  ),      

               // PE 3, Lane 31                 
               .pe3__std__lane31_strm0_ready         ( pe3__std__lane31_strm0_ready      ),      
               .std__pe3__lane31_strm0_cntl          ( std__pe3__lane31_strm0_cntl       ),      
               .std__pe3__lane31_strm0_data          ( std__pe3__lane31_strm0_data       ),      
               .std__pe3__lane31_strm0_data_valid    ( std__pe3__lane31_strm0_data_valid ),      
               .std__pe3__lane31_strm0_data_mask     ( std__pe3__lane31_strm0_data_mask  ),      

               .pe3__std__lane31_strm1_ready         ( pe3__std__lane31_strm1_ready      ),      
               .std__pe3__lane31_strm1_cntl          ( std__pe3__lane31_strm1_cntl       ),      
               .std__pe3__lane31_strm1_data          ( std__pe3__lane31_strm1_data       ),      
               .std__pe3__lane31_strm1_data_valid    ( std__pe3__lane31_strm1_data_valid ),      
               .std__pe3__lane31_strm1_data_mask     ( std__pe3__lane31_strm1_data_mask  ),      

               // PE 4, Lane 0                 
               .pe4__std__lane0_strm0_ready         ( pe4__std__lane0_strm0_ready      ),      
               .std__pe4__lane0_strm0_cntl          ( std__pe4__lane0_strm0_cntl       ),      
               .std__pe4__lane0_strm0_data          ( std__pe4__lane0_strm0_data       ),      
               .std__pe4__lane0_strm0_data_valid    ( std__pe4__lane0_strm0_data_valid ),      
               .std__pe4__lane0_strm0_data_mask     ( std__pe4__lane0_strm0_data_mask  ),      

               .pe4__std__lane0_strm1_ready         ( pe4__std__lane0_strm1_ready      ),      
               .std__pe4__lane0_strm1_cntl          ( std__pe4__lane0_strm1_cntl       ),      
               .std__pe4__lane0_strm1_data          ( std__pe4__lane0_strm1_data       ),      
               .std__pe4__lane0_strm1_data_valid    ( std__pe4__lane0_strm1_data_valid ),      
               .std__pe4__lane0_strm1_data_mask     ( std__pe4__lane0_strm1_data_mask  ),      

               // PE 4, Lane 1                 
               .pe4__std__lane1_strm0_ready         ( pe4__std__lane1_strm0_ready      ),      
               .std__pe4__lane1_strm0_cntl          ( std__pe4__lane1_strm0_cntl       ),      
               .std__pe4__lane1_strm0_data          ( std__pe4__lane1_strm0_data       ),      
               .std__pe4__lane1_strm0_data_valid    ( std__pe4__lane1_strm0_data_valid ),      
               .std__pe4__lane1_strm0_data_mask     ( std__pe4__lane1_strm0_data_mask  ),      

               .pe4__std__lane1_strm1_ready         ( pe4__std__lane1_strm1_ready      ),      
               .std__pe4__lane1_strm1_cntl          ( std__pe4__lane1_strm1_cntl       ),      
               .std__pe4__lane1_strm1_data          ( std__pe4__lane1_strm1_data       ),      
               .std__pe4__lane1_strm1_data_valid    ( std__pe4__lane1_strm1_data_valid ),      
               .std__pe4__lane1_strm1_data_mask     ( std__pe4__lane1_strm1_data_mask  ),      

               // PE 4, Lane 2                 
               .pe4__std__lane2_strm0_ready         ( pe4__std__lane2_strm0_ready      ),      
               .std__pe4__lane2_strm0_cntl          ( std__pe4__lane2_strm0_cntl       ),      
               .std__pe4__lane2_strm0_data          ( std__pe4__lane2_strm0_data       ),      
               .std__pe4__lane2_strm0_data_valid    ( std__pe4__lane2_strm0_data_valid ),      
               .std__pe4__lane2_strm0_data_mask     ( std__pe4__lane2_strm0_data_mask  ),      

               .pe4__std__lane2_strm1_ready         ( pe4__std__lane2_strm1_ready      ),      
               .std__pe4__lane2_strm1_cntl          ( std__pe4__lane2_strm1_cntl       ),      
               .std__pe4__lane2_strm1_data          ( std__pe4__lane2_strm1_data       ),      
               .std__pe4__lane2_strm1_data_valid    ( std__pe4__lane2_strm1_data_valid ),      
               .std__pe4__lane2_strm1_data_mask     ( std__pe4__lane2_strm1_data_mask  ),      

               // PE 4, Lane 3                 
               .pe4__std__lane3_strm0_ready         ( pe4__std__lane3_strm0_ready      ),      
               .std__pe4__lane3_strm0_cntl          ( std__pe4__lane3_strm0_cntl       ),      
               .std__pe4__lane3_strm0_data          ( std__pe4__lane3_strm0_data       ),      
               .std__pe4__lane3_strm0_data_valid    ( std__pe4__lane3_strm0_data_valid ),      
               .std__pe4__lane3_strm0_data_mask     ( std__pe4__lane3_strm0_data_mask  ),      

               .pe4__std__lane3_strm1_ready         ( pe4__std__lane3_strm1_ready      ),      
               .std__pe4__lane3_strm1_cntl          ( std__pe4__lane3_strm1_cntl       ),      
               .std__pe4__lane3_strm1_data          ( std__pe4__lane3_strm1_data       ),      
               .std__pe4__lane3_strm1_data_valid    ( std__pe4__lane3_strm1_data_valid ),      
               .std__pe4__lane3_strm1_data_mask     ( std__pe4__lane3_strm1_data_mask  ),      

               // PE 4, Lane 4                 
               .pe4__std__lane4_strm0_ready         ( pe4__std__lane4_strm0_ready      ),      
               .std__pe4__lane4_strm0_cntl          ( std__pe4__lane4_strm0_cntl       ),      
               .std__pe4__lane4_strm0_data          ( std__pe4__lane4_strm0_data       ),      
               .std__pe4__lane4_strm0_data_valid    ( std__pe4__lane4_strm0_data_valid ),      
               .std__pe4__lane4_strm0_data_mask     ( std__pe4__lane4_strm0_data_mask  ),      

               .pe4__std__lane4_strm1_ready         ( pe4__std__lane4_strm1_ready      ),      
               .std__pe4__lane4_strm1_cntl          ( std__pe4__lane4_strm1_cntl       ),      
               .std__pe4__lane4_strm1_data          ( std__pe4__lane4_strm1_data       ),      
               .std__pe4__lane4_strm1_data_valid    ( std__pe4__lane4_strm1_data_valid ),      
               .std__pe4__lane4_strm1_data_mask     ( std__pe4__lane4_strm1_data_mask  ),      

               // PE 4, Lane 5                 
               .pe4__std__lane5_strm0_ready         ( pe4__std__lane5_strm0_ready      ),      
               .std__pe4__lane5_strm0_cntl          ( std__pe4__lane5_strm0_cntl       ),      
               .std__pe4__lane5_strm0_data          ( std__pe4__lane5_strm0_data       ),      
               .std__pe4__lane5_strm0_data_valid    ( std__pe4__lane5_strm0_data_valid ),      
               .std__pe4__lane5_strm0_data_mask     ( std__pe4__lane5_strm0_data_mask  ),      

               .pe4__std__lane5_strm1_ready         ( pe4__std__lane5_strm1_ready      ),      
               .std__pe4__lane5_strm1_cntl          ( std__pe4__lane5_strm1_cntl       ),      
               .std__pe4__lane5_strm1_data          ( std__pe4__lane5_strm1_data       ),      
               .std__pe4__lane5_strm1_data_valid    ( std__pe4__lane5_strm1_data_valid ),      
               .std__pe4__lane5_strm1_data_mask     ( std__pe4__lane5_strm1_data_mask  ),      

               // PE 4, Lane 6                 
               .pe4__std__lane6_strm0_ready         ( pe4__std__lane6_strm0_ready      ),      
               .std__pe4__lane6_strm0_cntl          ( std__pe4__lane6_strm0_cntl       ),      
               .std__pe4__lane6_strm0_data          ( std__pe4__lane6_strm0_data       ),      
               .std__pe4__lane6_strm0_data_valid    ( std__pe4__lane6_strm0_data_valid ),      
               .std__pe4__lane6_strm0_data_mask     ( std__pe4__lane6_strm0_data_mask  ),      

               .pe4__std__lane6_strm1_ready         ( pe4__std__lane6_strm1_ready      ),      
               .std__pe4__lane6_strm1_cntl          ( std__pe4__lane6_strm1_cntl       ),      
               .std__pe4__lane6_strm1_data          ( std__pe4__lane6_strm1_data       ),      
               .std__pe4__lane6_strm1_data_valid    ( std__pe4__lane6_strm1_data_valid ),      
               .std__pe4__lane6_strm1_data_mask     ( std__pe4__lane6_strm1_data_mask  ),      

               // PE 4, Lane 7                 
               .pe4__std__lane7_strm0_ready         ( pe4__std__lane7_strm0_ready      ),      
               .std__pe4__lane7_strm0_cntl          ( std__pe4__lane7_strm0_cntl       ),      
               .std__pe4__lane7_strm0_data          ( std__pe4__lane7_strm0_data       ),      
               .std__pe4__lane7_strm0_data_valid    ( std__pe4__lane7_strm0_data_valid ),      
               .std__pe4__lane7_strm0_data_mask     ( std__pe4__lane7_strm0_data_mask  ),      

               .pe4__std__lane7_strm1_ready         ( pe4__std__lane7_strm1_ready      ),      
               .std__pe4__lane7_strm1_cntl          ( std__pe4__lane7_strm1_cntl       ),      
               .std__pe4__lane7_strm1_data          ( std__pe4__lane7_strm1_data       ),      
               .std__pe4__lane7_strm1_data_valid    ( std__pe4__lane7_strm1_data_valid ),      
               .std__pe4__lane7_strm1_data_mask     ( std__pe4__lane7_strm1_data_mask  ),      

               // PE 4, Lane 8                 
               .pe4__std__lane8_strm0_ready         ( pe4__std__lane8_strm0_ready      ),      
               .std__pe4__lane8_strm0_cntl          ( std__pe4__lane8_strm0_cntl       ),      
               .std__pe4__lane8_strm0_data          ( std__pe4__lane8_strm0_data       ),      
               .std__pe4__lane8_strm0_data_valid    ( std__pe4__lane8_strm0_data_valid ),      
               .std__pe4__lane8_strm0_data_mask     ( std__pe4__lane8_strm0_data_mask  ),      

               .pe4__std__lane8_strm1_ready         ( pe4__std__lane8_strm1_ready      ),      
               .std__pe4__lane8_strm1_cntl          ( std__pe4__lane8_strm1_cntl       ),      
               .std__pe4__lane8_strm1_data          ( std__pe4__lane8_strm1_data       ),      
               .std__pe4__lane8_strm1_data_valid    ( std__pe4__lane8_strm1_data_valid ),      
               .std__pe4__lane8_strm1_data_mask     ( std__pe4__lane8_strm1_data_mask  ),      

               // PE 4, Lane 9                 
               .pe4__std__lane9_strm0_ready         ( pe4__std__lane9_strm0_ready      ),      
               .std__pe4__lane9_strm0_cntl          ( std__pe4__lane9_strm0_cntl       ),      
               .std__pe4__lane9_strm0_data          ( std__pe4__lane9_strm0_data       ),      
               .std__pe4__lane9_strm0_data_valid    ( std__pe4__lane9_strm0_data_valid ),      
               .std__pe4__lane9_strm0_data_mask     ( std__pe4__lane9_strm0_data_mask  ),      

               .pe4__std__lane9_strm1_ready         ( pe4__std__lane9_strm1_ready      ),      
               .std__pe4__lane9_strm1_cntl          ( std__pe4__lane9_strm1_cntl       ),      
               .std__pe4__lane9_strm1_data          ( std__pe4__lane9_strm1_data       ),      
               .std__pe4__lane9_strm1_data_valid    ( std__pe4__lane9_strm1_data_valid ),      
               .std__pe4__lane9_strm1_data_mask     ( std__pe4__lane9_strm1_data_mask  ),      

               // PE 4, Lane 10                 
               .pe4__std__lane10_strm0_ready         ( pe4__std__lane10_strm0_ready      ),      
               .std__pe4__lane10_strm0_cntl          ( std__pe4__lane10_strm0_cntl       ),      
               .std__pe4__lane10_strm0_data          ( std__pe4__lane10_strm0_data       ),      
               .std__pe4__lane10_strm0_data_valid    ( std__pe4__lane10_strm0_data_valid ),      
               .std__pe4__lane10_strm0_data_mask     ( std__pe4__lane10_strm0_data_mask  ),      

               .pe4__std__lane10_strm1_ready         ( pe4__std__lane10_strm1_ready      ),      
               .std__pe4__lane10_strm1_cntl          ( std__pe4__lane10_strm1_cntl       ),      
               .std__pe4__lane10_strm1_data          ( std__pe4__lane10_strm1_data       ),      
               .std__pe4__lane10_strm1_data_valid    ( std__pe4__lane10_strm1_data_valid ),      
               .std__pe4__lane10_strm1_data_mask     ( std__pe4__lane10_strm1_data_mask  ),      

               // PE 4, Lane 11                 
               .pe4__std__lane11_strm0_ready         ( pe4__std__lane11_strm0_ready      ),      
               .std__pe4__lane11_strm0_cntl          ( std__pe4__lane11_strm0_cntl       ),      
               .std__pe4__lane11_strm0_data          ( std__pe4__lane11_strm0_data       ),      
               .std__pe4__lane11_strm0_data_valid    ( std__pe4__lane11_strm0_data_valid ),      
               .std__pe4__lane11_strm0_data_mask     ( std__pe4__lane11_strm0_data_mask  ),      

               .pe4__std__lane11_strm1_ready         ( pe4__std__lane11_strm1_ready      ),      
               .std__pe4__lane11_strm1_cntl          ( std__pe4__lane11_strm1_cntl       ),      
               .std__pe4__lane11_strm1_data          ( std__pe4__lane11_strm1_data       ),      
               .std__pe4__lane11_strm1_data_valid    ( std__pe4__lane11_strm1_data_valid ),      
               .std__pe4__lane11_strm1_data_mask     ( std__pe4__lane11_strm1_data_mask  ),      

               // PE 4, Lane 12                 
               .pe4__std__lane12_strm0_ready         ( pe4__std__lane12_strm0_ready      ),      
               .std__pe4__lane12_strm0_cntl          ( std__pe4__lane12_strm0_cntl       ),      
               .std__pe4__lane12_strm0_data          ( std__pe4__lane12_strm0_data       ),      
               .std__pe4__lane12_strm0_data_valid    ( std__pe4__lane12_strm0_data_valid ),      
               .std__pe4__lane12_strm0_data_mask     ( std__pe4__lane12_strm0_data_mask  ),      

               .pe4__std__lane12_strm1_ready         ( pe4__std__lane12_strm1_ready      ),      
               .std__pe4__lane12_strm1_cntl          ( std__pe4__lane12_strm1_cntl       ),      
               .std__pe4__lane12_strm1_data          ( std__pe4__lane12_strm1_data       ),      
               .std__pe4__lane12_strm1_data_valid    ( std__pe4__lane12_strm1_data_valid ),      
               .std__pe4__lane12_strm1_data_mask     ( std__pe4__lane12_strm1_data_mask  ),      

               // PE 4, Lane 13                 
               .pe4__std__lane13_strm0_ready         ( pe4__std__lane13_strm0_ready      ),      
               .std__pe4__lane13_strm0_cntl          ( std__pe4__lane13_strm0_cntl       ),      
               .std__pe4__lane13_strm0_data          ( std__pe4__lane13_strm0_data       ),      
               .std__pe4__lane13_strm0_data_valid    ( std__pe4__lane13_strm0_data_valid ),      
               .std__pe4__lane13_strm0_data_mask     ( std__pe4__lane13_strm0_data_mask  ),      

               .pe4__std__lane13_strm1_ready         ( pe4__std__lane13_strm1_ready      ),      
               .std__pe4__lane13_strm1_cntl          ( std__pe4__lane13_strm1_cntl       ),      
               .std__pe4__lane13_strm1_data          ( std__pe4__lane13_strm1_data       ),      
               .std__pe4__lane13_strm1_data_valid    ( std__pe4__lane13_strm1_data_valid ),      
               .std__pe4__lane13_strm1_data_mask     ( std__pe4__lane13_strm1_data_mask  ),      

               // PE 4, Lane 14                 
               .pe4__std__lane14_strm0_ready         ( pe4__std__lane14_strm0_ready      ),      
               .std__pe4__lane14_strm0_cntl          ( std__pe4__lane14_strm0_cntl       ),      
               .std__pe4__lane14_strm0_data          ( std__pe4__lane14_strm0_data       ),      
               .std__pe4__lane14_strm0_data_valid    ( std__pe4__lane14_strm0_data_valid ),      
               .std__pe4__lane14_strm0_data_mask     ( std__pe4__lane14_strm0_data_mask  ),      

               .pe4__std__lane14_strm1_ready         ( pe4__std__lane14_strm1_ready      ),      
               .std__pe4__lane14_strm1_cntl          ( std__pe4__lane14_strm1_cntl       ),      
               .std__pe4__lane14_strm1_data          ( std__pe4__lane14_strm1_data       ),      
               .std__pe4__lane14_strm1_data_valid    ( std__pe4__lane14_strm1_data_valid ),      
               .std__pe4__lane14_strm1_data_mask     ( std__pe4__lane14_strm1_data_mask  ),      

               // PE 4, Lane 15                 
               .pe4__std__lane15_strm0_ready         ( pe4__std__lane15_strm0_ready      ),      
               .std__pe4__lane15_strm0_cntl          ( std__pe4__lane15_strm0_cntl       ),      
               .std__pe4__lane15_strm0_data          ( std__pe4__lane15_strm0_data       ),      
               .std__pe4__lane15_strm0_data_valid    ( std__pe4__lane15_strm0_data_valid ),      
               .std__pe4__lane15_strm0_data_mask     ( std__pe4__lane15_strm0_data_mask  ),      

               .pe4__std__lane15_strm1_ready         ( pe4__std__lane15_strm1_ready      ),      
               .std__pe4__lane15_strm1_cntl          ( std__pe4__lane15_strm1_cntl       ),      
               .std__pe4__lane15_strm1_data          ( std__pe4__lane15_strm1_data       ),      
               .std__pe4__lane15_strm1_data_valid    ( std__pe4__lane15_strm1_data_valid ),      
               .std__pe4__lane15_strm1_data_mask     ( std__pe4__lane15_strm1_data_mask  ),      

               // PE 4, Lane 16                 
               .pe4__std__lane16_strm0_ready         ( pe4__std__lane16_strm0_ready      ),      
               .std__pe4__lane16_strm0_cntl          ( std__pe4__lane16_strm0_cntl       ),      
               .std__pe4__lane16_strm0_data          ( std__pe4__lane16_strm0_data       ),      
               .std__pe4__lane16_strm0_data_valid    ( std__pe4__lane16_strm0_data_valid ),      
               .std__pe4__lane16_strm0_data_mask     ( std__pe4__lane16_strm0_data_mask  ),      

               .pe4__std__lane16_strm1_ready         ( pe4__std__lane16_strm1_ready      ),      
               .std__pe4__lane16_strm1_cntl          ( std__pe4__lane16_strm1_cntl       ),      
               .std__pe4__lane16_strm1_data          ( std__pe4__lane16_strm1_data       ),      
               .std__pe4__lane16_strm1_data_valid    ( std__pe4__lane16_strm1_data_valid ),      
               .std__pe4__lane16_strm1_data_mask     ( std__pe4__lane16_strm1_data_mask  ),      

               // PE 4, Lane 17                 
               .pe4__std__lane17_strm0_ready         ( pe4__std__lane17_strm0_ready      ),      
               .std__pe4__lane17_strm0_cntl          ( std__pe4__lane17_strm0_cntl       ),      
               .std__pe4__lane17_strm0_data          ( std__pe4__lane17_strm0_data       ),      
               .std__pe4__lane17_strm0_data_valid    ( std__pe4__lane17_strm0_data_valid ),      
               .std__pe4__lane17_strm0_data_mask     ( std__pe4__lane17_strm0_data_mask  ),      

               .pe4__std__lane17_strm1_ready         ( pe4__std__lane17_strm1_ready      ),      
               .std__pe4__lane17_strm1_cntl          ( std__pe4__lane17_strm1_cntl       ),      
               .std__pe4__lane17_strm1_data          ( std__pe4__lane17_strm1_data       ),      
               .std__pe4__lane17_strm1_data_valid    ( std__pe4__lane17_strm1_data_valid ),      
               .std__pe4__lane17_strm1_data_mask     ( std__pe4__lane17_strm1_data_mask  ),      

               // PE 4, Lane 18                 
               .pe4__std__lane18_strm0_ready         ( pe4__std__lane18_strm0_ready      ),      
               .std__pe4__lane18_strm0_cntl          ( std__pe4__lane18_strm0_cntl       ),      
               .std__pe4__lane18_strm0_data          ( std__pe4__lane18_strm0_data       ),      
               .std__pe4__lane18_strm0_data_valid    ( std__pe4__lane18_strm0_data_valid ),      
               .std__pe4__lane18_strm0_data_mask     ( std__pe4__lane18_strm0_data_mask  ),      

               .pe4__std__lane18_strm1_ready         ( pe4__std__lane18_strm1_ready      ),      
               .std__pe4__lane18_strm1_cntl          ( std__pe4__lane18_strm1_cntl       ),      
               .std__pe4__lane18_strm1_data          ( std__pe4__lane18_strm1_data       ),      
               .std__pe4__lane18_strm1_data_valid    ( std__pe4__lane18_strm1_data_valid ),      
               .std__pe4__lane18_strm1_data_mask     ( std__pe4__lane18_strm1_data_mask  ),      

               // PE 4, Lane 19                 
               .pe4__std__lane19_strm0_ready         ( pe4__std__lane19_strm0_ready      ),      
               .std__pe4__lane19_strm0_cntl          ( std__pe4__lane19_strm0_cntl       ),      
               .std__pe4__lane19_strm0_data          ( std__pe4__lane19_strm0_data       ),      
               .std__pe4__lane19_strm0_data_valid    ( std__pe4__lane19_strm0_data_valid ),      
               .std__pe4__lane19_strm0_data_mask     ( std__pe4__lane19_strm0_data_mask  ),      

               .pe4__std__lane19_strm1_ready         ( pe4__std__lane19_strm1_ready      ),      
               .std__pe4__lane19_strm1_cntl          ( std__pe4__lane19_strm1_cntl       ),      
               .std__pe4__lane19_strm1_data          ( std__pe4__lane19_strm1_data       ),      
               .std__pe4__lane19_strm1_data_valid    ( std__pe4__lane19_strm1_data_valid ),      
               .std__pe4__lane19_strm1_data_mask     ( std__pe4__lane19_strm1_data_mask  ),      

               // PE 4, Lane 20                 
               .pe4__std__lane20_strm0_ready         ( pe4__std__lane20_strm0_ready      ),      
               .std__pe4__lane20_strm0_cntl          ( std__pe4__lane20_strm0_cntl       ),      
               .std__pe4__lane20_strm0_data          ( std__pe4__lane20_strm0_data       ),      
               .std__pe4__lane20_strm0_data_valid    ( std__pe4__lane20_strm0_data_valid ),      
               .std__pe4__lane20_strm0_data_mask     ( std__pe4__lane20_strm0_data_mask  ),      

               .pe4__std__lane20_strm1_ready         ( pe4__std__lane20_strm1_ready      ),      
               .std__pe4__lane20_strm1_cntl          ( std__pe4__lane20_strm1_cntl       ),      
               .std__pe4__lane20_strm1_data          ( std__pe4__lane20_strm1_data       ),      
               .std__pe4__lane20_strm1_data_valid    ( std__pe4__lane20_strm1_data_valid ),      
               .std__pe4__lane20_strm1_data_mask     ( std__pe4__lane20_strm1_data_mask  ),      

               // PE 4, Lane 21                 
               .pe4__std__lane21_strm0_ready         ( pe4__std__lane21_strm0_ready      ),      
               .std__pe4__lane21_strm0_cntl          ( std__pe4__lane21_strm0_cntl       ),      
               .std__pe4__lane21_strm0_data          ( std__pe4__lane21_strm0_data       ),      
               .std__pe4__lane21_strm0_data_valid    ( std__pe4__lane21_strm0_data_valid ),      
               .std__pe4__lane21_strm0_data_mask     ( std__pe4__lane21_strm0_data_mask  ),      

               .pe4__std__lane21_strm1_ready         ( pe4__std__lane21_strm1_ready      ),      
               .std__pe4__lane21_strm1_cntl          ( std__pe4__lane21_strm1_cntl       ),      
               .std__pe4__lane21_strm1_data          ( std__pe4__lane21_strm1_data       ),      
               .std__pe4__lane21_strm1_data_valid    ( std__pe4__lane21_strm1_data_valid ),      
               .std__pe4__lane21_strm1_data_mask     ( std__pe4__lane21_strm1_data_mask  ),      

               // PE 4, Lane 22                 
               .pe4__std__lane22_strm0_ready         ( pe4__std__lane22_strm0_ready      ),      
               .std__pe4__lane22_strm0_cntl          ( std__pe4__lane22_strm0_cntl       ),      
               .std__pe4__lane22_strm0_data          ( std__pe4__lane22_strm0_data       ),      
               .std__pe4__lane22_strm0_data_valid    ( std__pe4__lane22_strm0_data_valid ),      
               .std__pe4__lane22_strm0_data_mask     ( std__pe4__lane22_strm0_data_mask  ),      

               .pe4__std__lane22_strm1_ready         ( pe4__std__lane22_strm1_ready      ),      
               .std__pe4__lane22_strm1_cntl          ( std__pe4__lane22_strm1_cntl       ),      
               .std__pe4__lane22_strm1_data          ( std__pe4__lane22_strm1_data       ),      
               .std__pe4__lane22_strm1_data_valid    ( std__pe4__lane22_strm1_data_valid ),      
               .std__pe4__lane22_strm1_data_mask     ( std__pe4__lane22_strm1_data_mask  ),      

               // PE 4, Lane 23                 
               .pe4__std__lane23_strm0_ready         ( pe4__std__lane23_strm0_ready      ),      
               .std__pe4__lane23_strm0_cntl          ( std__pe4__lane23_strm0_cntl       ),      
               .std__pe4__lane23_strm0_data          ( std__pe4__lane23_strm0_data       ),      
               .std__pe4__lane23_strm0_data_valid    ( std__pe4__lane23_strm0_data_valid ),      
               .std__pe4__lane23_strm0_data_mask     ( std__pe4__lane23_strm0_data_mask  ),      

               .pe4__std__lane23_strm1_ready         ( pe4__std__lane23_strm1_ready      ),      
               .std__pe4__lane23_strm1_cntl          ( std__pe4__lane23_strm1_cntl       ),      
               .std__pe4__lane23_strm1_data          ( std__pe4__lane23_strm1_data       ),      
               .std__pe4__lane23_strm1_data_valid    ( std__pe4__lane23_strm1_data_valid ),      
               .std__pe4__lane23_strm1_data_mask     ( std__pe4__lane23_strm1_data_mask  ),      

               // PE 4, Lane 24                 
               .pe4__std__lane24_strm0_ready         ( pe4__std__lane24_strm0_ready      ),      
               .std__pe4__lane24_strm0_cntl          ( std__pe4__lane24_strm0_cntl       ),      
               .std__pe4__lane24_strm0_data          ( std__pe4__lane24_strm0_data       ),      
               .std__pe4__lane24_strm0_data_valid    ( std__pe4__lane24_strm0_data_valid ),      
               .std__pe4__lane24_strm0_data_mask     ( std__pe4__lane24_strm0_data_mask  ),      

               .pe4__std__lane24_strm1_ready         ( pe4__std__lane24_strm1_ready      ),      
               .std__pe4__lane24_strm1_cntl          ( std__pe4__lane24_strm1_cntl       ),      
               .std__pe4__lane24_strm1_data          ( std__pe4__lane24_strm1_data       ),      
               .std__pe4__lane24_strm1_data_valid    ( std__pe4__lane24_strm1_data_valid ),      
               .std__pe4__lane24_strm1_data_mask     ( std__pe4__lane24_strm1_data_mask  ),      

               // PE 4, Lane 25                 
               .pe4__std__lane25_strm0_ready         ( pe4__std__lane25_strm0_ready      ),      
               .std__pe4__lane25_strm0_cntl          ( std__pe4__lane25_strm0_cntl       ),      
               .std__pe4__lane25_strm0_data          ( std__pe4__lane25_strm0_data       ),      
               .std__pe4__lane25_strm0_data_valid    ( std__pe4__lane25_strm0_data_valid ),      
               .std__pe4__lane25_strm0_data_mask     ( std__pe4__lane25_strm0_data_mask  ),      

               .pe4__std__lane25_strm1_ready         ( pe4__std__lane25_strm1_ready      ),      
               .std__pe4__lane25_strm1_cntl          ( std__pe4__lane25_strm1_cntl       ),      
               .std__pe4__lane25_strm1_data          ( std__pe4__lane25_strm1_data       ),      
               .std__pe4__lane25_strm1_data_valid    ( std__pe4__lane25_strm1_data_valid ),      
               .std__pe4__lane25_strm1_data_mask     ( std__pe4__lane25_strm1_data_mask  ),      

               // PE 4, Lane 26                 
               .pe4__std__lane26_strm0_ready         ( pe4__std__lane26_strm0_ready      ),      
               .std__pe4__lane26_strm0_cntl          ( std__pe4__lane26_strm0_cntl       ),      
               .std__pe4__lane26_strm0_data          ( std__pe4__lane26_strm0_data       ),      
               .std__pe4__lane26_strm0_data_valid    ( std__pe4__lane26_strm0_data_valid ),      
               .std__pe4__lane26_strm0_data_mask     ( std__pe4__lane26_strm0_data_mask  ),      

               .pe4__std__lane26_strm1_ready         ( pe4__std__lane26_strm1_ready      ),      
               .std__pe4__lane26_strm1_cntl          ( std__pe4__lane26_strm1_cntl       ),      
               .std__pe4__lane26_strm1_data          ( std__pe4__lane26_strm1_data       ),      
               .std__pe4__lane26_strm1_data_valid    ( std__pe4__lane26_strm1_data_valid ),      
               .std__pe4__lane26_strm1_data_mask     ( std__pe4__lane26_strm1_data_mask  ),      

               // PE 4, Lane 27                 
               .pe4__std__lane27_strm0_ready         ( pe4__std__lane27_strm0_ready      ),      
               .std__pe4__lane27_strm0_cntl          ( std__pe4__lane27_strm0_cntl       ),      
               .std__pe4__lane27_strm0_data          ( std__pe4__lane27_strm0_data       ),      
               .std__pe4__lane27_strm0_data_valid    ( std__pe4__lane27_strm0_data_valid ),      
               .std__pe4__lane27_strm0_data_mask     ( std__pe4__lane27_strm0_data_mask  ),      

               .pe4__std__lane27_strm1_ready         ( pe4__std__lane27_strm1_ready      ),      
               .std__pe4__lane27_strm1_cntl          ( std__pe4__lane27_strm1_cntl       ),      
               .std__pe4__lane27_strm1_data          ( std__pe4__lane27_strm1_data       ),      
               .std__pe4__lane27_strm1_data_valid    ( std__pe4__lane27_strm1_data_valid ),      
               .std__pe4__lane27_strm1_data_mask     ( std__pe4__lane27_strm1_data_mask  ),      

               // PE 4, Lane 28                 
               .pe4__std__lane28_strm0_ready         ( pe4__std__lane28_strm0_ready      ),      
               .std__pe4__lane28_strm0_cntl          ( std__pe4__lane28_strm0_cntl       ),      
               .std__pe4__lane28_strm0_data          ( std__pe4__lane28_strm0_data       ),      
               .std__pe4__lane28_strm0_data_valid    ( std__pe4__lane28_strm0_data_valid ),      
               .std__pe4__lane28_strm0_data_mask     ( std__pe4__lane28_strm0_data_mask  ),      

               .pe4__std__lane28_strm1_ready         ( pe4__std__lane28_strm1_ready      ),      
               .std__pe4__lane28_strm1_cntl          ( std__pe4__lane28_strm1_cntl       ),      
               .std__pe4__lane28_strm1_data          ( std__pe4__lane28_strm1_data       ),      
               .std__pe4__lane28_strm1_data_valid    ( std__pe4__lane28_strm1_data_valid ),      
               .std__pe4__lane28_strm1_data_mask     ( std__pe4__lane28_strm1_data_mask  ),      

               // PE 4, Lane 29                 
               .pe4__std__lane29_strm0_ready         ( pe4__std__lane29_strm0_ready      ),      
               .std__pe4__lane29_strm0_cntl          ( std__pe4__lane29_strm0_cntl       ),      
               .std__pe4__lane29_strm0_data          ( std__pe4__lane29_strm0_data       ),      
               .std__pe4__lane29_strm0_data_valid    ( std__pe4__lane29_strm0_data_valid ),      
               .std__pe4__lane29_strm0_data_mask     ( std__pe4__lane29_strm0_data_mask  ),      

               .pe4__std__lane29_strm1_ready         ( pe4__std__lane29_strm1_ready      ),      
               .std__pe4__lane29_strm1_cntl          ( std__pe4__lane29_strm1_cntl       ),      
               .std__pe4__lane29_strm1_data          ( std__pe4__lane29_strm1_data       ),      
               .std__pe4__lane29_strm1_data_valid    ( std__pe4__lane29_strm1_data_valid ),      
               .std__pe4__lane29_strm1_data_mask     ( std__pe4__lane29_strm1_data_mask  ),      

               // PE 4, Lane 30                 
               .pe4__std__lane30_strm0_ready         ( pe4__std__lane30_strm0_ready      ),      
               .std__pe4__lane30_strm0_cntl          ( std__pe4__lane30_strm0_cntl       ),      
               .std__pe4__lane30_strm0_data          ( std__pe4__lane30_strm0_data       ),      
               .std__pe4__lane30_strm0_data_valid    ( std__pe4__lane30_strm0_data_valid ),      
               .std__pe4__lane30_strm0_data_mask     ( std__pe4__lane30_strm0_data_mask  ),      

               .pe4__std__lane30_strm1_ready         ( pe4__std__lane30_strm1_ready      ),      
               .std__pe4__lane30_strm1_cntl          ( std__pe4__lane30_strm1_cntl       ),      
               .std__pe4__lane30_strm1_data          ( std__pe4__lane30_strm1_data       ),      
               .std__pe4__lane30_strm1_data_valid    ( std__pe4__lane30_strm1_data_valid ),      
               .std__pe4__lane30_strm1_data_mask     ( std__pe4__lane30_strm1_data_mask  ),      

               // PE 4, Lane 31                 
               .pe4__std__lane31_strm0_ready         ( pe4__std__lane31_strm0_ready      ),      
               .std__pe4__lane31_strm0_cntl          ( std__pe4__lane31_strm0_cntl       ),      
               .std__pe4__lane31_strm0_data          ( std__pe4__lane31_strm0_data       ),      
               .std__pe4__lane31_strm0_data_valid    ( std__pe4__lane31_strm0_data_valid ),      
               .std__pe4__lane31_strm0_data_mask     ( std__pe4__lane31_strm0_data_mask  ),      

               .pe4__std__lane31_strm1_ready         ( pe4__std__lane31_strm1_ready      ),      
               .std__pe4__lane31_strm1_cntl          ( std__pe4__lane31_strm1_cntl       ),      
               .std__pe4__lane31_strm1_data          ( std__pe4__lane31_strm1_data       ),      
               .std__pe4__lane31_strm1_data_valid    ( std__pe4__lane31_strm1_data_valid ),      
               .std__pe4__lane31_strm1_data_mask     ( std__pe4__lane31_strm1_data_mask  ),      

               // PE 5, Lane 0                 
               .pe5__std__lane0_strm0_ready         ( pe5__std__lane0_strm0_ready      ),      
               .std__pe5__lane0_strm0_cntl          ( std__pe5__lane0_strm0_cntl       ),      
               .std__pe5__lane0_strm0_data          ( std__pe5__lane0_strm0_data       ),      
               .std__pe5__lane0_strm0_data_valid    ( std__pe5__lane0_strm0_data_valid ),      
               .std__pe5__lane0_strm0_data_mask     ( std__pe5__lane0_strm0_data_mask  ),      

               .pe5__std__lane0_strm1_ready         ( pe5__std__lane0_strm1_ready      ),      
               .std__pe5__lane0_strm1_cntl          ( std__pe5__lane0_strm1_cntl       ),      
               .std__pe5__lane0_strm1_data          ( std__pe5__lane0_strm1_data       ),      
               .std__pe5__lane0_strm1_data_valid    ( std__pe5__lane0_strm1_data_valid ),      
               .std__pe5__lane0_strm1_data_mask     ( std__pe5__lane0_strm1_data_mask  ),      

               // PE 5, Lane 1                 
               .pe5__std__lane1_strm0_ready         ( pe5__std__lane1_strm0_ready      ),      
               .std__pe5__lane1_strm0_cntl          ( std__pe5__lane1_strm0_cntl       ),      
               .std__pe5__lane1_strm0_data          ( std__pe5__lane1_strm0_data       ),      
               .std__pe5__lane1_strm0_data_valid    ( std__pe5__lane1_strm0_data_valid ),      
               .std__pe5__lane1_strm0_data_mask     ( std__pe5__lane1_strm0_data_mask  ),      

               .pe5__std__lane1_strm1_ready         ( pe5__std__lane1_strm1_ready      ),      
               .std__pe5__lane1_strm1_cntl          ( std__pe5__lane1_strm1_cntl       ),      
               .std__pe5__lane1_strm1_data          ( std__pe5__lane1_strm1_data       ),      
               .std__pe5__lane1_strm1_data_valid    ( std__pe5__lane1_strm1_data_valid ),      
               .std__pe5__lane1_strm1_data_mask     ( std__pe5__lane1_strm1_data_mask  ),      

               // PE 5, Lane 2                 
               .pe5__std__lane2_strm0_ready         ( pe5__std__lane2_strm0_ready      ),      
               .std__pe5__lane2_strm0_cntl          ( std__pe5__lane2_strm0_cntl       ),      
               .std__pe5__lane2_strm0_data          ( std__pe5__lane2_strm0_data       ),      
               .std__pe5__lane2_strm0_data_valid    ( std__pe5__lane2_strm0_data_valid ),      
               .std__pe5__lane2_strm0_data_mask     ( std__pe5__lane2_strm0_data_mask  ),      

               .pe5__std__lane2_strm1_ready         ( pe5__std__lane2_strm1_ready      ),      
               .std__pe5__lane2_strm1_cntl          ( std__pe5__lane2_strm1_cntl       ),      
               .std__pe5__lane2_strm1_data          ( std__pe5__lane2_strm1_data       ),      
               .std__pe5__lane2_strm1_data_valid    ( std__pe5__lane2_strm1_data_valid ),      
               .std__pe5__lane2_strm1_data_mask     ( std__pe5__lane2_strm1_data_mask  ),      

               // PE 5, Lane 3                 
               .pe5__std__lane3_strm0_ready         ( pe5__std__lane3_strm0_ready      ),      
               .std__pe5__lane3_strm0_cntl          ( std__pe5__lane3_strm0_cntl       ),      
               .std__pe5__lane3_strm0_data          ( std__pe5__lane3_strm0_data       ),      
               .std__pe5__lane3_strm0_data_valid    ( std__pe5__lane3_strm0_data_valid ),      
               .std__pe5__lane3_strm0_data_mask     ( std__pe5__lane3_strm0_data_mask  ),      

               .pe5__std__lane3_strm1_ready         ( pe5__std__lane3_strm1_ready      ),      
               .std__pe5__lane3_strm1_cntl          ( std__pe5__lane3_strm1_cntl       ),      
               .std__pe5__lane3_strm1_data          ( std__pe5__lane3_strm1_data       ),      
               .std__pe5__lane3_strm1_data_valid    ( std__pe5__lane3_strm1_data_valid ),      
               .std__pe5__lane3_strm1_data_mask     ( std__pe5__lane3_strm1_data_mask  ),      

               // PE 5, Lane 4                 
               .pe5__std__lane4_strm0_ready         ( pe5__std__lane4_strm0_ready      ),      
               .std__pe5__lane4_strm0_cntl          ( std__pe5__lane4_strm0_cntl       ),      
               .std__pe5__lane4_strm0_data          ( std__pe5__lane4_strm0_data       ),      
               .std__pe5__lane4_strm0_data_valid    ( std__pe5__lane4_strm0_data_valid ),      
               .std__pe5__lane4_strm0_data_mask     ( std__pe5__lane4_strm0_data_mask  ),      

               .pe5__std__lane4_strm1_ready         ( pe5__std__lane4_strm1_ready      ),      
               .std__pe5__lane4_strm1_cntl          ( std__pe5__lane4_strm1_cntl       ),      
               .std__pe5__lane4_strm1_data          ( std__pe5__lane4_strm1_data       ),      
               .std__pe5__lane4_strm1_data_valid    ( std__pe5__lane4_strm1_data_valid ),      
               .std__pe5__lane4_strm1_data_mask     ( std__pe5__lane4_strm1_data_mask  ),      

               // PE 5, Lane 5                 
               .pe5__std__lane5_strm0_ready         ( pe5__std__lane5_strm0_ready      ),      
               .std__pe5__lane5_strm0_cntl          ( std__pe5__lane5_strm0_cntl       ),      
               .std__pe5__lane5_strm0_data          ( std__pe5__lane5_strm0_data       ),      
               .std__pe5__lane5_strm0_data_valid    ( std__pe5__lane5_strm0_data_valid ),      
               .std__pe5__lane5_strm0_data_mask     ( std__pe5__lane5_strm0_data_mask  ),      

               .pe5__std__lane5_strm1_ready         ( pe5__std__lane5_strm1_ready      ),      
               .std__pe5__lane5_strm1_cntl          ( std__pe5__lane5_strm1_cntl       ),      
               .std__pe5__lane5_strm1_data          ( std__pe5__lane5_strm1_data       ),      
               .std__pe5__lane5_strm1_data_valid    ( std__pe5__lane5_strm1_data_valid ),      
               .std__pe5__lane5_strm1_data_mask     ( std__pe5__lane5_strm1_data_mask  ),      

               // PE 5, Lane 6                 
               .pe5__std__lane6_strm0_ready         ( pe5__std__lane6_strm0_ready      ),      
               .std__pe5__lane6_strm0_cntl          ( std__pe5__lane6_strm0_cntl       ),      
               .std__pe5__lane6_strm0_data          ( std__pe5__lane6_strm0_data       ),      
               .std__pe5__lane6_strm0_data_valid    ( std__pe5__lane6_strm0_data_valid ),      
               .std__pe5__lane6_strm0_data_mask     ( std__pe5__lane6_strm0_data_mask  ),      

               .pe5__std__lane6_strm1_ready         ( pe5__std__lane6_strm1_ready      ),      
               .std__pe5__lane6_strm1_cntl          ( std__pe5__lane6_strm1_cntl       ),      
               .std__pe5__lane6_strm1_data          ( std__pe5__lane6_strm1_data       ),      
               .std__pe5__lane6_strm1_data_valid    ( std__pe5__lane6_strm1_data_valid ),      
               .std__pe5__lane6_strm1_data_mask     ( std__pe5__lane6_strm1_data_mask  ),      

               // PE 5, Lane 7                 
               .pe5__std__lane7_strm0_ready         ( pe5__std__lane7_strm0_ready      ),      
               .std__pe5__lane7_strm0_cntl          ( std__pe5__lane7_strm0_cntl       ),      
               .std__pe5__lane7_strm0_data          ( std__pe5__lane7_strm0_data       ),      
               .std__pe5__lane7_strm0_data_valid    ( std__pe5__lane7_strm0_data_valid ),      
               .std__pe5__lane7_strm0_data_mask     ( std__pe5__lane7_strm0_data_mask  ),      

               .pe5__std__lane7_strm1_ready         ( pe5__std__lane7_strm1_ready      ),      
               .std__pe5__lane7_strm1_cntl          ( std__pe5__lane7_strm1_cntl       ),      
               .std__pe5__lane7_strm1_data          ( std__pe5__lane7_strm1_data       ),      
               .std__pe5__lane7_strm1_data_valid    ( std__pe5__lane7_strm1_data_valid ),      
               .std__pe5__lane7_strm1_data_mask     ( std__pe5__lane7_strm1_data_mask  ),      

               // PE 5, Lane 8                 
               .pe5__std__lane8_strm0_ready         ( pe5__std__lane8_strm0_ready      ),      
               .std__pe5__lane8_strm0_cntl          ( std__pe5__lane8_strm0_cntl       ),      
               .std__pe5__lane8_strm0_data          ( std__pe5__lane8_strm0_data       ),      
               .std__pe5__lane8_strm0_data_valid    ( std__pe5__lane8_strm0_data_valid ),      
               .std__pe5__lane8_strm0_data_mask     ( std__pe5__lane8_strm0_data_mask  ),      

               .pe5__std__lane8_strm1_ready         ( pe5__std__lane8_strm1_ready      ),      
               .std__pe5__lane8_strm1_cntl          ( std__pe5__lane8_strm1_cntl       ),      
               .std__pe5__lane8_strm1_data          ( std__pe5__lane8_strm1_data       ),      
               .std__pe5__lane8_strm1_data_valid    ( std__pe5__lane8_strm1_data_valid ),      
               .std__pe5__lane8_strm1_data_mask     ( std__pe5__lane8_strm1_data_mask  ),      

               // PE 5, Lane 9                 
               .pe5__std__lane9_strm0_ready         ( pe5__std__lane9_strm0_ready      ),      
               .std__pe5__lane9_strm0_cntl          ( std__pe5__lane9_strm0_cntl       ),      
               .std__pe5__lane9_strm0_data          ( std__pe5__lane9_strm0_data       ),      
               .std__pe5__lane9_strm0_data_valid    ( std__pe5__lane9_strm0_data_valid ),      
               .std__pe5__lane9_strm0_data_mask     ( std__pe5__lane9_strm0_data_mask  ),      

               .pe5__std__lane9_strm1_ready         ( pe5__std__lane9_strm1_ready      ),      
               .std__pe5__lane9_strm1_cntl          ( std__pe5__lane9_strm1_cntl       ),      
               .std__pe5__lane9_strm1_data          ( std__pe5__lane9_strm1_data       ),      
               .std__pe5__lane9_strm1_data_valid    ( std__pe5__lane9_strm1_data_valid ),      
               .std__pe5__lane9_strm1_data_mask     ( std__pe5__lane9_strm1_data_mask  ),      

               // PE 5, Lane 10                 
               .pe5__std__lane10_strm0_ready         ( pe5__std__lane10_strm0_ready      ),      
               .std__pe5__lane10_strm0_cntl          ( std__pe5__lane10_strm0_cntl       ),      
               .std__pe5__lane10_strm0_data          ( std__pe5__lane10_strm0_data       ),      
               .std__pe5__lane10_strm0_data_valid    ( std__pe5__lane10_strm0_data_valid ),      
               .std__pe5__lane10_strm0_data_mask     ( std__pe5__lane10_strm0_data_mask  ),      

               .pe5__std__lane10_strm1_ready         ( pe5__std__lane10_strm1_ready      ),      
               .std__pe5__lane10_strm1_cntl          ( std__pe5__lane10_strm1_cntl       ),      
               .std__pe5__lane10_strm1_data          ( std__pe5__lane10_strm1_data       ),      
               .std__pe5__lane10_strm1_data_valid    ( std__pe5__lane10_strm1_data_valid ),      
               .std__pe5__lane10_strm1_data_mask     ( std__pe5__lane10_strm1_data_mask  ),      

               // PE 5, Lane 11                 
               .pe5__std__lane11_strm0_ready         ( pe5__std__lane11_strm0_ready      ),      
               .std__pe5__lane11_strm0_cntl          ( std__pe5__lane11_strm0_cntl       ),      
               .std__pe5__lane11_strm0_data          ( std__pe5__lane11_strm0_data       ),      
               .std__pe5__lane11_strm0_data_valid    ( std__pe5__lane11_strm0_data_valid ),      
               .std__pe5__lane11_strm0_data_mask     ( std__pe5__lane11_strm0_data_mask  ),      

               .pe5__std__lane11_strm1_ready         ( pe5__std__lane11_strm1_ready      ),      
               .std__pe5__lane11_strm1_cntl          ( std__pe5__lane11_strm1_cntl       ),      
               .std__pe5__lane11_strm1_data          ( std__pe5__lane11_strm1_data       ),      
               .std__pe5__lane11_strm1_data_valid    ( std__pe5__lane11_strm1_data_valid ),      
               .std__pe5__lane11_strm1_data_mask     ( std__pe5__lane11_strm1_data_mask  ),      

               // PE 5, Lane 12                 
               .pe5__std__lane12_strm0_ready         ( pe5__std__lane12_strm0_ready      ),      
               .std__pe5__lane12_strm0_cntl          ( std__pe5__lane12_strm0_cntl       ),      
               .std__pe5__lane12_strm0_data          ( std__pe5__lane12_strm0_data       ),      
               .std__pe5__lane12_strm0_data_valid    ( std__pe5__lane12_strm0_data_valid ),      
               .std__pe5__lane12_strm0_data_mask     ( std__pe5__lane12_strm0_data_mask  ),      

               .pe5__std__lane12_strm1_ready         ( pe5__std__lane12_strm1_ready      ),      
               .std__pe5__lane12_strm1_cntl          ( std__pe5__lane12_strm1_cntl       ),      
               .std__pe5__lane12_strm1_data          ( std__pe5__lane12_strm1_data       ),      
               .std__pe5__lane12_strm1_data_valid    ( std__pe5__lane12_strm1_data_valid ),      
               .std__pe5__lane12_strm1_data_mask     ( std__pe5__lane12_strm1_data_mask  ),      

               // PE 5, Lane 13                 
               .pe5__std__lane13_strm0_ready         ( pe5__std__lane13_strm0_ready      ),      
               .std__pe5__lane13_strm0_cntl          ( std__pe5__lane13_strm0_cntl       ),      
               .std__pe5__lane13_strm0_data          ( std__pe5__lane13_strm0_data       ),      
               .std__pe5__lane13_strm0_data_valid    ( std__pe5__lane13_strm0_data_valid ),      
               .std__pe5__lane13_strm0_data_mask     ( std__pe5__lane13_strm0_data_mask  ),      

               .pe5__std__lane13_strm1_ready         ( pe5__std__lane13_strm1_ready      ),      
               .std__pe5__lane13_strm1_cntl          ( std__pe5__lane13_strm1_cntl       ),      
               .std__pe5__lane13_strm1_data          ( std__pe5__lane13_strm1_data       ),      
               .std__pe5__lane13_strm1_data_valid    ( std__pe5__lane13_strm1_data_valid ),      
               .std__pe5__lane13_strm1_data_mask     ( std__pe5__lane13_strm1_data_mask  ),      

               // PE 5, Lane 14                 
               .pe5__std__lane14_strm0_ready         ( pe5__std__lane14_strm0_ready      ),      
               .std__pe5__lane14_strm0_cntl          ( std__pe5__lane14_strm0_cntl       ),      
               .std__pe5__lane14_strm0_data          ( std__pe5__lane14_strm0_data       ),      
               .std__pe5__lane14_strm0_data_valid    ( std__pe5__lane14_strm0_data_valid ),      
               .std__pe5__lane14_strm0_data_mask     ( std__pe5__lane14_strm0_data_mask  ),      

               .pe5__std__lane14_strm1_ready         ( pe5__std__lane14_strm1_ready      ),      
               .std__pe5__lane14_strm1_cntl          ( std__pe5__lane14_strm1_cntl       ),      
               .std__pe5__lane14_strm1_data          ( std__pe5__lane14_strm1_data       ),      
               .std__pe5__lane14_strm1_data_valid    ( std__pe5__lane14_strm1_data_valid ),      
               .std__pe5__lane14_strm1_data_mask     ( std__pe5__lane14_strm1_data_mask  ),      

               // PE 5, Lane 15                 
               .pe5__std__lane15_strm0_ready         ( pe5__std__lane15_strm0_ready      ),      
               .std__pe5__lane15_strm0_cntl          ( std__pe5__lane15_strm0_cntl       ),      
               .std__pe5__lane15_strm0_data          ( std__pe5__lane15_strm0_data       ),      
               .std__pe5__lane15_strm0_data_valid    ( std__pe5__lane15_strm0_data_valid ),      
               .std__pe5__lane15_strm0_data_mask     ( std__pe5__lane15_strm0_data_mask  ),      

               .pe5__std__lane15_strm1_ready         ( pe5__std__lane15_strm1_ready      ),      
               .std__pe5__lane15_strm1_cntl          ( std__pe5__lane15_strm1_cntl       ),      
               .std__pe5__lane15_strm1_data          ( std__pe5__lane15_strm1_data       ),      
               .std__pe5__lane15_strm1_data_valid    ( std__pe5__lane15_strm1_data_valid ),      
               .std__pe5__lane15_strm1_data_mask     ( std__pe5__lane15_strm1_data_mask  ),      

               // PE 5, Lane 16                 
               .pe5__std__lane16_strm0_ready         ( pe5__std__lane16_strm0_ready      ),      
               .std__pe5__lane16_strm0_cntl          ( std__pe5__lane16_strm0_cntl       ),      
               .std__pe5__lane16_strm0_data          ( std__pe5__lane16_strm0_data       ),      
               .std__pe5__lane16_strm0_data_valid    ( std__pe5__lane16_strm0_data_valid ),      
               .std__pe5__lane16_strm0_data_mask     ( std__pe5__lane16_strm0_data_mask  ),      

               .pe5__std__lane16_strm1_ready         ( pe5__std__lane16_strm1_ready      ),      
               .std__pe5__lane16_strm1_cntl          ( std__pe5__lane16_strm1_cntl       ),      
               .std__pe5__lane16_strm1_data          ( std__pe5__lane16_strm1_data       ),      
               .std__pe5__lane16_strm1_data_valid    ( std__pe5__lane16_strm1_data_valid ),      
               .std__pe5__lane16_strm1_data_mask     ( std__pe5__lane16_strm1_data_mask  ),      

               // PE 5, Lane 17                 
               .pe5__std__lane17_strm0_ready         ( pe5__std__lane17_strm0_ready      ),      
               .std__pe5__lane17_strm0_cntl          ( std__pe5__lane17_strm0_cntl       ),      
               .std__pe5__lane17_strm0_data          ( std__pe5__lane17_strm0_data       ),      
               .std__pe5__lane17_strm0_data_valid    ( std__pe5__lane17_strm0_data_valid ),      
               .std__pe5__lane17_strm0_data_mask     ( std__pe5__lane17_strm0_data_mask  ),      

               .pe5__std__lane17_strm1_ready         ( pe5__std__lane17_strm1_ready      ),      
               .std__pe5__lane17_strm1_cntl          ( std__pe5__lane17_strm1_cntl       ),      
               .std__pe5__lane17_strm1_data          ( std__pe5__lane17_strm1_data       ),      
               .std__pe5__lane17_strm1_data_valid    ( std__pe5__lane17_strm1_data_valid ),      
               .std__pe5__lane17_strm1_data_mask     ( std__pe5__lane17_strm1_data_mask  ),      

               // PE 5, Lane 18                 
               .pe5__std__lane18_strm0_ready         ( pe5__std__lane18_strm0_ready      ),      
               .std__pe5__lane18_strm0_cntl          ( std__pe5__lane18_strm0_cntl       ),      
               .std__pe5__lane18_strm0_data          ( std__pe5__lane18_strm0_data       ),      
               .std__pe5__lane18_strm0_data_valid    ( std__pe5__lane18_strm0_data_valid ),      
               .std__pe5__lane18_strm0_data_mask     ( std__pe5__lane18_strm0_data_mask  ),      

               .pe5__std__lane18_strm1_ready         ( pe5__std__lane18_strm1_ready      ),      
               .std__pe5__lane18_strm1_cntl          ( std__pe5__lane18_strm1_cntl       ),      
               .std__pe5__lane18_strm1_data          ( std__pe5__lane18_strm1_data       ),      
               .std__pe5__lane18_strm1_data_valid    ( std__pe5__lane18_strm1_data_valid ),      
               .std__pe5__lane18_strm1_data_mask     ( std__pe5__lane18_strm1_data_mask  ),      

               // PE 5, Lane 19                 
               .pe5__std__lane19_strm0_ready         ( pe5__std__lane19_strm0_ready      ),      
               .std__pe5__lane19_strm0_cntl          ( std__pe5__lane19_strm0_cntl       ),      
               .std__pe5__lane19_strm0_data          ( std__pe5__lane19_strm0_data       ),      
               .std__pe5__lane19_strm0_data_valid    ( std__pe5__lane19_strm0_data_valid ),      
               .std__pe5__lane19_strm0_data_mask     ( std__pe5__lane19_strm0_data_mask  ),      

               .pe5__std__lane19_strm1_ready         ( pe5__std__lane19_strm1_ready      ),      
               .std__pe5__lane19_strm1_cntl          ( std__pe5__lane19_strm1_cntl       ),      
               .std__pe5__lane19_strm1_data          ( std__pe5__lane19_strm1_data       ),      
               .std__pe5__lane19_strm1_data_valid    ( std__pe5__lane19_strm1_data_valid ),      
               .std__pe5__lane19_strm1_data_mask     ( std__pe5__lane19_strm1_data_mask  ),      

               // PE 5, Lane 20                 
               .pe5__std__lane20_strm0_ready         ( pe5__std__lane20_strm0_ready      ),      
               .std__pe5__lane20_strm0_cntl          ( std__pe5__lane20_strm0_cntl       ),      
               .std__pe5__lane20_strm0_data          ( std__pe5__lane20_strm0_data       ),      
               .std__pe5__lane20_strm0_data_valid    ( std__pe5__lane20_strm0_data_valid ),      
               .std__pe5__lane20_strm0_data_mask     ( std__pe5__lane20_strm0_data_mask  ),      

               .pe5__std__lane20_strm1_ready         ( pe5__std__lane20_strm1_ready      ),      
               .std__pe5__lane20_strm1_cntl          ( std__pe5__lane20_strm1_cntl       ),      
               .std__pe5__lane20_strm1_data          ( std__pe5__lane20_strm1_data       ),      
               .std__pe5__lane20_strm1_data_valid    ( std__pe5__lane20_strm1_data_valid ),      
               .std__pe5__lane20_strm1_data_mask     ( std__pe5__lane20_strm1_data_mask  ),      

               // PE 5, Lane 21                 
               .pe5__std__lane21_strm0_ready         ( pe5__std__lane21_strm0_ready      ),      
               .std__pe5__lane21_strm0_cntl          ( std__pe5__lane21_strm0_cntl       ),      
               .std__pe5__lane21_strm0_data          ( std__pe5__lane21_strm0_data       ),      
               .std__pe5__lane21_strm0_data_valid    ( std__pe5__lane21_strm0_data_valid ),      
               .std__pe5__lane21_strm0_data_mask     ( std__pe5__lane21_strm0_data_mask  ),      

               .pe5__std__lane21_strm1_ready         ( pe5__std__lane21_strm1_ready      ),      
               .std__pe5__lane21_strm1_cntl          ( std__pe5__lane21_strm1_cntl       ),      
               .std__pe5__lane21_strm1_data          ( std__pe5__lane21_strm1_data       ),      
               .std__pe5__lane21_strm1_data_valid    ( std__pe5__lane21_strm1_data_valid ),      
               .std__pe5__lane21_strm1_data_mask     ( std__pe5__lane21_strm1_data_mask  ),      

               // PE 5, Lane 22                 
               .pe5__std__lane22_strm0_ready         ( pe5__std__lane22_strm0_ready      ),      
               .std__pe5__lane22_strm0_cntl          ( std__pe5__lane22_strm0_cntl       ),      
               .std__pe5__lane22_strm0_data          ( std__pe5__lane22_strm0_data       ),      
               .std__pe5__lane22_strm0_data_valid    ( std__pe5__lane22_strm0_data_valid ),      
               .std__pe5__lane22_strm0_data_mask     ( std__pe5__lane22_strm0_data_mask  ),      

               .pe5__std__lane22_strm1_ready         ( pe5__std__lane22_strm1_ready      ),      
               .std__pe5__lane22_strm1_cntl          ( std__pe5__lane22_strm1_cntl       ),      
               .std__pe5__lane22_strm1_data          ( std__pe5__lane22_strm1_data       ),      
               .std__pe5__lane22_strm1_data_valid    ( std__pe5__lane22_strm1_data_valid ),      
               .std__pe5__lane22_strm1_data_mask     ( std__pe5__lane22_strm1_data_mask  ),      

               // PE 5, Lane 23                 
               .pe5__std__lane23_strm0_ready         ( pe5__std__lane23_strm0_ready      ),      
               .std__pe5__lane23_strm0_cntl          ( std__pe5__lane23_strm0_cntl       ),      
               .std__pe5__lane23_strm0_data          ( std__pe5__lane23_strm0_data       ),      
               .std__pe5__lane23_strm0_data_valid    ( std__pe5__lane23_strm0_data_valid ),      
               .std__pe5__lane23_strm0_data_mask     ( std__pe5__lane23_strm0_data_mask  ),      

               .pe5__std__lane23_strm1_ready         ( pe5__std__lane23_strm1_ready      ),      
               .std__pe5__lane23_strm1_cntl          ( std__pe5__lane23_strm1_cntl       ),      
               .std__pe5__lane23_strm1_data          ( std__pe5__lane23_strm1_data       ),      
               .std__pe5__lane23_strm1_data_valid    ( std__pe5__lane23_strm1_data_valid ),      
               .std__pe5__lane23_strm1_data_mask     ( std__pe5__lane23_strm1_data_mask  ),      

               // PE 5, Lane 24                 
               .pe5__std__lane24_strm0_ready         ( pe5__std__lane24_strm0_ready      ),      
               .std__pe5__lane24_strm0_cntl          ( std__pe5__lane24_strm0_cntl       ),      
               .std__pe5__lane24_strm0_data          ( std__pe5__lane24_strm0_data       ),      
               .std__pe5__lane24_strm0_data_valid    ( std__pe5__lane24_strm0_data_valid ),      
               .std__pe5__lane24_strm0_data_mask     ( std__pe5__lane24_strm0_data_mask  ),      

               .pe5__std__lane24_strm1_ready         ( pe5__std__lane24_strm1_ready      ),      
               .std__pe5__lane24_strm1_cntl          ( std__pe5__lane24_strm1_cntl       ),      
               .std__pe5__lane24_strm1_data          ( std__pe5__lane24_strm1_data       ),      
               .std__pe5__lane24_strm1_data_valid    ( std__pe5__lane24_strm1_data_valid ),      
               .std__pe5__lane24_strm1_data_mask     ( std__pe5__lane24_strm1_data_mask  ),      

               // PE 5, Lane 25                 
               .pe5__std__lane25_strm0_ready         ( pe5__std__lane25_strm0_ready      ),      
               .std__pe5__lane25_strm0_cntl          ( std__pe5__lane25_strm0_cntl       ),      
               .std__pe5__lane25_strm0_data          ( std__pe5__lane25_strm0_data       ),      
               .std__pe5__lane25_strm0_data_valid    ( std__pe5__lane25_strm0_data_valid ),      
               .std__pe5__lane25_strm0_data_mask     ( std__pe5__lane25_strm0_data_mask  ),      

               .pe5__std__lane25_strm1_ready         ( pe5__std__lane25_strm1_ready      ),      
               .std__pe5__lane25_strm1_cntl          ( std__pe5__lane25_strm1_cntl       ),      
               .std__pe5__lane25_strm1_data          ( std__pe5__lane25_strm1_data       ),      
               .std__pe5__lane25_strm1_data_valid    ( std__pe5__lane25_strm1_data_valid ),      
               .std__pe5__lane25_strm1_data_mask     ( std__pe5__lane25_strm1_data_mask  ),      

               // PE 5, Lane 26                 
               .pe5__std__lane26_strm0_ready         ( pe5__std__lane26_strm0_ready      ),      
               .std__pe5__lane26_strm0_cntl          ( std__pe5__lane26_strm0_cntl       ),      
               .std__pe5__lane26_strm0_data          ( std__pe5__lane26_strm0_data       ),      
               .std__pe5__lane26_strm0_data_valid    ( std__pe5__lane26_strm0_data_valid ),      
               .std__pe5__lane26_strm0_data_mask     ( std__pe5__lane26_strm0_data_mask  ),      

               .pe5__std__lane26_strm1_ready         ( pe5__std__lane26_strm1_ready      ),      
               .std__pe5__lane26_strm1_cntl          ( std__pe5__lane26_strm1_cntl       ),      
               .std__pe5__lane26_strm1_data          ( std__pe5__lane26_strm1_data       ),      
               .std__pe5__lane26_strm1_data_valid    ( std__pe5__lane26_strm1_data_valid ),      
               .std__pe5__lane26_strm1_data_mask     ( std__pe5__lane26_strm1_data_mask  ),      

               // PE 5, Lane 27                 
               .pe5__std__lane27_strm0_ready         ( pe5__std__lane27_strm0_ready      ),      
               .std__pe5__lane27_strm0_cntl          ( std__pe5__lane27_strm0_cntl       ),      
               .std__pe5__lane27_strm0_data          ( std__pe5__lane27_strm0_data       ),      
               .std__pe5__lane27_strm0_data_valid    ( std__pe5__lane27_strm0_data_valid ),      
               .std__pe5__lane27_strm0_data_mask     ( std__pe5__lane27_strm0_data_mask  ),      

               .pe5__std__lane27_strm1_ready         ( pe5__std__lane27_strm1_ready      ),      
               .std__pe5__lane27_strm1_cntl          ( std__pe5__lane27_strm1_cntl       ),      
               .std__pe5__lane27_strm1_data          ( std__pe5__lane27_strm1_data       ),      
               .std__pe5__lane27_strm1_data_valid    ( std__pe5__lane27_strm1_data_valid ),      
               .std__pe5__lane27_strm1_data_mask     ( std__pe5__lane27_strm1_data_mask  ),      

               // PE 5, Lane 28                 
               .pe5__std__lane28_strm0_ready         ( pe5__std__lane28_strm0_ready      ),      
               .std__pe5__lane28_strm0_cntl          ( std__pe5__lane28_strm0_cntl       ),      
               .std__pe5__lane28_strm0_data          ( std__pe5__lane28_strm0_data       ),      
               .std__pe5__lane28_strm0_data_valid    ( std__pe5__lane28_strm0_data_valid ),      
               .std__pe5__lane28_strm0_data_mask     ( std__pe5__lane28_strm0_data_mask  ),      

               .pe5__std__lane28_strm1_ready         ( pe5__std__lane28_strm1_ready      ),      
               .std__pe5__lane28_strm1_cntl          ( std__pe5__lane28_strm1_cntl       ),      
               .std__pe5__lane28_strm1_data          ( std__pe5__lane28_strm1_data       ),      
               .std__pe5__lane28_strm1_data_valid    ( std__pe5__lane28_strm1_data_valid ),      
               .std__pe5__lane28_strm1_data_mask     ( std__pe5__lane28_strm1_data_mask  ),      

               // PE 5, Lane 29                 
               .pe5__std__lane29_strm0_ready         ( pe5__std__lane29_strm0_ready      ),      
               .std__pe5__lane29_strm0_cntl          ( std__pe5__lane29_strm0_cntl       ),      
               .std__pe5__lane29_strm0_data          ( std__pe5__lane29_strm0_data       ),      
               .std__pe5__lane29_strm0_data_valid    ( std__pe5__lane29_strm0_data_valid ),      
               .std__pe5__lane29_strm0_data_mask     ( std__pe5__lane29_strm0_data_mask  ),      

               .pe5__std__lane29_strm1_ready         ( pe5__std__lane29_strm1_ready      ),      
               .std__pe5__lane29_strm1_cntl          ( std__pe5__lane29_strm1_cntl       ),      
               .std__pe5__lane29_strm1_data          ( std__pe5__lane29_strm1_data       ),      
               .std__pe5__lane29_strm1_data_valid    ( std__pe5__lane29_strm1_data_valid ),      
               .std__pe5__lane29_strm1_data_mask     ( std__pe5__lane29_strm1_data_mask  ),      

               // PE 5, Lane 30                 
               .pe5__std__lane30_strm0_ready         ( pe5__std__lane30_strm0_ready      ),      
               .std__pe5__lane30_strm0_cntl          ( std__pe5__lane30_strm0_cntl       ),      
               .std__pe5__lane30_strm0_data          ( std__pe5__lane30_strm0_data       ),      
               .std__pe5__lane30_strm0_data_valid    ( std__pe5__lane30_strm0_data_valid ),      
               .std__pe5__lane30_strm0_data_mask     ( std__pe5__lane30_strm0_data_mask  ),      

               .pe5__std__lane30_strm1_ready         ( pe5__std__lane30_strm1_ready      ),      
               .std__pe5__lane30_strm1_cntl          ( std__pe5__lane30_strm1_cntl       ),      
               .std__pe5__lane30_strm1_data          ( std__pe5__lane30_strm1_data       ),      
               .std__pe5__lane30_strm1_data_valid    ( std__pe5__lane30_strm1_data_valid ),      
               .std__pe5__lane30_strm1_data_mask     ( std__pe5__lane30_strm1_data_mask  ),      

               // PE 5, Lane 31                 
               .pe5__std__lane31_strm0_ready         ( pe5__std__lane31_strm0_ready      ),      
               .std__pe5__lane31_strm0_cntl          ( std__pe5__lane31_strm0_cntl       ),      
               .std__pe5__lane31_strm0_data          ( std__pe5__lane31_strm0_data       ),      
               .std__pe5__lane31_strm0_data_valid    ( std__pe5__lane31_strm0_data_valid ),      
               .std__pe5__lane31_strm0_data_mask     ( std__pe5__lane31_strm0_data_mask  ),      

               .pe5__std__lane31_strm1_ready         ( pe5__std__lane31_strm1_ready      ),      
               .std__pe5__lane31_strm1_cntl          ( std__pe5__lane31_strm1_cntl       ),      
               .std__pe5__lane31_strm1_data          ( std__pe5__lane31_strm1_data       ),      
               .std__pe5__lane31_strm1_data_valid    ( std__pe5__lane31_strm1_data_valid ),      
               .std__pe5__lane31_strm1_data_mask     ( std__pe5__lane31_strm1_data_mask  ),      

               // PE 6, Lane 0                 
               .pe6__std__lane0_strm0_ready         ( pe6__std__lane0_strm0_ready      ),      
               .std__pe6__lane0_strm0_cntl          ( std__pe6__lane0_strm0_cntl       ),      
               .std__pe6__lane0_strm0_data          ( std__pe6__lane0_strm0_data       ),      
               .std__pe6__lane0_strm0_data_valid    ( std__pe6__lane0_strm0_data_valid ),      
               .std__pe6__lane0_strm0_data_mask     ( std__pe6__lane0_strm0_data_mask  ),      

               .pe6__std__lane0_strm1_ready         ( pe6__std__lane0_strm1_ready      ),      
               .std__pe6__lane0_strm1_cntl          ( std__pe6__lane0_strm1_cntl       ),      
               .std__pe6__lane0_strm1_data          ( std__pe6__lane0_strm1_data       ),      
               .std__pe6__lane0_strm1_data_valid    ( std__pe6__lane0_strm1_data_valid ),      
               .std__pe6__lane0_strm1_data_mask     ( std__pe6__lane0_strm1_data_mask  ),      

               // PE 6, Lane 1                 
               .pe6__std__lane1_strm0_ready         ( pe6__std__lane1_strm0_ready      ),      
               .std__pe6__lane1_strm0_cntl          ( std__pe6__lane1_strm0_cntl       ),      
               .std__pe6__lane1_strm0_data          ( std__pe6__lane1_strm0_data       ),      
               .std__pe6__lane1_strm0_data_valid    ( std__pe6__lane1_strm0_data_valid ),      
               .std__pe6__lane1_strm0_data_mask     ( std__pe6__lane1_strm0_data_mask  ),      

               .pe6__std__lane1_strm1_ready         ( pe6__std__lane1_strm1_ready      ),      
               .std__pe6__lane1_strm1_cntl          ( std__pe6__lane1_strm1_cntl       ),      
               .std__pe6__lane1_strm1_data          ( std__pe6__lane1_strm1_data       ),      
               .std__pe6__lane1_strm1_data_valid    ( std__pe6__lane1_strm1_data_valid ),      
               .std__pe6__lane1_strm1_data_mask     ( std__pe6__lane1_strm1_data_mask  ),      

               // PE 6, Lane 2                 
               .pe6__std__lane2_strm0_ready         ( pe6__std__lane2_strm0_ready      ),      
               .std__pe6__lane2_strm0_cntl          ( std__pe6__lane2_strm0_cntl       ),      
               .std__pe6__lane2_strm0_data          ( std__pe6__lane2_strm0_data       ),      
               .std__pe6__lane2_strm0_data_valid    ( std__pe6__lane2_strm0_data_valid ),      
               .std__pe6__lane2_strm0_data_mask     ( std__pe6__lane2_strm0_data_mask  ),      

               .pe6__std__lane2_strm1_ready         ( pe6__std__lane2_strm1_ready      ),      
               .std__pe6__lane2_strm1_cntl          ( std__pe6__lane2_strm1_cntl       ),      
               .std__pe6__lane2_strm1_data          ( std__pe6__lane2_strm1_data       ),      
               .std__pe6__lane2_strm1_data_valid    ( std__pe6__lane2_strm1_data_valid ),      
               .std__pe6__lane2_strm1_data_mask     ( std__pe6__lane2_strm1_data_mask  ),      

               // PE 6, Lane 3                 
               .pe6__std__lane3_strm0_ready         ( pe6__std__lane3_strm0_ready      ),      
               .std__pe6__lane3_strm0_cntl          ( std__pe6__lane3_strm0_cntl       ),      
               .std__pe6__lane3_strm0_data          ( std__pe6__lane3_strm0_data       ),      
               .std__pe6__lane3_strm0_data_valid    ( std__pe6__lane3_strm0_data_valid ),      
               .std__pe6__lane3_strm0_data_mask     ( std__pe6__lane3_strm0_data_mask  ),      

               .pe6__std__lane3_strm1_ready         ( pe6__std__lane3_strm1_ready      ),      
               .std__pe6__lane3_strm1_cntl          ( std__pe6__lane3_strm1_cntl       ),      
               .std__pe6__lane3_strm1_data          ( std__pe6__lane3_strm1_data       ),      
               .std__pe6__lane3_strm1_data_valid    ( std__pe6__lane3_strm1_data_valid ),      
               .std__pe6__lane3_strm1_data_mask     ( std__pe6__lane3_strm1_data_mask  ),      

               // PE 6, Lane 4                 
               .pe6__std__lane4_strm0_ready         ( pe6__std__lane4_strm0_ready      ),      
               .std__pe6__lane4_strm0_cntl          ( std__pe6__lane4_strm0_cntl       ),      
               .std__pe6__lane4_strm0_data          ( std__pe6__lane4_strm0_data       ),      
               .std__pe6__lane4_strm0_data_valid    ( std__pe6__lane4_strm0_data_valid ),      
               .std__pe6__lane4_strm0_data_mask     ( std__pe6__lane4_strm0_data_mask  ),      

               .pe6__std__lane4_strm1_ready         ( pe6__std__lane4_strm1_ready      ),      
               .std__pe6__lane4_strm1_cntl          ( std__pe6__lane4_strm1_cntl       ),      
               .std__pe6__lane4_strm1_data          ( std__pe6__lane4_strm1_data       ),      
               .std__pe6__lane4_strm1_data_valid    ( std__pe6__lane4_strm1_data_valid ),      
               .std__pe6__lane4_strm1_data_mask     ( std__pe6__lane4_strm1_data_mask  ),      

               // PE 6, Lane 5                 
               .pe6__std__lane5_strm0_ready         ( pe6__std__lane5_strm0_ready      ),      
               .std__pe6__lane5_strm0_cntl          ( std__pe6__lane5_strm0_cntl       ),      
               .std__pe6__lane5_strm0_data          ( std__pe6__lane5_strm0_data       ),      
               .std__pe6__lane5_strm0_data_valid    ( std__pe6__lane5_strm0_data_valid ),      
               .std__pe6__lane5_strm0_data_mask     ( std__pe6__lane5_strm0_data_mask  ),      

               .pe6__std__lane5_strm1_ready         ( pe6__std__lane5_strm1_ready      ),      
               .std__pe6__lane5_strm1_cntl          ( std__pe6__lane5_strm1_cntl       ),      
               .std__pe6__lane5_strm1_data          ( std__pe6__lane5_strm1_data       ),      
               .std__pe6__lane5_strm1_data_valid    ( std__pe6__lane5_strm1_data_valid ),      
               .std__pe6__lane5_strm1_data_mask     ( std__pe6__lane5_strm1_data_mask  ),      

               // PE 6, Lane 6                 
               .pe6__std__lane6_strm0_ready         ( pe6__std__lane6_strm0_ready      ),      
               .std__pe6__lane6_strm0_cntl          ( std__pe6__lane6_strm0_cntl       ),      
               .std__pe6__lane6_strm0_data          ( std__pe6__lane6_strm0_data       ),      
               .std__pe6__lane6_strm0_data_valid    ( std__pe6__lane6_strm0_data_valid ),      
               .std__pe6__lane6_strm0_data_mask     ( std__pe6__lane6_strm0_data_mask  ),      

               .pe6__std__lane6_strm1_ready         ( pe6__std__lane6_strm1_ready      ),      
               .std__pe6__lane6_strm1_cntl          ( std__pe6__lane6_strm1_cntl       ),      
               .std__pe6__lane6_strm1_data          ( std__pe6__lane6_strm1_data       ),      
               .std__pe6__lane6_strm1_data_valid    ( std__pe6__lane6_strm1_data_valid ),      
               .std__pe6__lane6_strm1_data_mask     ( std__pe6__lane6_strm1_data_mask  ),      

               // PE 6, Lane 7                 
               .pe6__std__lane7_strm0_ready         ( pe6__std__lane7_strm0_ready      ),      
               .std__pe6__lane7_strm0_cntl          ( std__pe6__lane7_strm0_cntl       ),      
               .std__pe6__lane7_strm0_data          ( std__pe6__lane7_strm0_data       ),      
               .std__pe6__lane7_strm0_data_valid    ( std__pe6__lane7_strm0_data_valid ),      
               .std__pe6__lane7_strm0_data_mask     ( std__pe6__lane7_strm0_data_mask  ),      

               .pe6__std__lane7_strm1_ready         ( pe6__std__lane7_strm1_ready      ),      
               .std__pe6__lane7_strm1_cntl          ( std__pe6__lane7_strm1_cntl       ),      
               .std__pe6__lane7_strm1_data          ( std__pe6__lane7_strm1_data       ),      
               .std__pe6__lane7_strm1_data_valid    ( std__pe6__lane7_strm1_data_valid ),      
               .std__pe6__lane7_strm1_data_mask     ( std__pe6__lane7_strm1_data_mask  ),      

               // PE 6, Lane 8                 
               .pe6__std__lane8_strm0_ready         ( pe6__std__lane8_strm0_ready      ),      
               .std__pe6__lane8_strm0_cntl          ( std__pe6__lane8_strm0_cntl       ),      
               .std__pe6__lane8_strm0_data          ( std__pe6__lane8_strm0_data       ),      
               .std__pe6__lane8_strm0_data_valid    ( std__pe6__lane8_strm0_data_valid ),      
               .std__pe6__lane8_strm0_data_mask     ( std__pe6__lane8_strm0_data_mask  ),      

               .pe6__std__lane8_strm1_ready         ( pe6__std__lane8_strm1_ready      ),      
               .std__pe6__lane8_strm1_cntl          ( std__pe6__lane8_strm1_cntl       ),      
               .std__pe6__lane8_strm1_data          ( std__pe6__lane8_strm1_data       ),      
               .std__pe6__lane8_strm1_data_valid    ( std__pe6__lane8_strm1_data_valid ),      
               .std__pe6__lane8_strm1_data_mask     ( std__pe6__lane8_strm1_data_mask  ),      

               // PE 6, Lane 9                 
               .pe6__std__lane9_strm0_ready         ( pe6__std__lane9_strm0_ready      ),      
               .std__pe6__lane9_strm0_cntl          ( std__pe6__lane9_strm0_cntl       ),      
               .std__pe6__lane9_strm0_data          ( std__pe6__lane9_strm0_data       ),      
               .std__pe6__lane9_strm0_data_valid    ( std__pe6__lane9_strm0_data_valid ),      
               .std__pe6__lane9_strm0_data_mask     ( std__pe6__lane9_strm0_data_mask  ),      

               .pe6__std__lane9_strm1_ready         ( pe6__std__lane9_strm1_ready      ),      
               .std__pe6__lane9_strm1_cntl          ( std__pe6__lane9_strm1_cntl       ),      
               .std__pe6__lane9_strm1_data          ( std__pe6__lane9_strm1_data       ),      
               .std__pe6__lane9_strm1_data_valid    ( std__pe6__lane9_strm1_data_valid ),      
               .std__pe6__lane9_strm1_data_mask     ( std__pe6__lane9_strm1_data_mask  ),      

               // PE 6, Lane 10                 
               .pe6__std__lane10_strm0_ready         ( pe6__std__lane10_strm0_ready      ),      
               .std__pe6__lane10_strm0_cntl          ( std__pe6__lane10_strm0_cntl       ),      
               .std__pe6__lane10_strm0_data          ( std__pe6__lane10_strm0_data       ),      
               .std__pe6__lane10_strm0_data_valid    ( std__pe6__lane10_strm0_data_valid ),      
               .std__pe6__lane10_strm0_data_mask     ( std__pe6__lane10_strm0_data_mask  ),      

               .pe6__std__lane10_strm1_ready         ( pe6__std__lane10_strm1_ready      ),      
               .std__pe6__lane10_strm1_cntl          ( std__pe6__lane10_strm1_cntl       ),      
               .std__pe6__lane10_strm1_data          ( std__pe6__lane10_strm1_data       ),      
               .std__pe6__lane10_strm1_data_valid    ( std__pe6__lane10_strm1_data_valid ),      
               .std__pe6__lane10_strm1_data_mask     ( std__pe6__lane10_strm1_data_mask  ),      

               // PE 6, Lane 11                 
               .pe6__std__lane11_strm0_ready         ( pe6__std__lane11_strm0_ready      ),      
               .std__pe6__lane11_strm0_cntl          ( std__pe6__lane11_strm0_cntl       ),      
               .std__pe6__lane11_strm0_data          ( std__pe6__lane11_strm0_data       ),      
               .std__pe6__lane11_strm0_data_valid    ( std__pe6__lane11_strm0_data_valid ),      
               .std__pe6__lane11_strm0_data_mask     ( std__pe6__lane11_strm0_data_mask  ),      

               .pe6__std__lane11_strm1_ready         ( pe6__std__lane11_strm1_ready      ),      
               .std__pe6__lane11_strm1_cntl          ( std__pe6__lane11_strm1_cntl       ),      
               .std__pe6__lane11_strm1_data          ( std__pe6__lane11_strm1_data       ),      
               .std__pe6__lane11_strm1_data_valid    ( std__pe6__lane11_strm1_data_valid ),      
               .std__pe6__lane11_strm1_data_mask     ( std__pe6__lane11_strm1_data_mask  ),      

               // PE 6, Lane 12                 
               .pe6__std__lane12_strm0_ready         ( pe6__std__lane12_strm0_ready      ),      
               .std__pe6__lane12_strm0_cntl          ( std__pe6__lane12_strm0_cntl       ),      
               .std__pe6__lane12_strm0_data          ( std__pe6__lane12_strm0_data       ),      
               .std__pe6__lane12_strm0_data_valid    ( std__pe6__lane12_strm0_data_valid ),      
               .std__pe6__lane12_strm0_data_mask     ( std__pe6__lane12_strm0_data_mask  ),      

               .pe6__std__lane12_strm1_ready         ( pe6__std__lane12_strm1_ready      ),      
               .std__pe6__lane12_strm1_cntl          ( std__pe6__lane12_strm1_cntl       ),      
               .std__pe6__lane12_strm1_data          ( std__pe6__lane12_strm1_data       ),      
               .std__pe6__lane12_strm1_data_valid    ( std__pe6__lane12_strm1_data_valid ),      
               .std__pe6__lane12_strm1_data_mask     ( std__pe6__lane12_strm1_data_mask  ),      

               // PE 6, Lane 13                 
               .pe6__std__lane13_strm0_ready         ( pe6__std__lane13_strm0_ready      ),      
               .std__pe6__lane13_strm0_cntl          ( std__pe6__lane13_strm0_cntl       ),      
               .std__pe6__lane13_strm0_data          ( std__pe6__lane13_strm0_data       ),      
               .std__pe6__lane13_strm0_data_valid    ( std__pe6__lane13_strm0_data_valid ),      
               .std__pe6__lane13_strm0_data_mask     ( std__pe6__lane13_strm0_data_mask  ),      

               .pe6__std__lane13_strm1_ready         ( pe6__std__lane13_strm1_ready      ),      
               .std__pe6__lane13_strm1_cntl          ( std__pe6__lane13_strm1_cntl       ),      
               .std__pe6__lane13_strm1_data          ( std__pe6__lane13_strm1_data       ),      
               .std__pe6__lane13_strm1_data_valid    ( std__pe6__lane13_strm1_data_valid ),      
               .std__pe6__lane13_strm1_data_mask     ( std__pe6__lane13_strm1_data_mask  ),      

               // PE 6, Lane 14                 
               .pe6__std__lane14_strm0_ready         ( pe6__std__lane14_strm0_ready      ),      
               .std__pe6__lane14_strm0_cntl          ( std__pe6__lane14_strm0_cntl       ),      
               .std__pe6__lane14_strm0_data          ( std__pe6__lane14_strm0_data       ),      
               .std__pe6__lane14_strm0_data_valid    ( std__pe6__lane14_strm0_data_valid ),      
               .std__pe6__lane14_strm0_data_mask     ( std__pe6__lane14_strm0_data_mask  ),      

               .pe6__std__lane14_strm1_ready         ( pe6__std__lane14_strm1_ready      ),      
               .std__pe6__lane14_strm1_cntl          ( std__pe6__lane14_strm1_cntl       ),      
               .std__pe6__lane14_strm1_data          ( std__pe6__lane14_strm1_data       ),      
               .std__pe6__lane14_strm1_data_valid    ( std__pe6__lane14_strm1_data_valid ),      
               .std__pe6__lane14_strm1_data_mask     ( std__pe6__lane14_strm1_data_mask  ),      

               // PE 6, Lane 15                 
               .pe6__std__lane15_strm0_ready         ( pe6__std__lane15_strm0_ready      ),      
               .std__pe6__lane15_strm0_cntl          ( std__pe6__lane15_strm0_cntl       ),      
               .std__pe6__lane15_strm0_data          ( std__pe6__lane15_strm0_data       ),      
               .std__pe6__lane15_strm0_data_valid    ( std__pe6__lane15_strm0_data_valid ),      
               .std__pe6__lane15_strm0_data_mask     ( std__pe6__lane15_strm0_data_mask  ),      

               .pe6__std__lane15_strm1_ready         ( pe6__std__lane15_strm1_ready      ),      
               .std__pe6__lane15_strm1_cntl          ( std__pe6__lane15_strm1_cntl       ),      
               .std__pe6__lane15_strm1_data          ( std__pe6__lane15_strm1_data       ),      
               .std__pe6__lane15_strm1_data_valid    ( std__pe6__lane15_strm1_data_valid ),      
               .std__pe6__lane15_strm1_data_mask     ( std__pe6__lane15_strm1_data_mask  ),      

               // PE 6, Lane 16                 
               .pe6__std__lane16_strm0_ready         ( pe6__std__lane16_strm0_ready      ),      
               .std__pe6__lane16_strm0_cntl          ( std__pe6__lane16_strm0_cntl       ),      
               .std__pe6__lane16_strm0_data          ( std__pe6__lane16_strm0_data       ),      
               .std__pe6__lane16_strm0_data_valid    ( std__pe6__lane16_strm0_data_valid ),      
               .std__pe6__lane16_strm0_data_mask     ( std__pe6__lane16_strm0_data_mask  ),      

               .pe6__std__lane16_strm1_ready         ( pe6__std__lane16_strm1_ready      ),      
               .std__pe6__lane16_strm1_cntl          ( std__pe6__lane16_strm1_cntl       ),      
               .std__pe6__lane16_strm1_data          ( std__pe6__lane16_strm1_data       ),      
               .std__pe6__lane16_strm1_data_valid    ( std__pe6__lane16_strm1_data_valid ),      
               .std__pe6__lane16_strm1_data_mask     ( std__pe6__lane16_strm1_data_mask  ),      

               // PE 6, Lane 17                 
               .pe6__std__lane17_strm0_ready         ( pe6__std__lane17_strm0_ready      ),      
               .std__pe6__lane17_strm0_cntl          ( std__pe6__lane17_strm0_cntl       ),      
               .std__pe6__lane17_strm0_data          ( std__pe6__lane17_strm0_data       ),      
               .std__pe6__lane17_strm0_data_valid    ( std__pe6__lane17_strm0_data_valid ),      
               .std__pe6__lane17_strm0_data_mask     ( std__pe6__lane17_strm0_data_mask  ),      

               .pe6__std__lane17_strm1_ready         ( pe6__std__lane17_strm1_ready      ),      
               .std__pe6__lane17_strm1_cntl          ( std__pe6__lane17_strm1_cntl       ),      
               .std__pe6__lane17_strm1_data          ( std__pe6__lane17_strm1_data       ),      
               .std__pe6__lane17_strm1_data_valid    ( std__pe6__lane17_strm1_data_valid ),      
               .std__pe6__lane17_strm1_data_mask     ( std__pe6__lane17_strm1_data_mask  ),      

               // PE 6, Lane 18                 
               .pe6__std__lane18_strm0_ready         ( pe6__std__lane18_strm0_ready      ),      
               .std__pe6__lane18_strm0_cntl          ( std__pe6__lane18_strm0_cntl       ),      
               .std__pe6__lane18_strm0_data          ( std__pe6__lane18_strm0_data       ),      
               .std__pe6__lane18_strm0_data_valid    ( std__pe6__lane18_strm0_data_valid ),      
               .std__pe6__lane18_strm0_data_mask     ( std__pe6__lane18_strm0_data_mask  ),      

               .pe6__std__lane18_strm1_ready         ( pe6__std__lane18_strm1_ready      ),      
               .std__pe6__lane18_strm1_cntl          ( std__pe6__lane18_strm1_cntl       ),      
               .std__pe6__lane18_strm1_data          ( std__pe6__lane18_strm1_data       ),      
               .std__pe6__lane18_strm1_data_valid    ( std__pe6__lane18_strm1_data_valid ),      
               .std__pe6__lane18_strm1_data_mask     ( std__pe6__lane18_strm1_data_mask  ),      

               // PE 6, Lane 19                 
               .pe6__std__lane19_strm0_ready         ( pe6__std__lane19_strm0_ready      ),      
               .std__pe6__lane19_strm0_cntl          ( std__pe6__lane19_strm0_cntl       ),      
               .std__pe6__lane19_strm0_data          ( std__pe6__lane19_strm0_data       ),      
               .std__pe6__lane19_strm0_data_valid    ( std__pe6__lane19_strm0_data_valid ),      
               .std__pe6__lane19_strm0_data_mask     ( std__pe6__lane19_strm0_data_mask  ),      

               .pe6__std__lane19_strm1_ready         ( pe6__std__lane19_strm1_ready      ),      
               .std__pe6__lane19_strm1_cntl          ( std__pe6__lane19_strm1_cntl       ),      
               .std__pe6__lane19_strm1_data          ( std__pe6__lane19_strm1_data       ),      
               .std__pe6__lane19_strm1_data_valid    ( std__pe6__lane19_strm1_data_valid ),      
               .std__pe6__lane19_strm1_data_mask     ( std__pe6__lane19_strm1_data_mask  ),      

               // PE 6, Lane 20                 
               .pe6__std__lane20_strm0_ready         ( pe6__std__lane20_strm0_ready      ),      
               .std__pe6__lane20_strm0_cntl          ( std__pe6__lane20_strm0_cntl       ),      
               .std__pe6__lane20_strm0_data          ( std__pe6__lane20_strm0_data       ),      
               .std__pe6__lane20_strm0_data_valid    ( std__pe6__lane20_strm0_data_valid ),      
               .std__pe6__lane20_strm0_data_mask     ( std__pe6__lane20_strm0_data_mask  ),      

               .pe6__std__lane20_strm1_ready         ( pe6__std__lane20_strm1_ready      ),      
               .std__pe6__lane20_strm1_cntl          ( std__pe6__lane20_strm1_cntl       ),      
               .std__pe6__lane20_strm1_data          ( std__pe6__lane20_strm1_data       ),      
               .std__pe6__lane20_strm1_data_valid    ( std__pe6__lane20_strm1_data_valid ),      
               .std__pe6__lane20_strm1_data_mask     ( std__pe6__lane20_strm1_data_mask  ),      

               // PE 6, Lane 21                 
               .pe6__std__lane21_strm0_ready         ( pe6__std__lane21_strm0_ready      ),      
               .std__pe6__lane21_strm0_cntl          ( std__pe6__lane21_strm0_cntl       ),      
               .std__pe6__lane21_strm0_data          ( std__pe6__lane21_strm0_data       ),      
               .std__pe6__lane21_strm0_data_valid    ( std__pe6__lane21_strm0_data_valid ),      
               .std__pe6__lane21_strm0_data_mask     ( std__pe6__lane21_strm0_data_mask  ),      

               .pe6__std__lane21_strm1_ready         ( pe6__std__lane21_strm1_ready      ),      
               .std__pe6__lane21_strm1_cntl          ( std__pe6__lane21_strm1_cntl       ),      
               .std__pe6__lane21_strm1_data          ( std__pe6__lane21_strm1_data       ),      
               .std__pe6__lane21_strm1_data_valid    ( std__pe6__lane21_strm1_data_valid ),      
               .std__pe6__lane21_strm1_data_mask     ( std__pe6__lane21_strm1_data_mask  ),      

               // PE 6, Lane 22                 
               .pe6__std__lane22_strm0_ready         ( pe6__std__lane22_strm0_ready      ),      
               .std__pe6__lane22_strm0_cntl          ( std__pe6__lane22_strm0_cntl       ),      
               .std__pe6__lane22_strm0_data          ( std__pe6__lane22_strm0_data       ),      
               .std__pe6__lane22_strm0_data_valid    ( std__pe6__lane22_strm0_data_valid ),      
               .std__pe6__lane22_strm0_data_mask     ( std__pe6__lane22_strm0_data_mask  ),      

               .pe6__std__lane22_strm1_ready         ( pe6__std__lane22_strm1_ready      ),      
               .std__pe6__lane22_strm1_cntl          ( std__pe6__lane22_strm1_cntl       ),      
               .std__pe6__lane22_strm1_data          ( std__pe6__lane22_strm1_data       ),      
               .std__pe6__lane22_strm1_data_valid    ( std__pe6__lane22_strm1_data_valid ),      
               .std__pe6__lane22_strm1_data_mask     ( std__pe6__lane22_strm1_data_mask  ),      

               // PE 6, Lane 23                 
               .pe6__std__lane23_strm0_ready         ( pe6__std__lane23_strm0_ready      ),      
               .std__pe6__lane23_strm0_cntl          ( std__pe6__lane23_strm0_cntl       ),      
               .std__pe6__lane23_strm0_data          ( std__pe6__lane23_strm0_data       ),      
               .std__pe6__lane23_strm0_data_valid    ( std__pe6__lane23_strm0_data_valid ),      
               .std__pe6__lane23_strm0_data_mask     ( std__pe6__lane23_strm0_data_mask  ),      

               .pe6__std__lane23_strm1_ready         ( pe6__std__lane23_strm1_ready      ),      
               .std__pe6__lane23_strm1_cntl          ( std__pe6__lane23_strm1_cntl       ),      
               .std__pe6__lane23_strm1_data          ( std__pe6__lane23_strm1_data       ),      
               .std__pe6__lane23_strm1_data_valid    ( std__pe6__lane23_strm1_data_valid ),      
               .std__pe6__lane23_strm1_data_mask     ( std__pe6__lane23_strm1_data_mask  ),      

               // PE 6, Lane 24                 
               .pe6__std__lane24_strm0_ready         ( pe6__std__lane24_strm0_ready      ),      
               .std__pe6__lane24_strm0_cntl          ( std__pe6__lane24_strm0_cntl       ),      
               .std__pe6__lane24_strm0_data          ( std__pe6__lane24_strm0_data       ),      
               .std__pe6__lane24_strm0_data_valid    ( std__pe6__lane24_strm0_data_valid ),      
               .std__pe6__lane24_strm0_data_mask     ( std__pe6__lane24_strm0_data_mask  ),      

               .pe6__std__lane24_strm1_ready         ( pe6__std__lane24_strm1_ready      ),      
               .std__pe6__lane24_strm1_cntl          ( std__pe6__lane24_strm1_cntl       ),      
               .std__pe6__lane24_strm1_data          ( std__pe6__lane24_strm1_data       ),      
               .std__pe6__lane24_strm1_data_valid    ( std__pe6__lane24_strm1_data_valid ),      
               .std__pe6__lane24_strm1_data_mask     ( std__pe6__lane24_strm1_data_mask  ),      

               // PE 6, Lane 25                 
               .pe6__std__lane25_strm0_ready         ( pe6__std__lane25_strm0_ready      ),      
               .std__pe6__lane25_strm0_cntl          ( std__pe6__lane25_strm0_cntl       ),      
               .std__pe6__lane25_strm0_data          ( std__pe6__lane25_strm0_data       ),      
               .std__pe6__lane25_strm0_data_valid    ( std__pe6__lane25_strm0_data_valid ),      
               .std__pe6__lane25_strm0_data_mask     ( std__pe6__lane25_strm0_data_mask  ),      

               .pe6__std__lane25_strm1_ready         ( pe6__std__lane25_strm1_ready      ),      
               .std__pe6__lane25_strm1_cntl          ( std__pe6__lane25_strm1_cntl       ),      
               .std__pe6__lane25_strm1_data          ( std__pe6__lane25_strm1_data       ),      
               .std__pe6__lane25_strm1_data_valid    ( std__pe6__lane25_strm1_data_valid ),      
               .std__pe6__lane25_strm1_data_mask     ( std__pe6__lane25_strm1_data_mask  ),      

               // PE 6, Lane 26                 
               .pe6__std__lane26_strm0_ready         ( pe6__std__lane26_strm0_ready      ),      
               .std__pe6__lane26_strm0_cntl          ( std__pe6__lane26_strm0_cntl       ),      
               .std__pe6__lane26_strm0_data          ( std__pe6__lane26_strm0_data       ),      
               .std__pe6__lane26_strm0_data_valid    ( std__pe6__lane26_strm0_data_valid ),      
               .std__pe6__lane26_strm0_data_mask     ( std__pe6__lane26_strm0_data_mask  ),      

               .pe6__std__lane26_strm1_ready         ( pe6__std__lane26_strm1_ready      ),      
               .std__pe6__lane26_strm1_cntl          ( std__pe6__lane26_strm1_cntl       ),      
               .std__pe6__lane26_strm1_data          ( std__pe6__lane26_strm1_data       ),      
               .std__pe6__lane26_strm1_data_valid    ( std__pe6__lane26_strm1_data_valid ),      
               .std__pe6__lane26_strm1_data_mask     ( std__pe6__lane26_strm1_data_mask  ),      

               // PE 6, Lane 27                 
               .pe6__std__lane27_strm0_ready         ( pe6__std__lane27_strm0_ready      ),      
               .std__pe6__lane27_strm0_cntl          ( std__pe6__lane27_strm0_cntl       ),      
               .std__pe6__lane27_strm0_data          ( std__pe6__lane27_strm0_data       ),      
               .std__pe6__lane27_strm0_data_valid    ( std__pe6__lane27_strm0_data_valid ),      
               .std__pe6__lane27_strm0_data_mask     ( std__pe6__lane27_strm0_data_mask  ),      

               .pe6__std__lane27_strm1_ready         ( pe6__std__lane27_strm1_ready      ),      
               .std__pe6__lane27_strm1_cntl          ( std__pe6__lane27_strm1_cntl       ),      
               .std__pe6__lane27_strm1_data          ( std__pe6__lane27_strm1_data       ),      
               .std__pe6__lane27_strm1_data_valid    ( std__pe6__lane27_strm1_data_valid ),      
               .std__pe6__lane27_strm1_data_mask     ( std__pe6__lane27_strm1_data_mask  ),      

               // PE 6, Lane 28                 
               .pe6__std__lane28_strm0_ready         ( pe6__std__lane28_strm0_ready      ),      
               .std__pe6__lane28_strm0_cntl          ( std__pe6__lane28_strm0_cntl       ),      
               .std__pe6__lane28_strm0_data          ( std__pe6__lane28_strm0_data       ),      
               .std__pe6__lane28_strm0_data_valid    ( std__pe6__lane28_strm0_data_valid ),      
               .std__pe6__lane28_strm0_data_mask     ( std__pe6__lane28_strm0_data_mask  ),      

               .pe6__std__lane28_strm1_ready         ( pe6__std__lane28_strm1_ready      ),      
               .std__pe6__lane28_strm1_cntl          ( std__pe6__lane28_strm1_cntl       ),      
               .std__pe6__lane28_strm1_data          ( std__pe6__lane28_strm1_data       ),      
               .std__pe6__lane28_strm1_data_valid    ( std__pe6__lane28_strm1_data_valid ),      
               .std__pe6__lane28_strm1_data_mask     ( std__pe6__lane28_strm1_data_mask  ),      

               // PE 6, Lane 29                 
               .pe6__std__lane29_strm0_ready         ( pe6__std__lane29_strm0_ready      ),      
               .std__pe6__lane29_strm0_cntl          ( std__pe6__lane29_strm0_cntl       ),      
               .std__pe6__lane29_strm0_data          ( std__pe6__lane29_strm0_data       ),      
               .std__pe6__lane29_strm0_data_valid    ( std__pe6__lane29_strm0_data_valid ),      
               .std__pe6__lane29_strm0_data_mask     ( std__pe6__lane29_strm0_data_mask  ),      

               .pe6__std__lane29_strm1_ready         ( pe6__std__lane29_strm1_ready      ),      
               .std__pe6__lane29_strm1_cntl          ( std__pe6__lane29_strm1_cntl       ),      
               .std__pe6__lane29_strm1_data          ( std__pe6__lane29_strm1_data       ),      
               .std__pe6__lane29_strm1_data_valid    ( std__pe6__lane29_strm1_data_valid ),      
               .std__pe6__lane29_strm1_data_mask     ( std__pe6__lane29_strm1_data_mask  ),      

               // PE 6, Lane 30                 
               .pe6__std__lane30_strm0_ready         ( pe6__std__lane30_strm0_ready      ),      
               .std__pe6__lane30_strm0_cntl          ( std__pe6__lane30_strm0_cntl       ),      
               .std__pe6__lane30_strm0_data          ( std__pe6__lane30_strm0_data       ),      
               .std__pe6__lane30_strm0_data_valid    ( std__pe6__lane30_strm0_data_valid ),      
               .std__pe6__lane30_strm0_data_mask     ( std__pe6__lane30_strm0_data_mask  ),      

               .pe6__std__lane30_strm1_ready         ( pe6__std__lane30_strm1_ready      ),      
               .std__pe6__lane30_strm1_cntl          ( std__pe6__lane30_strm1_cntl       ),      
               .std__pe6__lane30_strm1_data          ( std__pe6__lane30_strm1_data       ),      
               .std__pe6__lane30_strm1_data_valid    ( std__pe6__lane30_strm1_data_valid ),      
               .std__pe6__lane30_strm1_data_mask     ( std__pe6__lane30_strm1_data_mask  ),      

               // PE 6, Lane 31                 
               .pe6__std__lane31_strm0_ready         ( pe6__std__lane31_strm0_ready      ),      
               .std__pe6__lane31_strm0_cntl          ( std__pe6__lane31_strm0_cntl       ),      
               .std__pe6__lane31_strm0_data          ( std__pe6__lane31_strm0_data       ),      
               .std__pe6__lane31_strm0_data_valid    ( std__pe6__lane31_strm0_data_valid ),      
               .std__pe6__lane31_strm0_data_mask     ( std__pe6__lane31_strm0_data_mask  ),      

               .pe6__std__lane31_strm1_ready         ( pe6__std__lane31_strm1_ready      ),      
               .std__pe6__lane31_strm1_cntl          ( std__pe6__lane31_strm1_cntl       ),      
               .std__pe6__lane31_strm1_data          ( std__pe6__lane31_strm1_data       ),      
               .std__pe6__lane31_strm1_data_valid    ( std__pe6__lane31_strm1_data_valid ),      
               .std__pe6__lane31_strm1_data_mask     ( std__pe6__lane31_strm1_data_mask  ),      

               // PE 7, Lane 0                 
               .pe7__std__lane0_strm0_ready         ( pe7__std__lane0_strm0_ready      ),      
               .std__pe7__lane0_strm0_cntl          ( std__pe7__lane0_strm0_cntl       ),      
               .std__pe7__lane0_strm0_data          ( std__pe7__lane0_strm0_data       ),      
               .std__pe7__lane0_strm0_data_valid    ( std__pe7__lane0_strm0_data_valid ),      
               .std__pe7__lane0_strm0_data_mask     ( std__pe7__lane0_strm0_data_mask  ),      

               .pe7__std__lane0_strm1_ready         ( pe7__std__lane0_strm1_ready      ),      
               .std__pe7__lane0_strm1_cntl          ( std__pe7__lane0_strm1_cntl       ),      
               .std__pe7__lane0_strm1_data          ( std__pe7__lane0_strm1_data       ),      
               .std__pe7__lane0_strm1_data_valid    ( std__pe7__lane0_strm1_data_valid ),      
               .std__pe7__lane0_strm1_data_mask     ( std__pe7__lane0_strm1_data_mask  ),      

               // PE 7, Lane 1                 
               .pe7__std__lane1_strm0_ready         ( pe7__std__lane1_strm0_ready      ),      
               .std__pe7__lane1_strm0_cntl          ( std__pe7__lane1_strm0_cntl       ),      
               .std__pe7__lane1_strm0_data          ( std__pe7__lane1_strm0_data       ),      
               .std__pe7__lane1_strm0_data_valid    ( std__pe7__lane1_strm0_data_valid ),      
               .std__pe7__lane1_strm0_data_mask     ( std__pe7__lane1_strm0_data_mask  ),      

               .pe7__std__lane1_strm1_ready         ( pe7__std__lane1_strm1_ready      ),      
               .std__pe7__lane1_strm1_cntl          ( std__pe7__lane1_strm1_cntl       ),      
               .std__pe7__lane1_strm1_data          ( std__pe7__lane1_strm1_data       ),      
               .std__pe7__lane1_strm1_data_valid    ( std__pe7__lane1_strm1_data_valid ),      
               .std__pe7__lane1_strm1_data_mask     ( std__pe7__lane1_strm1_data_mask  ),      

               // PE 7, Lane 2                 
               .pe7__std__lane2_strm0_ready         ( pe7__std__lane2_strm0_ready      ),      
               .std__pe7__lane2_strm0_cntl          ( std__pe7__lane2_strm0_cntl       ),      
               .std__pe7__lane2_strm0_data          ( std__pe7__lane2_strm0_data       ),      
               .std__pe7__lane2_strm0_data_valid    ( std__pe7__lane2_strm0_data_valid ),      
               .std__pe7__lane2_strm0_data_mask     ( std__pe7__lane2_strm0_data_mask  ),      

               .pe7__std__lane2_strm1_ready         ( pe7__std__lane2_strm1_ready      ),      
               .std__pe7__lane2_strm1_cntl          ( std__pe7__lane2_strm1_cntl       ),      
               .std__pe7__lane2_strm1_data          ( std__pe7__lane2_strm1_data       ),      
               .std__pe7__lane2_strm1_data_valid    ( std__pe7__lane2_strm1_data_valid ),      
               .std__pe7__lane2_strm1_data_mask     ( std__pe7__lane2_strm1_data_mask  ),      

               // PE 7, Lane 3                 
               .pe7__std__lane3_strm0_ready         ( pe7__std__lane3_strm0_ready      ),      
               .std__pe7__lane3_strm0_cntl          ( std__pe7__lane3_strm0_cntl       ),      
               .std__pe7__lane3_strm0_data          ( std__pe7__lane3_strm0_data       ),      
               .std__pe7__lane3_strm0_data_valid    ( std__pe7__lane3_strm0_data_valid ),      
               .std__pe7__lane3_strm0_data_mask     ( std__pe7__lane3_strm0_data_mask  ),      

               .pe7__std__lane3_strm1_ready         ( pe7__std__lane3_strm1_ready      ),      
               .std__pe7__lane3_strm1_cntl          ( std__pe7__lane3_strm1_cntl       ),      
               .std__pe7__lane3_strm1_data          ( std__pe7__lane3_strm1_data       ),      
               .std__pe7__lane3_strm1_data_valid    ( std__pe7__lane3_strm1_data_valid ),      
               .std__pe7__lane3_strm1_data_mask     ( std__pe7__lane3_strm1_data_mask  ),      

               // PE 7, Lane 4                 
               .pe7__std__lane4_strm0_ready         ( pe7__std__lane4_strm0_ready      ),      
               .std__pe7__lane4_strm0_cntl          ( std__pe7__lane4_strm0_cntl       ),      
               .std__pe7__lane4_strm0_data          ( std__pe7__lane4_strm0_data       ),      
               .std__pe7__lane4_strm0_data_valid    ( std__pe7__lane4_strm0_data_valid ),      
               .std__pe7__lane4_strm0_data_mask     ( std__pe7__lane4_strm0_data_mask  ),      

               .pe7__std__lane4_strm1_ready         ( pe7__std__lane4_strm1_ready      ),      
               .std__pe7__lane4_strm1_cntl          ( std__pe7__lane4_strm1_cntl       ),      
               .std__pe7__lane4_strm1_data          ( std__pe7__lane4_strm1_data       ),      
               .std__pe7__lane4_strm1_data_valid    ( std__pe7__lane4_strm1_data_valid ),      
               .std__pe7__lane4_strm1_data_mask     ( std__pe7__lane4_strm1_data_mask  ),      

               // PE 7, Lane 5                 
               .pe7__std__lane5_strm0_ready         ( pe7__std__lane5_strm0_ready      ),      
               .std__pe7__lane5_strm0_cntl          ( std__pe7__lane5_strm0_cntl       ),      
               .std__pe7__lane5_strm0_data          ( std__pe7__lane5_strm0_data       ),      
               .std__pe7__lane5_strm0_data_valid    ( std__pe7__lane5_strm0_data_valid ),      
               .std__pe7__lane5_strm0_data_mask     ( std__pe7__lane5_strm0_data_mask  ),      

               .pe7__std__lane5_strm1_ready         ( pe7__std__lane5_strm1_ready      ),      
               .std__pe7__lane5_strm1_cntl          ( std__pe7__lane5_strm1_cntl       ),      
               .std__pe7__lane5_strm1_data          ( std__pe7__lane5_strm1_data       ),      
               .std__pe7__lane5_strm1_data_valid    ( std__pe7__lane5_strm1_data_valid ),      
               .std__pe7__lane5_strm1_data_mask     ( std__pe7__lane5_strm1_data_mask  ),      

               // PE 7, Lane 6                 
               .pe7__std__lane6_strm0_ready         ( pe7__std__lane6_strm0_ready      ),      
               .std__pe7__lane6_strm0_cntl          ( std__pe7__lane6_strm0_cntl       ),      
               .std__pe7__lane6_strm0_data          ( std__pe7__lane6_strm0_data       ),      
               .std__pe7__lane6_strm0_data_valid    ( std__pe7__lane6_strm0_data_valid ),      
               .std__pe7__lane6_strm0_data_mask     ( std__pe7__lane6_strm0_data_mask  ),      

               .pe7__std__lane6_strm1_ready         ( pe7__std__lane6_strm1_ready      ),      
               .std__pe7__lane6_strm1_cntl          ( std__pe7__lane6_strm1_cntl       ),      
               .std__pe7__lane6_strm1_data          ( std__pe7__lane6_strm1_data       ),      
               .std__pe7__lane6_strm1_data_valid    ( std__pe7__lane6_strm1_data_valid ),      
               .std__pe7__lane6_strm1_data_mask     ( std__pe7__lane6_strm1_data_mask  ),      

               // PE 7, Lane 7                 
               .pe7__std__lane7_strm0_ready         ( pe7__std__lane7_strm0_ready      ),      
               .std__pe7__lane7_strm0_cntl          ( std__pe7__lane7_strm0_cntl       ),      
               .std__pe7__lane7_strm0_data          ( std__pe7__lane7_strm0_data       ),      
               .std__pe7__lane7_strm0_data_valid    ( std__pe7__lane7_strm0_data_valid ),      
               .std__pe7__lane7_strm0_data_mask     ( std__pe7__lane7_strm0_data_mask  ),      

               .pe7__std__lane7_strm1_ready         ( pe7__std__lane7_strm1_ready      ),      
               .std__pe7__lane7_strm1_cntl          ( std__pe7__lane7_strm1_cntl       ),      
               .std__pe7__lane7_strm1_data          ( std__pe7__lane7_strm1_data       ),      
               .std__pe7__lane7_strm1_data_valid    ( std__pe7__lane7_strm1_data_valid ),      
               .std__pe7__lane7_strm1_data_mask     ( std__pe7__lane7_strm1_data_mask  ),      

               // PE 7, Lane 8                 
               .pe7__std__lane8_strm0_ready         ( pe7__std__lane8_strm0_ready      ),      
               .std__pe7__lane8_strm0_cntl          ( std__pe7__lane8_strm0_cntl       ),      
               .std__pe7__lane8_strm0_data          ( std__pe7__lane8_strm0_data       ),      
               .std__pe7__lane8_strm0_data_valid    ( std__pe7__lane8_strm0_data_valid ),      
               .std__pe7__lane8_strm0_data_mask     ( std__pe7__lane8_strm0_data_mask  ),      

               .pe7__std__lane8_strm1_ready         ( pe7__std__lane8_strm1_ready      ),      
               .std__pe7__lane8_strm1_cntl          ( std__pe7__lane8_strm1_cntl       ),      
               .std__pe7__lane8_strm1_data          ( std__pe7__lane8_strm1_data       ),      
               .std__pe7__lane8_strm1_data_valid    ( std__pe7__lane8_strm1_data_valid ),      
               .std__pe7__lane8_strm1_data_mask     ( std__pe7__lane8_strm1_data_mask  ),      

               // PE 7, Lane 9                 
               .pe7__std__lane9_strm0_ready         ( pe7__std__lane9_strm0_ready      ),      
               .std__pe7__lane9_strm0_cntl          ( std__pe7__lane9_strm0_cntl       ),      
               .std__pe7__lane9_strm0_data          ( std__pe7__lane9_strm0_data       ),      
               .std__pe7__lane9_strm0_data_valid    ( std__pe7__lane9_strm0_data_valid ),      
               .std__pe7__lane9_strm0_data_mask     ( std__pe7__lane9_strm0_data_mask  ),      

               .pe7__std__lane9_strm1_ready         ( pe7__std__lane9_strm1_ready      ),      
               .std__pe7__lane9_strm1_cntl          ( std__pe7__lane9_strm1_cntl       ),      
               .std__pe7__lane9_strm1_data          ( std__pe7__lane9_strm1_data       ),      
               .std__pe7__lane9_strm1_data_valid    ( std__pe7__lane9_strm1_data_valid ),      
               .std__pe7__lane9_strm1_data_mask     ( std__pe7__lane9_strm1_data_mask  ),      

               // PE 7, Lane 10                 
               .pe7__std__lane10_strm0_ready         ( pe7__std__lane10_strm0_ready      ),      
               .std__pe7__lane10_strm0_cntl          ( std__pe7__lane10_strm0_cntl       ),      
               .std__pe7__lane10_strm0_data          ( std__pe7__lane10_strm0_data       ),      
               .std__pe7__lane10_strm0_data_valid    ( std__pe7__lane10_strm0_data_valid ),      
               .std__pe7__lane10_strm0_data_mask     ( std__pe7__lane10_strm0_data_mask  ),      

               .pe7__std__lane10_strm1_ready         ( pe7__std__lane10_strm1_ready      ),      
               .std__pe7__lane10_strm1_cntl          ( std__pe7__lane10_strm1_cntl       ),      
               .std__pe7__lane10_strm1_data          ( std__pe7__lane10_strm1_data       ),      
               .std__pe7__lane10_strm1_data_valid    ( std__pe7__lane10_strm1_data_valid ),      
               .std__pe7__lane10_strm1_data_mask     ( std__pe7__lane10_strm1_data_mask  ),      

               // PE 7, Lane 11                 
               .pe7__std__lane11_strm0_ready         ( pe7__std__lane11_strm0_ready      ),      
               .std__pe7__lane11_strm0_cntl          ( std__pe7__lane11_strm0_cntl       ),      
               .std__pe7__lane11_strm0_data          ( std__pe7__lane11_strm0_data       ),      
               .std__pe7__lane11_strm0_data_valid    ( std__pe7__lane11_strm0_data_valid ),      
               .std__pe7__lane11_strm0_data_mask     ( std__pe7__lane11_strm0_data_mask  ),      

               .pe7__std__lane11_strm1_ready         ( pe7__std__lane11_strm1_ready      ),      
               .std__pe7__lane11_strm1_cntl          ( std__pe7__lane11_strm1_cntl       ),      
               .std__pe7__lane11_strm1_data          ( std__pe7__lane11_strm1_data       ),      
               .std__pe7__lane11_strm1_data_valid    ( std__pe7__lane11_strm1_data_valid ),      
               .std__pe7__lane11_strm1_data_mask     ( std__pe7__lane11_strm1_data_mask  ),      

               // PE 7, Lane 12                 
               .pe7__std__lane12_strm0_ready         ( pe7__std__lane12_strm0_ready      ),      
               .std__pe7__lane12_strm0_cntl          ( std__pe7__lane12_strm0_cntl       ),      
               .std__pe7__lane12_strm0_data          ( std__pe7__lane12_strm0_data       ),      
               .std__pe7__lane12_strm0_data_valid    ( std__pe7__lane12_strm0_data_valid ),      
               .std__pe7__lane12_strm0_data_mask     ( std__pe7__lane12_strm0_data_mask  ),      

               .pe7__std__lane12_strm1_ready         ( pe7__std__lane12_strm1_ready      ),      
               .std__pe7__lane12_strm1_cntl          ( std__pe7__lane12_strm1_cntl       ),      
               .std__pe7__lane12_strm1_data          ( std__pe7__lane12_strm1_data       ),      
               .std__pe7__lane12_strm1_data_valid    ( std__pe7__lane12_strm1_data_valid ),      
               .std__pe7__lane12_strm1_data_mask     ( std__pe7__lane12_strm1_data_mask  ),      

               // PE 7, Lane 13                 
               .pe7__std__lane13_strm0_ready         ( pe7__std__lane13_strm0_ready      ),      
               .std__pe7__lane13_strm0_cntl          ( std__pe7__lane13_strm0_cntl       ),      
               .std__pe7__lane13_strm0_data          ( std__pe7__lane13_strm0_data       ),      
               .std__pe7__lane13_strm0_data_valid    ( std__pe7__lane13_strm0_data_valid ),      
               .std__pe7__lane13_strm0_data_mask     ( std__pe7__lane13_strm0_data_mask  ),      

               .pe7__std__lane13_strm1_ready         ( pe7__std__lane13_strm1_ready      ),      
               .std__pe7__lane13_strm1_cntl          ( std__pe7__lane13_strm1_cntl       ),      
               .std__pe7__lane13_strm1_data          ( std__pe7__lane13_strm1_data       ),      
               .std__pe7__lane13_strm1_data_valid    ( std__pe7__lane13_strm1_data_valid ),      
               .std__pe7__lane13_strm1_data_mask     ( std__pe7__lane13_strm1_data_mask  ),      

               // PE 7, Lane 14                 
               .pe7__std__lane14_strm0_ready         ( pe7__std__lane14_strm0_ready      ),      
               .std__pe7__lane14_strm0_cntl          ( std__pe7__lane14_strm0_cntl       ),      
               .std__pe7__lane14_strm0_data          ( std__pe7__lane14_strm0_data       ),      
               .std__pe7__lane14_strm0_data_valid    ( std__pe7__lane14_strm0_data_valid ),      
               .std__pe7__lane14_strm0_data_mask     ( std__pe7__lane14_strm0_data_mask  ),      

               .pe7__std__lane14_strm1_ready         ( pe7__std__lane14_strm1_ready      ),      
               .std__pe7__lane14_strm1_cntl          ( std__pe7__lane14_strm1_cntl       ),      
               .std__pe7__lane14_strm1_data          ( std__pe7__lane14_strm1_data       ),      
               .std__pe7__lane14_strm1_data_valid    ( std__pe7__lane14_strm1_data_valid ),      
               .std__pe7__lane14_strm1_data_mask     ( std__pe7__lane14_strm1_data_mask  ),      

               // PE 7, Lane 15                 
               .pe7__std__lane15_strm0_ready         ( pe7__std__lane15_strm0_ready      ),      
               .std__pe7__lane15_strm0_cntl          ( std__pe7__lane15_strm0_cntl       ),      
               .std__pe7__lane15_strm0_data          ( std__pe7__lane15_strm0_data       ),      
               .std__pe7__lane15_strm0_data_valid    ( std__pe7__lane15_strm0_data_valid ),      
               .std__pe7__lane15_strm0_data_mask     ( std__pe7__lane15_strm0_data_mask  ),      

               .pe7__std__lane15_strm1_ready         ( pe7__std__lane15_strm1_ready      ),      
               .std__pe7__lane15_strm1_cntl          ( std__pe7__lane15_strm1_cntl       ),      
               .std__pe7__lane15_strm1_data          ( std__pe7__lane15_strm1_data       ),      
               .std__pe7__lane15_strm1_data_valid    ( std__pe7__lane15_strm1_data_valid ),      
               .std__pe7__lane15_strm1_data_mask     ( std__pe7__lane15_strm1_data_mask  ),      

               // PE 7, Lane 16                 
               .pe7__std__lane16_strm0_ready         ( pe7__std__lane16_strm0_ready      ),      
               .std__pe7__lane16_strm0_cntl          ( std__pe7__lane16_strm0_cntl       ),      
               .std__pe7__lane16_strm0_data          ( std__pe7__lane16_strm0_data       ),      
               .std__pe7__lane16_strm0_data_valid    ( std__pe7__lane16_strm0_data_valid ),      
               .std__pe7__lane16_strm0_data_mask     ( std__pe7__lane16_strm0_data_mask  ),      

               .pe7__std__lane16_strm1_ready         ( pe7__std__lane16_strm1_ready      ),      
               .std__pe7__lane16_strm1_cntl          ( std__pe7__lane16_strm1_cntl       ),      
               .std__pe7__lane16_strm1_data          ( std__pe7__lane16_strm1_data       ),      
               .std__pe7__lane16_strm1_data_valid    ( std__pe7__lane16_strm1_data_valid ),      
               .std__pe7__lane16_strm1_data_mask     ( std__pe7__lane16_strm1_data_mask  ),      

               // PE 7, Lane 17                 
               .pe7__std__lane17_strm0_ready         ( pe7__std__lane17_strm0_ready      ),      
               .std__pe7__lane17_strm0_cntl          ( std__pe7__lane17_strm0_cntl       ),      
               .std__pe7__lane17_strm0_data          ( std__pe7__lane17_strm0_data       ),      
               .std__pe7__lane17_strm0_data_valid    ( std__pe7__lane17_strm0_data_valid ),      
               .std__pe7__lane17_strm0_data_mask     ( std__pe7__lane17_strm0_data_mask  ),      

               .pe7__std__lane17_strm1_ready         ( pe7__std__lane17_strm1_ready      ),      
               .std__pe7__lane17_strm1_cntl          ( std__pe7__lane17_strm1_cntl       ),      
               .std__pe7__lane17_strm1_data          ( std__pe7__lane17_strm1_data       ),      
               .std__pe7__lane17_strm1_data_valid    ( std__pe7__lane17_strm1_data_valid ),      
               .std__pe7__lane17_strm1_data_mask     ( std__pe7__lane17_strm1_data_mask  ),      

               // PE 7, Lane 18                 
               .pe7__std__lane18_strm0_ready         ( pe7__std__lane18_strm0_ready      ),      
               .std__pe7__lane18_strm0_cntl          ( std__pe7__lane18_strm0_cntl       ),      
               .std__pe7__lane18_strm0_data          ( std__pe7__lane18_strm0_data       ),      
               .std__pe7__lane18_strm0_data_valid    ( std__pe7__lane18_strm0_data_valid ),      
               .std__pe7__lane18_strm0_data_mask     ( std__pe7__lane18_strm0_data_mask  ),      

               .pe7__std__lane18_strm1_ready         ( pe7__std__lane18_strm1_ready      ),      
               .std__pe7__lane18_strm1_cntl          ( std__pe7__lane18_strm1_cntl       ),      
               .std__pe7__lane18_strm1_data          ( std__pe7__lane18_strm1_data       ),      
               .std__pe7__lane18_strm1_data_valid    ( std__pe7__lane18_strm1_data_valid ),      
               .std__pe7__lane18_strm1_data_mask     ( std__pe7__lane18_strm1_data_mask  ),      

               // PE 7, Lane 19                 
               .pe7__std__lane19_strm0_ready         ( pe7__std__lane19_strm0_ready      ),      
               .std__pe7__lane19_strm0_cntl          ( std__pe7__lane19_strm0_cntl       ),      
               .std__pe7__lane19_strm0_data          ( std__pe7__lane19_strm0_data       ),      
               .std__pe7__lane19_strm0_data_valid    ( std__pe7__lane19_strm0_data_valid ),      
               .std__pe7__lane19_strm0_data_mask     ( std__pe7__lane19_strm0_data_mask  ),      

               .pe7__std__lane19_strm1_ready         ( pe7__std__lane19_strm1_ready      ),      
               .std__pe7__lane19_strm1_cntl          ( std__pe7__lane19_strm1_cntl       ),      
               .std__pe7__lane19_strm1_data          ( std__pe7__lane19_strm1_data       ),      
               .std__pe7__lane19_strm1_data_valid    ( std__pe7__lane19_strm1_data_valid ),      
               .std__pe7__lane19_strm1_data_mask     ( std__pe7__lane19_strm1_data_mask  ),      

               // PE 7, Lane 20                 
               .pe7__std__lane20_strm0_ready         ( pe7__std__lane20_strm0_ready      ),      
               .std__pe7__lane20_strm0_cntl          ( std__pe7__lane20_strm0_cntl       ),      
               .std__pe7__lane20_strm0_data          ( std__pe7__lane20_strm0_data       ),      
               .std__pe7__lane20_strm0_data_valid    ( std__pe7__lane20_strm0_data_valid ),      
               .std__pe7__lane20_strm0_data_mask     ( std__pe7__lane20_strm0_data_mask  ),      

               .pe7__std__lane20_strm1_ready         ( pe7__std__lane20_strm1_ready      ),      
               .std__pe7__lane20_strm1_cntl          ( std__pe7__lane20_strm1_cntl       ),      
               .std__pe7__lane20_strm1_data          ( std__pe7__lane20_strm1_data       ),      
               .std__pe7__lane20_strm1_data_valid    ( std__pe7__lane20_strm1_data_valid ),      
               .std__pe7__lane20_strm1_data_mask     ( std__pe7__lane20_strm1_data_mask  ),      

               // PE 7, Lane 21                 
               .pe7__std__lane21_strm0_ready         ( pe7__std__lane21_strm0_ready      ),      
               .std__pe7__lane21_strm0_cntl          ( std__pe7__lane21_strm0_cntl       ),      
               .std__pe7__lane21_strm0_data          ( std__pe7__lane21_strm0_data       ),      
               .std__pe7__lane21_strm0_data_valid    ( std__pe7__lane21_strm0_data_valid ),      
               .std__pe7__lane21_strm0_data_mask     ( std__pe7__lane21_strm0_data_mask  ),      

               .pe7__std__lane21_strm1_ready         ( pe7__std__lane21_strm1_ready      ),      
               .std__pe7__lane21_strm1_cntl          ( std__pe7__lane21_strm1_cntl       ),      
               .std__pe7__lane21_strm1_data          ( std__pe7__lane21_strm1_data       ),      
               .std__pe7__lane21_strm1_data_valid    ( std__pe7__lane21_strm1_data_valid ),      
               .std__pe7__lane21_strm1_data_mask     ( std__pe7__lane21_strm1_data_mask  ),      

               // PE 7, Lane 22                 
               .pe7__std__lane22_strm0_ready         ( pe7__std__lane22_strm0_ready      ),      
               .std__pe7__lane22_strm0_cntl          ( std__pe7__lane22_strm0_cntl       ),      
               .std__pe7__lane22_strm0_data          ( std__pe7__lane22_strm0_data       ),      
               .std__pe7__lane22_strm0_data_valid    ( std__pe7__lane22_strm0_data_valid ),      
               .std__pe7__lane22_strm0_data_mask     ( std__pe7__lane22_strm0_data_mask  ),      

               .pe7__std__lane22_strm1_ready         ( pe7__std__lane22_strm1_ready      ),      
               .std__pe7__lane22_strm1_cntl          ( std__pe7__lane22_strm1_cntl       ),      
               .std__pe7__lane22_strm1_data          ( std__pe7__lane22_strm1_data       ),      
               .std__pe7__lane22_strm1_data_valid    ( std__pe7__lane22_strm1_data_valid ),      
               .std__pe7__lane22_strm1_data_mask     ( std__pe7__lane22_strm1_data_mask  ),      

               // PE 7, Lane 23                 
               .pe7__std__lane23_strm0_ready         ( pe7__std__lane23_strm0_ready      ),      
               .std__pe7__lane23_strm0_cntl          ( std__pe7__lane23_strm0_cntl       ),      
               .std__pe7__lane23_strm0_data          ( std__pe7__lane23_strm0_data       ),      
               .std__pe7__lane23_strm0_data_valid    ( std__pe7__lane23_strm0_data_valid ),      
               .std__pe7__lane23_strm0_data_mask     ( std__pe7__lane23_strm0_data_mask  ),      

               .pe7__std__lane23_strm1_ready         ( pe7__std__lane23_strm1_ready      ),      
               .std__pe7__lane23_strm1_cntl          ( std__pe7__lane23_strm1_cntl       ),      
               .std__pe7__lane23_strm1_data          ( std__pe7__lane23_strm1_data       ),      
               .std__pe7__lane23_strm1_data_valid    ( std__pe7__lane23_strm1_data_valid ),      
               .std__pe7__lane23_strm1_data_mask     ( std__pe7__lane23_strm1_data_mask  ),      

               // PE 7, Lane 24                 
               .pe7__std__lane24_strm0_ready         ( pe7__std__lane24_strm0_ready      ),      
               .std__pe7__lane24_strm0_cntl          ( std__pe7__lane24_strm0_cntl       ),      
               .std__pe7__lane24_strm0_data          ( std__pe7__lane24_strm0_data       ),      
               .std__pe7__lane24_strm0_data_valid    ( std__pe7__lane24_strm0_data_valid ),      
               .std__pe7__lane24_strm0_data_mask     ( std__pe7__lane24_strm0_data_mask  ),      

               .pe7__std__lane24_strm1_ready         ( pe7__std__lane24_strm1_ready      ),      
               .std__pe7__lane24_strm1_cntl          ( std__pe7__lane24_strm1_cntl       ),      
               .std__pe7__lane24_strm1_data          ( std__pe7__lane24_strm1_data       ),      
               .std__pe7__lane24_strm1_data_valid    ( std__pe7__lane24_strm1_data_valid ),      
               .std__pe7__lane24_strm1_data_mask     ( std__pe7__lane24_strm1_data_mask  ),      

               // PE 7, Lane 25                 
               .pe7__std__lane25_strm0_ready         ( pe7__std__lane25_strm0_ready      ),      
               .std__pe7__lane25_strm0_cntl          ( std__pe7__lane25_strm0_cntl       ),      
               .std__pe7__lane25_strm0_data          ( std__pe7__lane25_strm0_data       ),      
               .std__pe7__lane25_strm0_data_valid    ( std__pe7__lane25_strm0_data_valid ),      
               .std__pe7__lane25_strm0_data_mask     ( std__pe7__lane25_strm0_data_mask  ),      

               .pe7__std__lane25_strm1_ready         ( pe7__std__lane25_strm1_ready      ),      
               .std__pe7__lane25_strm1_cntl          ( std__pe7__lane25_strm1_cntl       ),      
               .std__pe7__lane25_strm1_data          ( std__pe7__lane25_strm1_data       ),      
               .std__pe7__lane25_strm1_data_valid    ( std__pe7__lane25_strm1_data_valid ),      
               .std__pe7__lane25_strm1_data_mask     ( std__pe7__lane25_strm1_data_mask  ),      

               // PE 7, Lane 26                 
               .pe7__std__lane26_strm0_ready         ( pe7__std__lane26_strm0_ready      ),      
               .std__pe7__lane26_strm0_cntl          ( std__pe7__lane26_strm0_cntl       ),      
               .std__pe7__lane26_strm0_data          ( std__pe7__lane26_strm0_data       ),      
               .std__pe7__lane26_strm0_data_valid    ( std__pe7__lane26_strm0_data_valid ),      
               .std__pe7__lane26_strm0_data_mask     ( std__pe7__lane26_strm0_data_mask  ),      

               .pe7__std__lane26_strm1_ready         ( pe7__std__lane26_strm1_ready      ),      
               .std__pe7__lane26_strm1_cntl          ( std__pe7__lane26_strm1_cntl       ),      
               .std__pe7__lane26_strm1_data          ( std__pe7__lane26_strm1_data       ),      
               .std__pe7__lane26_strm1_data_valid    ( std__pe7__lane26_strm1_data_valid ),      
               .std__pe7__lane26_strm1_data_mask     ( std__pe7__lane26_strm1_data_mask  ),      

               // PE 7, Lane 27                 
               .pe7__std__lane27_strm0_ready         ( pe7__std__lane27_strm0_ready      ),      
               .std__pe7__lane27_strm0_cntl          ( std__pe7__lane27_strm0_cntl       ),      
               .std__pe7__lane27_strm0_data          ( std__pe7__lane27_strm0_data       ),      
               .std__pe7__lane27_strm0_data_valid    ( std__pe7__lane27_strm0_data_valid ),      
               .std__pe7__lane27_strm0_data_mask     ( std__pe7__lane27_strm0_data_mask  ),      

               .pe7__std__lane27_strm1_ready         ( pe7__std__lane27_strm1_ready      ),      
               .std__pe7__lane27_strm1_cntl          ( std__pe7__lane27_strm1_cntl       ),      
               .std__pe7__lane27_strm1_data          ( std__pe7__lane27_strm1_data       ),      
               .std__pe7__lane27_strm1_data_valid    ( std__pe7__lane27_strm1_data_valid ),      
               .std__pe7__lane27_strm1_data_mask     ( std__pe7__lane27_strm1_data_mask  ),      

               // PE 7, Lane 28                 
               .pe7__std__lane28_strm0_ready         ( pe7__std__lane28_strm0_ready      ),      
               .std__pe7__lane28_strm0_cntl          ( std__pe7__lane28_strm0_cntl       ),      
               .std__pe7__lane28_strm0_data          ( std__pe7__lane28_strm0_data       ),      
               .std__pe7__lane28_strm0_data_valid    ( std__pe7__lane28_strm0_data_valid ),      
               .std__pe7__lane28_strm0_data_mask     ( std__pe7__lane28_strm0_data_mask  ),      

               .pe7__std__lane28_strm1_ready         ( pe7__std__lane28_strm1_ready      ),      
               .std__pe7__lane28_strm1_cntl          ( std__pe7__lane28_strm1_cntl       ),      
               .std__pe7__lane28_strm1_data          ( std__pe7__lane28_strm1_data       ),      
               .std__pe7__lane28_strm1_data_valid    ( std__pe7__lane28_strm1_data_valid ),      
               .std__pe7__lane28_strm1_data_mask     ( std__pe7__lane28_strm1_data_mask  ),      

               // PE 7, Lane 29                 
               .pe7__std__lane29_strm0_ready         ( pe7__std__lane29_strm0_ready      ),      
               .std__pe7__lane29_strm0_cntl          ( std__pe7__lane29_strm0_cntl       ),      
               .std__pe7__lane29_strm0_data          ( std__pe7__lane29_strm0_data       ),      
               .std__pe7__lane29_strm0_data_valid    ( std__pe7__lane29_strm0_data_valid ),      
               .std__pe7__lane29_strm0_data_mask     ( std__pe7__lane29_strm0_data_mask  ),      

               .pe7__std__lane29_strm1_ready         ( pe7__std__lane29_strm1_ready      ),      
               .std__pe7__lane29_strm1_cntl          ( std__pe7__lane29_strm1_cntl       ),      
               .std__pe7__lane29_strm1_data          ( std__pe7__lane29_strm1_data       ),      
               .std__pe7__lane29_strm1_data_valid    ( std__pe7__lane29_strm1_data_valid ),      
               .std__pe7__lane29_strm1_data_mask     ( std__pe7__lane29_strm1_data_mask  ),      

               // PE 7, Lane 30                 
               .pe7__std__lane30_strm0_ready         ( pe7__std__lane30_strm0_ready      ),      
               .std__pe7__lane30_strm0_cntl          ( std__pe7__lane30_strm0_cntl       ),      
               .std__pe7__lane30_strm0_data          ( std__pe7__lane30_strm0_data       ),      
               .std__pe7__lane30_strm0_data_valid    ( std__pe7__lane30_strm0_data_valid ),      
               .std__pe7__lane30_strm0_data_mask     ( std__pe7__lane30_strm0_data_mask  ),      

               .pe7__std__lane30_strm1_ready         ( pe7__std__lane30_strm1_ready      ),      
               .std__pe7__lane30_strm1_cntl          ( std__pe7__lane30_strm1_cntl       ),      
               .std__pe7__lane30_strm1_data          ( std__pe7__lane30_strm1_data       ),      
               .std__pe7__lane30_strm1_data_valid    ( std__pe7__lane30_strm1_data_valid ),      
               .std__pe7__lane30_strm1_data_mask     ( std__pe7__lane30_strm1_data_mask  ),      

               // PE 7, Lane 31                 
               .pe7__std__lane31_strm0_ready         ( pe7__std__lane31_strm0_ready      ),      
               .std__pe7__lane31_strm0_cntl          ( std__pe7__lane31_strm0_cntl       ),      
               .std__pe7__lane31_strm0_data          ( std__pe7__lane31_strm0_data       ),      
               .std__pe7__lane31_strm0_data_valid    ( std__pe7__lane31_strm0_data_valid ),      
               .std__pe7__lane31_strm0_data_mask     ( std__pe7__lane31_strm0_data_mask  ),      

               .pe7__std__lane31_strm1_ready         ( pe7__std__lane31_strm1_ready      ),      
               .std__pe7__lane31_strm1_cntl          ( std__pe7__lane31_strm1_cntl       ),      
               .std__pe7__lane31_strm1_data          ( std__pe7__lane31_strm1_data       ),      
               .std__pe7__lane31_strm1_data_valid    ( std__pe7__lane31_strm1_data_valid ),      
               .std__pe7__lane31_strm1_data_mask     ( std__pe7__lane31_strm1_data_mask  ),      

               // PE 8, Lane 0                 
               .pe8__std__lane0_strm0_ready         ( pe8__std__lane0_strm0_ready      ),      
               .std__pe8__lane0_strm0_cntl          ( std__pe8__lane0_strm0_cntl       ),      
               .std__pe8__lane0_strm0_data          ( std__pe8__lane0_strm0_data       ),      
               .std__pe8__lane0_strm0_data_valid    ( std__pe8__lane0_strm0_data_valid ),      
               .std__pe8__lane0_strm0_data_mask     ( std__pe8__lane0_strm0_data_mask  ),      

               .pe8__std__lane0_strm1_ready         ( pe8__std__lane0_strm1_ready      ),      
               .std__pe8__lane0_strm1_cntl          ( std__pe8__lane0_strm1_cntl       ),      
               .std__pe8__lane0_strm1_data          ( std__pe8__lane0_strm1_data       ),      
               .std__pe8__lane0_strm1_data_valid    ( std__pe8__lane0_strm1_data_valid ),      
               .std__pe8__lane0_strm1_data_mask     ( std__pe8__lane0_strm1_data_mask  ),      

               // PE 8, Lane 1                 
               .pe8__std__lane1_strm0_ready         ( pe8__std__lane1_strm0_ready      ),      
               .std__pe8__lane1_strm0_cntl          ( std__pe8__lane1_strm0_cntl       ),      
               .std__pe8__lane1_strm0_data          ( std__pe8__lane1_strm0_data       ),      
               .std__pe8__lane1_strm0_data_valid    ( std__pe8__lane1_strm0_data_valid ),      
               .std__pe8__lane1_strm0_data_mask     ( std__pe8__lane1_strm0_data_mask  ),      

               .pe8__std__lane1_strm1_ready         ( pe8__std__lane1_strm1_ready      ),      
               .std__pe8__lane1_strm1_cntl          ( std__pe8__lane1_strm1_cntl       ),      
               .std__pe8__lane1_strm1_data          ( std__pe8__lane1_strm1_data       ),      
               .std__pe8__lane1_strm1_data_valid    ( std__pe8__lane1_strm1_data_valid ),      
               .std__pe8__lane1_strm1_data_mask     ( std__pe8__lane1_strm1_data_mask  ),      

               // PE 8, Lane 2                 
               .pe8__std__lane2_strm0_ready         ( pe8__std__lane2_strm0_ready      ),      
               .std__pe8__lane2_strm0_cntl          ( std__pe8__lane2_strm0_cntl       ),      
               .std__pe8__lane2_strm0_data          ( std__pe8__lane2_strm0_data       ),      
               .std__pe8__lane2_strm0_data_valid    ( std__pe8__lane2_strm0_data_valid ),      
               .std__pe8__lane2_strm0_data_mask     ( std__pe8__lane2_strm0_data_mask  ),      

               .pe8__std__lane2_strm1_ready         ( pe8__std__lane2_strm1_ready      ),      
               .std__pe8__lane2_strm1_cntl          ( std__pe8__lane2_strm1_cntl       ),      
               .std__pe8__lane2_strm1_data          ( std__pe8__lane2_strm1_data       ),      
               .std__pe8__lane2_strm1_data_valid    ( std__pe8__lane2_strm1_data_valid ),      
               .std__pe8__lane2_strm1_data_mask     ( std__pe8__lane2_strm1_data_mask  ),      

               // PE 8, Lane 3                 
               .pe8__std__lane3_strm0_ready         ( pe8__std__lane3_strm0_ready      ),      
               .std__pe8__lane3_strm0_cntl          ( std__pe8__lane3_strm0_cntl       ),      
               .std__pe8__lane3_strm0_data          ( std__pe8__lane3_strm0_data       ),      
               .std__pe8__lane3_strm0_data_valid    ( std__pe8__lane3_strm0_data_valid ),      
               .std__pe8__lane3_strm0_data_mask     ( std__pe8__lane3_strm0_data_mask  ),      

               .pe8__std__lane3_strm1_ready         ( pe8__std__lane3_strm1_ready      ),      
               .std__pe8__lane3_strm1_cntl          ( std__pe8__lane3_strm1_cntl       ),      
               .std__pe8__lane3_strm1_data          ( std__pe8__lane3_strm1_data       ),      
               .std__pe8__lane3_strm1_data_valid    ( std__pe8__lane3_strm1_data_valid ),      
               .std__pe8__lane3_strm1_data_mask     ( std__pe8__lane3_strm1_data_mask  ),      

               // PE 8, Lane 4                 
               .pe8__std__lane4_strm0_ready         ( pe8__std__lane4_strm0_ready      ),      
               .std__pe8__lane4_strm0_cntl          ( std__pe8__lane4_strm0_cntl       ),      
               .std__pe8__lane4_strm0_data          ( std__pe8__lane4_strm0_data       ),      
               .std__pe8__lane4_strm0_data_valid    ( std__pe8__lane4_strm0_data_valid ),      
               .std__pe8__lane4_strm0_data_mask     ( std__pe8__lane4_strm0_data_mask  ),      

               .pe8__std__lane4_strm1_ready         ( pe8__std__lane4_strm1_ready      ),      
               .std__pe8__lane4_strm1_cntl          ( std__pe8__lane4_strm1_cntl       ),      
               .std__pe8__lane4_strm1_data          ( std__pe8__lane4_strm1_data       ),      
               .std__pe8__lane4_strm1_data_valid    ( std__pe8__lane4_strm1_data_valid ),      
               .std__pe8__lane4_strm1_data_mask     ( std__pe8__lane4_strm1_data_mask  ),      

               // PE 8, Lane 5                 
               .pe8__std__lane5_strm0_ready         ( pe8__std__lane5_strm0_ready      ),      
               .std__pe8__lane5_strm0_cntl          ( std__pe8__lane5_strm0_cntl       ),      
               .std__pe8__lane5_strm0_data          ( std__pe8__lane5_strm0_data       ),      
               .std__pe8__lane5_strm0_data_valid    ( std__pe8__lane5_strm0_data_valid ),      
               .std__pe8__lane5_strm0_data_mask     ( std__pe8__lane5_strm0_data_mask  ),      

               .pe8__std__lane5_strm1_ready         ( pe8__std__lane5_strm1_ready      ),      
               .std__pe8__lane5_strm1_cntl          ( std__pe8__lane5_strm1_cntl       ),      
               .std__pe8__lane5_strm1_data          ( std__pe8__lane5_strm1_data       ),      
               .std__pe8__lane5_strm1_data_valid    ( std__pe8__lane5_strm1_data_valid ),      
               .std__pe8__lane5_strm1_data_mask     ( std__pe8__lane5_strm1_data_mask  ),      

               // PE 8, Lane 6                 
               .pe8__std__lane6_strm0_ready         ( pe8__std__lane6_strm0_ready      ),      
               .std__pe8__lane6_strm0_cntl          ( std__pe8__lane6_strm0_cntl       ),      
               .std__pe8__lane6_strm0_data          ( std__pe8__lane6_strm0_data       ),      
               .std__pe8__lane6_strm0_data_valid    ( std__pe8__lane6_strm0_data_valid ),      
               .std__pe8__lane6_strm0_data_mask     ( std__pe8__lane6_strm0_data_mask  ),      

               .pe8__std__lane6_strm1_ready         ( pe8__std__lane6_strm1_ready      ),      
               .std__pe8__lane6_strm1_cntl          ( std__pe8__lane6_strm1_cntl       ),      
               .std__pe8__lane6_strm1_data          ( std__pe8__lane6_strm1_data       ),      
               .std__pe8__lane6_strm1_data_valid    ( std__pe8__lane6_strm1_data_valid ),      
               .std__pe8__lane6_strm1_data_mask     ( std__pe8__lane6_strm1_data_mask  ),      

               // PE 8, Lane 7                 
               .pe8__std__lane7_strm0_ready         ( pe8__std__lane7_strm0_ready      ),      
               .std__pe8__lane7_strm0_cntl          ( std__pe8__lane7_strm0_cntl       ),      
               .std__pe8__lane7_strm0_data          ( std__pe8__lane7_strm0_data       ),      
               .std__pe8__lane7_strm0_data_valid    ( std__pe8__lane7_strm0_data_valid ),      
               .std__pe8__lane7_strm0_data_mask     ( std__pe8__lane7_strm0_data_mask  ),      

               .pe8__std__lane7_strm1_ready         ( pe8__std__lane7_strm1_ready      ),      
               .std__pe8__lane7_strm1_cntl          ( std__pe8__lane7_strm1_cntl       ),      
               .std__pe8__lane7_strm1_data          ( std__pe8__lane7_strm1_data       ),      
               .std__pe8__lane7_strm1_data_valid    ( std__pe8__lane7_strm1_data_valid ),      
               .std__pe8__lane7_strm1_data_mask     ( std__pe8__lane7_strm1_data_mask  ),      

               // PE 8, Lane 8                 
               .pe8__std__lane8_strm0_ready         ( pe8__std__lane8_strm0_ready      ),      
               .std__pe8__lane8_strm0_cntl          ( std__pe8__lane8_strm0_cntl       ),      
               .std__pe8__lane8_strm0_data          ( std__pe8__lane8_strm0_data       ),      
               .std__pe8__lane8_strm0_data_valid    ( std__pe8__lane8_strm0_data_valid ),      
               .std__pe8__lane8_strm0_data_mask     ( std__pe8__lane8_strm0_data_mask  ),      

               .pe8__std__lane8_strm1_ready         ( pe8__std__lane8_strm1_ready      ),      
               .std__pe8__lane8_strm1_cntl          ( std__pe8__lane8_strm1_cntl       ),      
               .std__pe8__lane8_strm1_data          ( std__pe8__lane8_strm1_data       ),      
               .std__pe8__lane8_strm1_data_valid    ( std__pe8__lane8_strm1_data_valid ),      
               .std__pe8__lane8_strm1_data_mask     ( std__pe8__lane8_strm1_data_mask  ),      

               // PE 8, Lane 9                 
               .pe8__std__lane9_strm0_ready         ( pe8__std__lane9_strm0_ready      ),      
               .std__pe8__lane9_strm0_cntl          ( std__pe8__lane9_strm0_cntl       ),      
               .std__pe8__lane9_strm0_data          ( std__pe8__lane9_strm0_data       ),      
               .std__pe8__lane9_strm0_data_valid    ( std__pe8__lane9_strm0_data_valid ),      
               .std__pe8__lane9_strm0_data_mask     ( std__pe8__lane9_strm0_data_mask  ),      

               .pe8__std__lane9_strm1_ready         ( pe8__std__lane9_strm1_ready      ),      
               .std__pe8__lane9_strm1_cntl          ( std__pe8__lane9_strm1_cntl       ),      
               .std__pe8__lane9_strm1_data          ( std__pe8__lane9_strm1_data       ),      
               .std__pe8__lane9_strm1_data_valid    ( std__pe8__lane9_strm1_data_valid ),      
               .std__pe8__lane9_strm1_data_mask     ( std__pe8__lane9_strm1_data_mask  ),      

               // PE 8, Lane 10                 
               .pe8__std__lane10_strm0_ready         ( pe8__std__lane10_strm0_ready      ),      
               .std__pe8__lane10_strm0_cntl          ( std__pe8__lane10_strm0_cntl       ),      
               .std__pe8__lane10_strm0_data          ( std__pe8__lane10_strm0_data       ),      
               .std__pe8__lane10_strm0_data_valid    ( std__pe8__lane10_strm0_data_valid ),      
               .std__pe8__lane10_strm0_data_mask     ( std__pe8__lane10_strm0_data_mask  ),      

               .pe8__std__lane10_strm1_ready         ( pe8__std__lane10_strm1_ready      ),      
               .std__pe8__lane10_strm1_cntl          ( std__pe8__lane10_strm1_cntl       ),      
               .std__pe8__lane10_strm1_data          ( std__pe8__lane10_strm1_data       ),      
               .std__pe8__lane10_strm1_data_valid    ( std__pe8__lane10_strm1_data_valid ),      
               .std__pe8__lane10_strm1_data_mask     ( std__pe8__lane10_strm1_data_mask  ),      

               // PE 8, Lane 11                 
               .pe8__std__lane11_strm0_ready         ( pe8__std__lane11_strm0_ready      ),      
               .std__pe8__lane11_strm0_cntl          ( std__pe8__lane11_strm0_cntl       ),      
               .std__pe8__lane11_strm0_data          ( std__pe8__lane11_strm0_data       ),      
               .std__pe8__lane11_strm0_data_valid    ( std__pe8__lane11_strm0_data_valid ),      
               .std__pe8__lane11_strm0_data_mask     ( std__pe8__lane11_strm0_data_mask  ),      

               .pe8__std__lane11_strm1_ready         ( pe8__std__lane11_strm1_ready      ),      
               .std__pe8__lane11_strm1_cntl          ( std__pe8__lane11_strm1_cntl       ),      
               .std__pe8__lane11_strm1_data          ( std__pe8__lane11_strm1_data       ),      
               .std__pe8__lane11_strm1_data_valid    ( std__pe8__lane11_strm1_data_valid ),      
               .std__pe8__lane11_strm1_data_mask     ( std__pe8__lane11_strm1_data_mask  ),      

               // PE 8, Lane 12                 
               .pe8__std__lane12_strm0_ready         ( pe8__std__lane12_strm0_ready      ),      
               .std__pe8__lane12_strm0_cntl          ( std__pe8__lane12_strm0_cntl       ),      
               .std__pe8__lane12_strm0_data          ( std__pe8__lane12_strm0_data       ),      
               .std__pe8__lane12_strm0_data_valid    ( std__pe8__lane12_strm0_data_valid ),      
               .std__pe8__lane12_strm0_data_mask     ( std__pe8__lane12_strm0_data_mask  ),      

               .pe8__std__lane12_strm1_ready         ( pe8__std__lane12_strm1_ready      ),      
               .std__pe8__lane12_strm1_cntl          ( std__pe8__lane12_strm1_cntl       ),      
               .std__pe8__lane12_strm1_data          ( std__pe8__lane12_strm1_data       ),      
               .std__pe8__lane12_strm1_data_valid    ( std__pe8__lane12_strm1_data_valid ),      
               .std__pe8__lane12_strm1_data_mask     ( std__pe8__lane12_strm1_data_mask  ),      

               // PE 8, Lane 13                 
               .pe8__std__lane13_strm0_ready         ( pe8__std__lane13_strm0_ready      ),      
               .std__pe8__lane13_strm0_cntl          ( std__pe8__lane13_strm0_cntl       ),      
               .std__pe8__lane13_strm0_data          ( std__pe8__lane13_strm0_data       ),      
               .std__pe8__lane13_strm0_data_valid    ( std__pe8__lane13_strm0_data_valid ),      
               .std__pe8__lane13_strm0_data_mask     ( std__pe8__lane13_strm0_data_mask  ),      

               .pe8__std__lane13_strm1_ready         ( pe8__std__lane13_strm1_ready      ),      
               .std__pe8__lane13_strm1_cntl          ( std__pe8__lane13_strm1_cntl       ),      
               .std__pe8__lane13_strm1_data          ( std__pe8__lane13_strm1_data       ),      
               .std__pe8__lane13_strm1_data_valid    ( std__pe8__lane13_strm1_data_valid ),      
               .std__pe8__lane13_strm1_data_mask     ( std__pe8__lane13_strm1_data_mask  ),      

               // PE 8, Lane 14                 
               .pe8__std__lane14_strm0_ready         ( pe8__std__lane14_strm0_ready      ),      
               .std__pe8__lane14_strm0_cntl          ( std__pe8__lane14_strm0_cntl       ),      
               .std__pe8__lane14_strm0_data          ( std__pe8__lane14_strm0_data       ),      
               .std__pe8__lane14_strm0_data_valid    ( std__pe8__lane14_strm0_data_valid ),      
               .std__pe8__lane14_strm0_data_mask     ( std__pe8__lane14_strm0_data_mask  ),      

               .pe8__std__lane14_strm1_ready         ( pe8__std__lane14_strm1_ready      ),      
               .std__pe8__lane14_strm1_cntl          ( std__pe8__lane14_strm1_cntl       ),      
               .std__pe8__lane14_strm1_data          ( std__pe8__lane14_strm1_data       ),      
               .std__pe8__lane14_strm1_data_valid    ( std__pe8__lane14_strm1_data_valid ),      
               .std__pe8__lane14_strm1_data_mask     ( std__pe8__lane14_strm1_data_mask  ),      

               // PE 8, Lane 15                 
               .pe8__std__lane15_strm0_ready         ( pe8__std__lane15_strm0_ready      ),      
               .std__pe8__lane15_strm0_cntl          ( std__pe8__lane15_strm0_cntl       ),      
               .std__pe8__lane15_strm0_data          ( std__pe8__lane15_strm0_data       ),      
               .std__pe8__lane15_strm0_data_valid    ( std__pe8__lane15_strm0_data_valid ),      
               .std__pe8__lane15_strm0_data_mask     ( std__pe8__lane15_strm0_data_mask  ),      

               .pe8__std__lane15_strm1_ready         ( pe8__std__lane15_strm1_ready      ),      
               .std__pe8__lane15_strm1_cntl          ( std__pe8__lane15_strm1_cntl       ),      
               .std__pe8__lane15_strm1_data          ( std__pe8__lane15_strm1_data       ),      
               .std__pe8__lane15_strm1_data_valid    ( std__pe8__lane15_strm1_data_valid ),      
               .std__pe8__lane15_strm1_data_mask     ( std__pe8__lane15_strm1_data_mask  ),      

               // PE 8, Lane 16                 
               .pe8__std__lane16_strm0_ready         ( pe8__std__lane16_strm0_ready      ),      
               .std__pe8__lane16_strm0_cntl          ( std__pe8__lane16_strm0_cntl       ),      
               .std__pe8__lane16_strm0_data          ( std__pe8__lane16_strm0_data       ),      
               .std__pe8__lane16_strm0_data_valid    ( std__pe8__lane16_strm0_data_valid ),      
               .std__pe8__lane16_strm0_data_mask     ( std__pe8__lane16_strm0_data_mask  ),      

               .pe8__std__lane16_strm1_ready         ( pe8__std__lane16_strm1_ready      ),      
               .std__pe8__lane16_strm1_cntl          ( std__pe8__lane16_strm1_cntl       ),      
               .std__pe8__lane16_strm1_data          ( std__pe8__lane16_strm1_data       ),      
               .std__pe8__lane16_strm1_data_valid    ( std__pe8__lane16_strm1_data_valid ),      
               .std__pe8__lane16_strm1_data_mask     ( std__pe8__lane16_strm1_data_mask  ),      

               // PE 8, Lane 17                 
               .pe8__std__lane17_strm0_ready         ( pe8__std__lane17_strm0_ready      ),      
               .std__pe8__lane17_strm0_cntl          ( std__pe8__lane17_strm0_cntl       ),      
               .std__pe8__lane17_strm0_data          ( std__pe8__lane17_strm0_data       ),      
               .std__pe8__lane17_strm0_data_valid    ( std__pe8__lane17_strm0_data_valid ),      
               .std__pe8__lane17_strm0_data_mask     ( std__pe8__lane17_strm0_data_mask  ),      

               .pe8__std__lane17_strm1_ready         ( pe8__std__lane17_strm1_ready      ),      
               .std__pe8__lane17_strm1_cntl          ( std__pe8__lane17_strm1_cntl       ),      
               .std__pe8__lane17_strm1_data          ( std__pe8__lane17_strm1_data       ),      
               .std__pe8__lane17_strm1_data_valid    ( std__pe8__lane17_strm1_data_valid ),      
               .std__pe8__lane17_strm1_data_mask     ( std__pe8__lane17_strm1_data_mask  ),      

               // PE 8, Lane 18                 
               .pe8__std__lane18_strm0_ready         ( pe8__std__lane18_strm0_ready      ),      
               .std__pe8__lane18_strm0_cntl          ( std__pe8__lane18_strm0_cntl       ),      
               .std__pe8__lane18_strm0_data          ( std__pe8__lane18_strm0_data       ),      
               .std__pe8__lane18_strm0_data_valid    ( std__pe8__lane18_strm0_data_valid ),      
               .std__pe8__lane18_strm0_data_mask     ( std__pe8__lane18_strm0_data_mask  ),      

               .pe8__std__lane18_strm1_ready         ( pe8__std__lane18_strm1_ready      ),      
               .std__pe8__lane18_strm1_cntl          ( std__pe8__lane18_strm1_cntl       ),      
               .std__pe8__lane18_strm1_data          ( std__pe8__lane18_strm1_data       ),      
               .std__pe8__lane18_strm1_data_valid    ( std__pe8__lane18_strm1_data_valid ),      
               .std__pe8__lane18_strm1_data_mask     ( std__pe8__lane18_strm1_data_mask  ),      

               // PE 8, Lane 19                 
               .pe8__std__lane19_strm0_ready         ( pe8__std__lane19_strm0_ready      ),      
               .std__pe8__lane19_strm0_cntl          ( std__pe8__lane19_strm0_cntl       ),      
               .std__pe8__lane19_strm0_data          ( std__pe8__lane19_strm0_data       ),      
               .std__pe8__lane19_strm0_data_valid    ( std__pe8__lane19_strm0_data_valid ),      
               .std__pe8__lane19_strm0_data_mask     ( std__pe8__lane19_strm0_data_mask  ),      

               .pe8__std__lane19_strm1_ready         ( pe8__std__lane19_strm1_ready      ),      
               .std__pe8__lane19_strm1_cntl          ( std__pe8__lane19_strm1_cntl       ),      
               .std__pe8__lane19_strm1_data          ( std__pe8__lane19_strm1_data       ),      
               .std__pe8__lane19_strm1_data_valid    ( std__pe8__lane19_strm1_data_valid ),      
               .std__pe8__lane19_strm1_data_mask     ( std__pe8__lane19_strm1_data_mask  ),      

               // PE 8, Lane 20                 
               .pe8__std__lane20_strm0_ready         ( pe8__std__lane20_strm0_ready      ),      
               .std__pe8__lane20_strm0_cntl          ( std__pe8__lane20_strm0_cntl       ),      
               .std__pe8__lane20_strm0_data          ( std__pe8__lane20_strm0_data       ),      
               .std__pe8__lane20_strm0_data_valid    ( std__pe8__lane20_strm0_data_valid ),      
               .std__pe8__lane20_strm0_data_mask     ( std__pe8__lane20_strm0_data_mask  ),      

               .pe8__std__lane20_strm1_ready         ( pe8__std__lane20_strm1_ready      ),      
               .std__pe8__lane20_strm1_cntl          ( std__pe8__lane20_strm1_cntl       ),      
               .std__pe8__lane20_strm1_data          ( std__pe8__lane20_strm1_data       ),      
               .std__pe8__lane20_strm1_data_valid    ( std__pe8__lane20_strm1_data_valid ),      
               .std__pe8__lane20_strm1_data_mask     ( std__pe8__lane20_strm1_data_mask  ),      

               // PE 8, Lane 21                 
               .pe8__std__lane21_strm0_ready         ( pe8__std__lane21_strm0_ready      ),      
               .std__pe8__lane21_strm0_cntl          ( std__pe8__lane21_strm0_cntl       ),      
               .std__pe8__lane21_strm0_data          ( std__pe8__lane21_strm0_data       ),      
               .std__pe8__lane21_strm0_data_valid    ( std__pe8__lane21_strm0_data_valid ),      
               .std__pe8__lane21_strm0_data_mask     ( std__pe8__lane21_strm0_data_mask  ),      

               .pe8__std__lane21_strm1_ready         ( pe8__std__lane21_strm1_ready      ),      
               .std__pe8__lane21_strm1_cntl          ( std__pe8__lane21_strm1_cntl       ),      
               .std__pe8__lane21_strm1_data          ( std__pe8__lane21_strm1_data       ),      
               .std__pe8__lane21_strm1_data_valid    ( std__pe8__lane21_strm1_data_valid ),      
               .std__pe8__lane21_strm1_data_mask     ( std__pe8__lane21_strm1_data_mask  ),      

               // PE 8, Lane 22                 
               .pe8__std__lane22_strm0_ready         ( pe8__std__lane22_strm0_ready      ),      
               .std__pe8__lane22_strm0_cntl          ( std__pe8__lane22_strm0_cntl       ),      
               .std__pe8__lane22_strm0_data          ( std__pe8__lane22_strm0_data       ),      
               .std__pe8__lane22_strm0_data_valid    ( std__pe8__lane22_strm0_data_valid ),      
               .std__pe8__lane22_strm0_data_mask     ( std__pe8__lane22_strm0_data_mask  ),      

               .pe8__std__lane22_strm1_ready         ( pe8__std__lane22_strm1_ready      ),      
               .std__pe8__lane22_strm1_cntl          ( std__pe8__lane22_strm1_cntl       ),      
               .std__pe8__lane22_strm1_data          ( std__pe8__lane22_strm1_data       ),      
               .std__pe8__lane22_strm1_data_valid    ( std__pe8__lane22_strm1_data_valid ),      
               .std__pe8__lane22_strm1_data_mask     ( std__pe8__lane22_strm1_data_mask  ),      

               // PE 8, Lane 23                 
               .pe8__std__lane23_strm0_ready         ( pe8__std__lane23_strm0_ready      ),      
               .std__pe8__lane23_strm0_cntl          ( std__pe8__lane23_strm0_cntl       ),      
               .std__pe8__lane23_strm0_data          ( std__pe8__lane23_strm0_data       ),      
               .std__pe8__lane23_strm0_data_valid    ( std__pe8__lane23_strm0_data_valid ),      
               .std__pe8__lane23_strm0_data_mask     ( std__pe8__lane23_strm0_data_mask  ),      

               .pe8__std__lane23_strm1_ready         ( pe8__std__lane23_strm1_ready      ),      
               .std__pe8__lane23_strm1_cntl          ( std__pe8__lane23_strm1_cntl       ),      
               .std__pe8__lane23_strm1_data          ( std__pe8__lane23_strm1_data       ),      
               .std__pe8__lane23_strm1_data_valid    ( std__pe8__lane23_strm1_data_valid ),      
               .std__pe8__lane23_strm1_data_mask     ( std__pe8__lane23_strm1_data_mask  ),      

               // PE 8, Lane 24                 
               .pe8__std__lane24_strm0_ready         ( pe8__std__lane24_strm0_ready      ),      
               .std__pe8__lane24_strm0_cntl          ( std__pe8__lane24_strm0_cntl       ),      
               .std__pe8__lane24_strm0_data          ( std__pe8__lane24_strm0_data       ),      
               .std__pe8__lane24_strm0_data_valid    ( std__pe8__lane24_strm0_data_valid ),      
               .std__pe8__lane24_strm0_data_mask     ( std__pe8__lane24_strm0_data_mask  ),      

               .pe8__std__lane24_strm1_ready         ( pe8__std__lane24_strm1_ready      ),      
               .std__pe8__lane24_strm1_cntl          ( std__pe8__lane24_strm1_cntl       ),      
               .std__pe8__lane24_strm1_data          ( std__pe8__lane24_strm1_data       ),      
               .std__pe8__lane24_strm1_data_valid    ( std__pe8__lane24_strm1_data_valid ),      
               .std__pe8__lane24_strm1_data_mask     ( std__pe8__lane24_strm1_data_mask  ),      

               // PE 8, Lane 25                 
               .pe8__std__lane25_strm0_ready         ( pe8__std__lane25_strm0_ready      ),      
               .std__pe8__lane25_strm0_cntl          ( std__pe8__lane25_strm0_cntl       ),      
               .std__pe8__lane25_strm0_data          ( std__pe8__lane25_strm0_data       ),      
               .std__pe8__lane25_strm0_data_valid    ( std__pe8__lane25_strm0_data_valid ),      
               .std__pe8__lane25_strm0_data_mask     ( std__pe8__lane25_strm0_data_mask  ),      

               .pe8__std__lane25_strm1_ready         ( pe8__std__lane25_strm1_ready      ),      
               .std__pe8__lane25_strm1_cntl          ( std__pe8__lane25_strm1_cntl       ),      
               .std__pe8__lane25_strm1_data          ( std__pe8__lane25_strm1_data       ),      
               .std__pe8__lane25_strm1_data_valid    ( std__pe8__lane25_strm1_data_valid ),      
               .std__pe8__lane25_strm1_data_mask     ( std__pe8__lane25_strm1_data_mask  ),      

               // PE 8, Lane 26                 
               .pe8__std__lane26_strm0_ready         ( pe8__std__lane26_strm0_ready      ),      
               .std__pe8__lane26_strm0_cntl          ( std__pe8__lane26_strm0_cntl       ),      
               .std__pe8__lane26_strm0_data          ( std__pe8__lane26_strm0_data       ),      
               .std__pe8__lane26_strm0_data_valid    ( std__pe8__lane26_strm0_data_valid ),      
               .std__pe8__lane26_strm0_data_mask     ( std__pe8__lane26_strm0_data_mask  ),      

               .pe8__std__lane26_strm1_ready         ( pe8__std__lane26_strm1_ready      ),      
               .std__pe8__lane26_strm1_cntl          ( std__pe8__lane26_strm1_cntl       ),      
               .std__pe8__lane26_strm1_data          ( std__pe8__lane26_strm1_data       ),      
               .std__pe8__lane26_strm1_data_valid    ( std__pe8__lane26_strm1_data_valid ),      
               .std__pe8__lane26_strm1_data_mask     ( std__pe8__lane26_strm1_data_mask  ),      

               // PE 8, Lane 27                 
               .pe8__std__lane27_strm0_ready         ( pe8__std__lane27_strm0_ready      ),      
               .std__pe8__lane27_strm0_cntl          ( std__pe8__lane27_strm0_cntl       ),      
               .std__pe8__lane27_strm0_data          ( std__pe8__lane27_strm0_data       ),      
               .std__pe8__lane27_strm0_data_valid    ( std__pe8__lane27_strm0_data_valid ),      
               .std__pe8__lane27_strm0_data_mask     ( std__pe8__lane27_strm0_data_mask  ),      

               .pe8__std__lane27_strm1_ready         ( pe8__std__lane27_strm1_ready      ),      
               .std__pe8__lane27_strm1_cntl          ( std__pe8__lane27_strm1_cntl       ),      
               .std__pe8__lane27_strm1_data          ( std__pe8__lane27_strm1_data       ),      
               .std__pe8__lane27_strm1_data_valid    ( std__pe8__lane27_strm1_data_valid ),      
               .std__pe8__lane27_strm1_data_mask     ( std__pe8__lane27_strm1_data_mask  ),      

               // PE 8, Lane 28                 
               .pe8__std__lane28_strm0_ready         ( pe8__std__lane28_strm0_ready      ),      
               .std__pe8__lane28_strm0_cntl          ( std__pe8__lane28_strm0_cntl       ),      
               .std__pe8__lane28_strm0_data          ( std__pe8__lane28_strm0_data       ),      
               .std__pe8__lane28_strm0_data_valid    ( std__pe8__lane28_strm0_data_valid ),      
               .std__pe8__lane28_strm0_data_mask     ( std__pe8__lane28_strm0_data_mask  ),      

               .pe8__std__lane28_strm1_ready         ( pe8__std__lane28_strm1_ready      ),      
               .std__pe8__lane28_strm1_cntl          ( std__pe8__lane28_strm1_cntl       ),      
               .std__pe8__lane28_strm1_data          ( std__pe8__lane28_strm1_data       ),      
               .std__pe8__lane28_strm1_data_valid    ( std__pe8__lane28_strm1_data_valid ),      
               .std__pe8__lane28_strm1_data_mask     ( std__pe8__lane28_strm1_data_mask  ),      

               // PE 8, Lane 29                 
               .pe8__std__lane29_strm0_ready         ( pe8__std__lane29_strm0_ready      ),      
               .std__pe8__lane29_strm0_cntl          ( std__pe8__lane29_strm0_cntl       ),      
               .std__pe8__lane29_strm0_data          ( std__pe8__lane29_strm0_data       ),      
               .std__pe8__lane29_strm0_data_valid    ( std__pe8__lane29_strm0_data_valid ),      
               .std__pe8__lane29_strm0_data_mask     ( std__pe8__lane29_strm0_data_mask  ),      

               .pe8__std__lane29_strm1_ready         ( pe8__std__lane29_strm1_ready      ),      
               .std__pe8__lane29_strm1_cntl          ( std__pe8__lane29_strm1_cntl       ),      
               .std__pe8__lane29_strm1_data          ( std__pe8__lane29_strm1_data       ),      
               .std__pe8__lane29_strm1_data_valid    ( std__pe8__lane29_strm1_data_valid ),      
               .std__pe8__lane29_strm1_data_mask     ( std__pe8__lane29_strm1_data_mask  ),      

               // PE 8, Lane 30                 
               .pe8__std__lane30_strm0_ready         ( pe8__std__lane30_strm0_ready      ),      
               .std__pe8__lane30_strm0_cntl          ( std__pe8__lane30_strm0_cntl       ),      
               .std__pe8__lane30_strm0_data          ( std__pe8__lane30_strm0_data       ),      
               .std__pe8__lane30_strm0_data_valid    ( std__pe8__lane30_strm0_data_valid ),      
               .std__pe8__lane30_strm0_data_mask     ( std__pe8__lane30_strm0_data_mask  ),      

               .pe8__std__lane30_strm1_ready         ( pe8__std__lane30_strm1_ready      ),      
               .std__pe8__lane30_strm1_cntl          ( std__pe8__lane30_strm1_cntl       ),      
               .std__pe8__lane30_strm1_data          ( std__pe8__lane30_strm1_data       ),      
               .std__pe8__lane30_strm1_data_valid    ( std__pe8__lane30_strm1_data_valid ),      
               .std__pe8__lane30_strm1_data_mask     ( std__pe8__lane30_strm1_data_mask  ),      

               // PE 8, Lane 31                 
               .pe8__std__lane31_strm0_ready         ( pe8__std__lane31_strm0_ready      ),      
               .std__pe8__lane31_strm0_cntl          ( std__pe8__lane31_strm0_cntl       ),      
               .std__pe8__lane31_strm0_data          ( std__pe8__lane31_strm0_data       ),      
               .std__pe8__lane31_strm0_data_valid    ( std__pe8__lane31_strm0_data_valid ),      
               .std__pe8__lane31_strm0_data_mask     ( std__pe8__lane31_strm0_data_mask  ),      

               .pe8__std__lane31_strm1_ready         ( pe8__std__lane31_strm1_ready      ),      
               .std__pe8__lane31_strm1_cntl          ( std__pe8__lane31_strm1_cntl       ),      
               .std__pe8__lane31_strm1_data          ( std__pe8__lane31_strm1_data       ),      
               .std__pe8__lane31_strm1_data_valid    ( std__pe8__lane31_strm1_data_valid ),      
               .std__pe8__lane31_strm1_data_mask     ( std__pe8__lane31_strm1_data_mask  ),      

               // PE 9, Lane 0                 
               .pe9__std__lane0_strm0_ready         ( pe9__std__lane0_strm0_ready      ),      
               .std__pe9__lane0_strm0_cntl          ( std__pe9__lane0_strm0_cntl       ),      
               .std__pe9__lane0_strm0_data          ( std__pe9__lane0_strm0_data       ),      
               .std__pe9__lane0_strm0_data_valid    ( std__pe9__lane0_strm0_data_valid ),      
               .std__pe9__lane0_strm0_data_mask     ( std__pe9__lane0_strm0_data_mask  ),      

               .pe9__std__lane0_strm1_ready         ( pe9__std__lane0_strm1_ready      ),      
               .std__pe9__lane0_strm1_cntl          ( std__pe9__lane0_strm1_cntl       ),      
               .std__pe9__lane0_strm1_data          ( std__pe9__lane0_strm1_data       ),      
               .std__pe9__lane0_strm1_data_valid    ( std__pe9__lane0_strm1_data_valid ),      
               .std__pe9__lane0_strm1_data_mask     ( std__pe9__lane0_strm1_data_mask  ),      

               // PE 9, Lane 1                 
               .pe9__std__lane1_strm0_ready         ( pe9__std__lane1_strm0_ready      ),      
               .std__pe9__lane1_strm0_cntl          ( std__pe9__lane1_strm0_cntl       ),      
               .std__pe9__lane1_strm0_data          ( std__pe9__lane1_strm0_data       ),      
               .std__pe9__lane1_strm0_data_valid    ( std__pe9__lane1_strm0_data_valid ),      
               .std__pe9__lane1_strm0_data_mask     ( std__pe9__lane1_strm0_data_mask  ),      

               .pe9__std__lane1_strm1_ready         ( pe9__std__lane1_strm1_ready      ),      
               .std__pe9__lane1_strm1_cntl          ( std__pe9__lane1_strm1_cntl       ),      
               .std__pe9__lane1_strm1_data          ( std__pe9__lane1_strm1_data       ),      
               .std__pe9__lane1_strm1_data_valid    ( std__pe9__lane1_strm1_data_valid ),      
               .std__pe9__lane1_strm1_data_mask     ( std__pe9__lane1_strm1_data_mask  ),      

               // PE 9, Lane 2                 
               .pe9__std__lane2_strm0_ready         ( pe9__std__lane2_strm0_ready      ),      
               .std__pe9__lane2_strm0_cntl          ( std__pe9__lane2_strm0_cntl       ),      
               .std__pe9__lane2_strm0_data          ( std__pe9__lane2_strm0_data       ),      
               .std__pe9__lane2_strm0_data_valid    ( std__pe9__lane2_strm0_data_valid ),      
               .std__pe9__lane2_strm0_data_mask     ( std__pe9__lane2_strm0_data_mask  ),      

               .pe9__std__lane2_strm1_ready         ( pe9__std__lane2_strm1_ready      ),      
               .std__pe9__lane2_strm1_cntl          ( std__pe9__lane2_strm1_cntl       ),      
               .std__pe9__lane2_strm1_data          ( std__pe9__lane2_strm1_data       ),      
               .std__pe9__lane2_strm1_data_valid    ( std__pe9__lane2_strm1_data_valid ),      
               .std__pe9__lane2_strm1_data_mask     ( std__pe9__lane2_strm1_data_mask  ),      

               // PE 9, Lane 3                 
               .pe9__std__lane3_strm0_ready         ( pe9__std__lane3_strm0_ready      ),      
               .std__pe9__lane3_strm0_cntl          ( std__pe9__lane3_strm0_cntl       ),      
               .std__pe9__lane3_strm0_data          ( std__pe9__lane3_strm0_data       ),      
               .std__pe9__lane3_strm0_data_valid    ( std__pe9__lane3_strm0_data_valid ),      
               .std__pe9__lane3_strm0_data_mask     ( std__pe9__lane3_strm0_data_mask  ),      

               .pe9__std__lane3_strm1_ready         ( pe9__std__lane3_strm1_ready      ),      
               .std__pe9__lane3_strm1_cntl          ( std__pe9__lane3_strm1_cntl       ),      
               .std__pe9__lane3_strm1_data          ( std__pe9__lane3_strm1_data       ),      
               .std__pe9__lane3_strm1_data_valid    ( std__pe9__lane3_strm1_data_valid ),      
               .std__pe9__lane3_strm1_data_mask     ( std__pe9__lane3_strm1_data_mask  ),      

               // PE 9, Lane 4                 
               .pe9__std__lane4_strm0_ready         ( pe9__std__lane4_strm0_ready      ),      
               .std__pe9__lane4_strm0_cntl          ( std__pe9__lane4_strm0_cntl       ),      
               .std__pe9__lane4_strm0_data          ( std__pe9__lane4_strm0_data       ),      
               .std__pe9__lane4_strm0_data_valid    ( std__pe9__lane4_strm0_data_valid ),      
               .std__pe9__lane4_strm0_data_mask     ( std__pe9__lane4_strm0_data_mask  ),      

               .pe9__std__lane4_strm1_ready         ( pe9__std__lane4_strm1_ready      ),      
               .std__pe9__lane4_strm1_cntl          ( std__pe9__lane4_strm1_cntl       ),      
               .std__pe9__lane4_strm1_data          ( std__pe9__lane4_strm1_data       ),      
               .std__pe9__lane4_strm1_data_valid    ( std__pe9__lane4_strm1_data_valid ),      
               .std__pe9__lane4_strm1_data_mask     ( std__pe9__lane4_strm1_data_mask  ),      

               // PE 9, Lane 5                 
               .pe9__std__lane5_strm0_ready         ( pe9__std__lane5_strm0_ready      ),      
               .std__pe9__lane5_strm0_cntl          ( std__pe9__lane5_strm0_cntl       ),      
               .std__pe9__lane5_strm0_data          ( std__pe9__lane5_strm0_data       ),      
               .std__pe9__lane5_strm0_data_valid    ( std__pe9__lane5_strm0_data_valid ),      
               .std__pe9__lane5_strm0_data_mask     ( std__pe9__lane5_strm0_data_mask  ),      

               .pe9__std__lane5_strm1_ready         ( pe9__std__lane5_strm1_ready      ),      
               .std__pe9__lane5_strm1_cntl          ( std__pe9__lane5_strm1_cntl       ),      
               .std__pe9__lane5_strm1_data          ( std__pe9__lane5_strm1_data       ),      
               .std__pe9__lane5_strm1_data_valid    ( std__pe9__lane5_strm1_data_valid ),      
               .std__pe9__lane5_strm1_data_mask     ( std__pe9__lane5_strm1_data_mask  ),      

               // PE 9, Lane 6                 
               .pe9__std__lane6_strm0_ready         ( pe9__std__lane6_strm0_ready      ),      
               .std__pe9__lane6_strm0_cntl          ( std__pe9__lane6_strm0_cntl       ),      
               .std__pe9__lane6_strm0_data          ( std__pe9__lane6_strm0_data       ),      
               .std__pe9__lane6_strm0_data_valid    ( std__pe9__lane6_strm0_data_valid ),      
               .std__pe9__lane6_strm0_data_mask     ( std__pe9__lane6_strm0_data_mask  ),      

               .pe9__std__lane6_strm1_ready         ( pe9__std__lane6_strm1_ready      ),      
               .std__pe9__lane6_strm1_cntl          ( std__pe9__lane6_strm1_cntl       ),      
               .std__pe9__lane6_strm1_data          ( std__pe9__lane6_strm1_data       ),      
               .std__pe9__lane6_strm1_data_valid    ( std__pe9__lane6_strm1_data_valid ),      
               .std__pe9__lane6_strm1_data_mask     ( std__pe9__lane6_strm1_data_mask  ),      

               // PE 9, Lane 7                 
               .pe9__std__lane7_strm0_ready         ( pe9__std__lane7_strm0_ready      ),      
               .std__pe9__lane7_strm0_cntl          ( std__pe9__lane7_strm0_cntl       ),      
               .std__pe9__lane7_strm0_data          ( std__pe9__lane7_strm0_data       ),      
               .std__pe9__lane7_strm0_data_valid    ( std__pe9__lane7_strm0_data_valid ),      
               .std__pe9__lane7_strm0_data_mask     ( std__pe9__lane7_strm0_data_mask  ),      

               .pe9__std__lane7_strm1_ready         ( pe9__std__lane7_strm1_ready      ),      
               .std__pe9__lane7_strm1_cntl          ( std__pe9__lane7_strm1_cntl       ),      
               .std__pe9__lane7_strm1_data          ( std__pe9__lane7_strm1_data       ),      
               .std__pe9__lane7_strm1_data_valid    ( std__pe9__lane7_strm1_data_valid ),      
               .std__pe9__lane7_strm1_data_mask     ( std__pe9__lane7_strm1_data_mask  ),      

               // PE 9, Lane 8                 
               .pe9__std__lane8_strm0_ready         ( pe9__std__lane8_strm0_ready      ),      
               .std__pe9__lane8_strm0_cntl          ( std__pe9__lane8_strm0_cntl       ),      
               .std__pe9__lane8_strm0_data          ( std__pe9__lane8_strm0_data       ),      
               .std__pe9__lane8_strm0_data_valid    ( std__pe9__lane8_strm0_data_valid ),      
               .std__pe9__lane8_strm0_data_mask     ( std__pe9__lane8_strm0_data_mask  ),      

               .pe9__std__lane8_strm1_ready         ( pe9__std__lane8_strm1_ready      ),      
               .std__pe9__lane8_strm1_cntl          ( std__pe9__lane8_strm1_cntl       ),      
               .std__pe9__lane8_strm1_data          ( std__pe9__lane8_strm1_data       ),      
               .std__pe9__lane8_strm1_data_valid    ( std__pe9__lane8_strm1_data_valid ),      
               .std__pe9__lane8_strm1_data_mask     ( std__pe9__lane8_strm1_data_mask  ),      

               // PE 9, Lane 9                 
               .pe9__std__lane9_strm0_ready         ( pe9__std__lane9_strm0_ready      ),      
               .std__pe9__lane9_strm0_cntl          ( std__pe9__lane9_strm0_cntl       ),      
               .std__pe9__lane9_strm0_data          ( std__pe9__lane9_strm0_data       ),      
               .std__pe9__lane9_strm0_data_valid    ( std__pe9__lane9_strm0_data_valid ),      
               .std__pe9__lane9_strm0_data_mask     ( std__pe9__lane9_strm0_data_mask  ),      

               .pe9__std__lane9_strm1_ready         ( pe9__std__lane9_strm1_ready      ),      
               .std__pe9__lane9_strm1_cntl          ( std__pe9__lane9_strm1_cntl       ),      
               .std__pe9__lane9_strm1_data          ( std__pe9__lane9_strm1_data       ),      
               .std__pe9__lane9_strm1_data_valid    ( std__pe9__lane9_strm1_data_valid ),      
               .std__pe9__lane9_strm1_data_mask     ( std__pe9__lane9_strm1_data_mask  ),      

               // PE 9, Lane 10                 
               .pe9__std__lane10_strm0_ready         ( pe9__std__lane10_strm0_ready      ),      
               .std__pe9__lane10_strm0_cntl          ( std__pe9__lane10_strm0_cntl       ),      
               .std__pe9__lane10_strm0_data          ( std__pe9__lane10_strm0_data       ),      
               .std__pe9__lane10_strm0_data_valid    ( std__pe9__lane10_strm0_data_valid ),      
               .std__pe9__lane10_strm0_data_mask     ( std__pe9__lane10_strm0_data_mask  ),      

               .pe9__std__lane10_strm1_ready         ( pe9__std__lane10_strm1_ready      ),      
               .std__pe9__lane10_strm1_cntl          ( std__pe9__lane10_strm1_cntl       ),      
               .std__pe9__lane10_strm1_data          ( std__pe9__lane10_strm1_data       ),      
               .std__pe9__lane10_strm1_data_valid    ( std__pe9__lane10_strm1_data_valid ),      
               .std__pe9__lane10_strm1_data_mask     ( std__pe9__lane10_strm1_data_mask  ),      

               // PE 9, Lane 11                 
               .pe9__std__lane11_strm0_ready         ( pe9__std__lane11_strm0_ready      ),      
               .std__pe9__lane11_strm0_cntl          ( std__pe9__lane11_strm0_cntl       ),      
               .std__pe9__lane11_strm0_data          ( std__pe9__lane11_strm0_data       ),      
               .std__pe9__lane11_strm0_data_valid    ( std__pe9__lane11_strm0_data_valid ),      
               .std__pe9__lane11_strm0_data_mask     ( std__pe9__lane11_strm0_data_mask  ),      

               .pe9__std__lane11_strm1_ready         ( pe9__std__lane11_strm1_ready      ),      
               .std__pe9__lane11_strm1_cntl          ( std__pe9__lane11_strm1_cntl       ),      
               .std__pe9__lane11_strm1_data          ( std__pe9__lane11_strm1_data       ),      
               .std__pe9__lane11_strm1_data_valid    ( std__pe9__lane11_strm1_data_valid ),      
               .std__pe9__lane11_strm1_data_mask     ( std__pe9__lane11_strm1_data_mask  ),      

               // PE 9, Lane 12                 
               .pe9__std__lane12_strm0_ready         ( pe9__std__lane12_strm0_ready      ),      
               .std__pe9__lane12_strm0_cntl          ( std__pe9__lane12_strm0_cntl       ),      
               .std__pe9__lane12_strm0_data          ( std__pe9__lane12_strm0_data       ),      
               .std__pe9__lane12_strm0_data_valid    ( std__pe9__lane12_strm0_data_valid ),      
               .std__pe9__lane12_strm0_data_mask     ( std__pe9__lane12_strm0_data_mask  ),      

               .pe9__std__lane12_strm1_ready         ( pe9__std__lane12_strm1_ready      ),      
               .std__pe9__lane12_strm1_cntl          ( std__pe9__lane12_strm1_cntl       ),      
               .std__pe9__lane12_strm1_data          ( std__pe9__lane12_strm1_data       ),      
               .std__pe9__lane12_strm1_data_valid    ( std__pe9__lane12_strm1_data_valid ),      
               .std__pe9__lane12_strm1_data_mask     ( std__pe9__lane12_strm1_data_mask  ),      

               // PE 9, Lane 13                 
               .pe9__std__lane13_strm0_ready         ( pe9__std__lane13_strm0_ready      ),      
               .std__pe9__lane13_strm0_cntl          ( std__pe9__lane13_strm0_cntl       ),      
               .std__pe9__lane13_strm0_data          ( std__pe9__lane13_strm0_data       ),      
               .std__pe9__lane13_strm0_data_valid    ( std__pe9__lane13_strm0_data_valid ),      
               .std__pe9__lane13_strm0_data_mask     ( std__pe9__lane13_strm0_data_mask  ),      

               .pe9__std__lane13_strm1_ready         ( pe9__std__lane13_strm1_ready      ),      
               .std__pe9__lane13_strm1_cntl          ( std__pe9__lane13_strm1_cntl       ),      
               .std__pe9__lane13_strm1_data          ( std__pe9__lane13_strm1_data       ),      
               .std__pe9__lane13_strm1_data_valid    ( std__pe9__lane13_strm1_data_valid ),      
               .std__pe9__lane13_strm1_data_mask     ( std__pe9__lane13_strm1_data_mask  ),      

               // PE 9, Lane 14                 
               .pe9__std__lane14_strm0_ready         ( pe9__std__lane14_strm0_ready      ),      
               .std__pe9__lane14_strm0_cntl          ( std__pe9__lane14_strm0_cntl       ),      
               .std__pe9__lane14_strm0_data          ( std__pe9__lane14_strm0_data       ),      
               .std__pe9__lane14_strm0_data_valid    ( std__pe9__lane14_strm0_data_valid ),      
               .std__pe9__lane14_strm0_data_mask     ( std__pe9__lane14_strm0_data_mask  ),      

               .pe9__std__lane14_strm1_ready         ( pe9__std__lane14_strm1_ready      ),      
               .std__pe9__lane14_strm1_cntl          ( std__pe9__lane14_strm1_cntl       ),      
               .std__pe9__lane14_strm1_data          ( std__pe9__lane14_strm1_data       ),      
               .std__pe9__lane14_strm1_data_valid    ( std__pe9__lane14_strm1_data_valid ),      
               .std__pe9__lane14_strm1_data_mask     ( std__pe9__lane14_strm1_data_mask  ),      

               // PE 9, Lane 15                 
               .pe9__std__lane15_strm0_ready         ( pe9__std__lane15_strm0_ready      ),      
               .std__pe9__lane15_strm0_cntl          ( std__pe9__lane15_strm0_cntl       ),      
               .std__pe9__lane15_strm0_data          ( std__pe9__lane15_strm0_data       ),      
               .std__pe9__lane15_strm0_data_valid    ( std__pe9__lane15_strm0_data_valid ),      
               .std__pe9__lane15_strm0_data_mask     ( std__pe9__lane15_strm0_data_mask  ),      

               .pe9__std__lane15_strm1_ready         ( pe9__std__lane15_strm1_ready      ),      
               .std__pe9__lane15_strm1_cntl          ( std__pe9__lane15_strm1_cntl       ),      
               .std__pe9__lane15_strm1_data          ( std__pe9__lane15_strm1_data       ),      
               .std__pe9__lane15_strm1_data_valid    ( std__pe9__lane15_strm1_data_valid ),      
               .std__pe9__lane15_strm1_data_mask     ( std__pe9__lane15_strm1_data_mask  ),      

               // PE 9, Lane 16                 
               .pe9__std__lane16_strm0_ready         ( pe9__std__lane16_strm0_ready      ),      
               .std__pe9__lane16_strm0_cntl          ( std__pe9__lane16_strm0_cntl       ),      
               .std__pe9__lane16_strm0_data          ( std__pe9__lane16_strm0_data       ),      
               .std__pe9__lane16_strm0_data_valid    ( std__pe9__lane16_strm0_data_valid ),      
               .std__pe9__lane16_strm0_data_mask     ( std__pe9__lane16_strm0_data_mask  ),      

               .pe9__std__lane16_strm1_ready         ( pe9__std__lane16_strm1_ready      ),      
               .std__pe9__lane16_strm1_cntl          ( std__pe9__lane16_strm1_cntl       ),      
               .std__pe9__lane16_strm1_data          ( std__pe9__lane16_strm1_data       ),      
               .std__pe9__lane16_strm1_data_valid    ( std__pe9__lane16_strm1_data_valid ),      
               .std__pe9__lane16_strm1_data_mask     ( std__pe9__lane16_strm1_data_mask  ),      

               // PE 9, Lane 17                 
               .pe9__std__lane17_strm0_ready         ( pe9__std__lane17_strm0_ready      ),      
               .std__pe9__lane17_strm0_cntl          ( std__pe9__lane17_strm0_cntl       ),      
               .std__pe9__lane17_strm0_data          ( std__pe9__lane17_strm0_data       ),      
               .std__pe9__lane17_strm0_data_valid    ( std__pe9__lane17_strm0_data_valid ),      
               .std__pe9__lane17_strm0_data_mask     ( std__pe9__lane17_strm0_data_mask  ),      

               .pe9__std__lane17_strm1_ready         ( pe9__std__lane17_strm1_ready      ),      
               .std__pe9__lane17_strm1_cntl          ( std__pe9__lane17_strm1_cntl       ),      
               .std__pe9__lane17_strm1_data          ( std__pe9__lane17_strm1_data       ),      
               .std__pe9__lane17_strm1_data_valid    ( std__pe9__lane17_strm1_data_valid ),      
               .std__pe9__lane17_strm1_data_mask     ( std__pe9__lane17_strm1_data_mask  ),      

               // PE 9, Lane 18                 
               .pe9__std__lane18_strm0_ready         ( pe9__std__lane18_strm0_ready      ),      
               .std__pe9__lane18_strm0_cntl          ( std__pe9__lane18_strm0_cntl       ),      
               .std__pe9__lane18_strm0_data          ( std__pe9__lane18_strm0_data       ),      
               .std__pe9__lane18_strm0_data_valid    ( std__pe9__lane18_strm0_data_valid ),      
               .std__pe9__lane18_strm0_data_mask     ( std__pe9__lane18_strm0_data_mask  ),      

               .pe9__std__lane18_strm1_ready         ( pe9__std__lane18_strm1_ready      ),      
               .std__pe9__lane18_strm1_cntl          ( std__pe9__lane18_strm1_cntl       ),      
               .std__pe9__lane18_strm1_data          ( std__pe9__lane18_strm1_data       ),      
               .std__pe9__lane18_strm1_data_valid    ( std__pe9__lane18_strm1_data_valid ),      
               .std__pe9__lane18_strm1_data_mask     ( std__pe9__lane18_strm1_data_mask  ),      

               // PE 9, Lane 19                 
               .pe9__std__lane19_strm0_ready         ( pe9__std__lane19_strm0_ready      ),      
               .std__pe9__lane19_strm0_cntl          ( std__pe9__lane19_strm0_cntl       ),      
               .std__pe9__lane19_strm0_data          ( std__pe9__lane19_strm0_data       ),      
               .std__pe9__lane19_strm0_data_valid    ( std__pe9__lane19_strm0_data_valid ),      
               .std__pe9__lane19_strm0_data_mask     ( std__pe9__lane19_strm0_data_mask  ),      

               .pe9__std__lane19_strm1_ready         ( pe9__std__lane19_strm1_ready      ),      
               .std__pe9__lane19_strm1_cntl          ( std__pe9__lane19_strm1_cntl       ),      
               .std__pe9__lane19_strm1_data          ( std__pe9__lane19_strm1_data       ),      
               .std__pe9__lane19_strm1_data_valid    ( std__pe9__lane19_strm1_data_valid ),      
               .std__pe9__lane19_strm1_data_mask     ( std__pe9__lane19_strm1_data_mask  ),      

               // PE 9, Lane 20                 
               .pe9__std__lane20_strm0_ready         ( pe9__std__lane20_strm0_ready      ),      
               .std__pe9__lane20_strm0_cntl          ( std__pe9__lane20_strm0_cntl       ),      
               .std__pe9__lane20_strm0_data          ( std__pe9__lane20_strm0_data       ),      
               .std__pe9__lane20_strm0_data_valid    ( std__pe9__lane20_strm0_data_valid ),      
               .std__pe9__lane20_strm0_data_mask     ( std__pe9__lane20_strm0_data_mask  ),      

               .pe9__std__lane20_strm1_ready         ( pe9__std__lane20_strm1_ready      ),      
               .std__pe9__lane20_strm1_cntl          ( std__pe9__lane20_strm1_cntl       ),      
               .std__pe9__lane20_strm1_data          ( std__pe9__lane20_strm1_data       ),      
               .std__pe9__lane20_strm1_data_valid    ( std__pe9__lane20_strm1_data_valid ),      
               .std__pe9__lane20_strm1_data_mask     ( std__pe9__lane20_strm1_data_mask  ),      

               // PE 9, Lane 21                 
               .pe9__std__lane21_strm0_ready         ( pe9__std__lane21_strm0_ready      ),      
               .std__pe9__lane21_strm0_cntl          ( std__pe9__lane21_strm0_cntl       ),      
               .std__pe9__lane21_strm0_data          ( std__pe9__lane21_strm0_data       ),      
               .std__pe9__lane21_strm0_data_valid    ( std__pe9__lane21_strm0_data_valid ),      
               .std__pe9__lane21_strm0_data_mask     ( std__pe9__lane21_strm0_data_mask  ),      

               .pe9__std__lane21_strm1_ready         ( pe9__std__lane21_strm1_ready      ),      
               .std__pe9__lane21_strm1_cntl          ( std__pe9__lane21_strm1_cntl       ),      
               .std__pe9__lane21_strm1_data          ( std__pe9__lane21_strm1_data       ),      
               .std__pe9__lane21_strm1_data_valid    ( std__pe9__lane21_strm1_data_valid ),      
               .std__pe9__lane21_strm1_data_mask     ( std__pe9__lane21_strm1_data_mask  ),      

               // PE 9, Lane 22                 
               .pe9__std__lane22_strm0_ready         ( pe9__std__lane22_strm0_ready      ),      
               .std__pe9__lane22_strm0_cntl          ( std__pe9__lane22_strm0_cntl       ),      
               .std__pe9__lane22_strm0_data          ( std__pe9__lane22_strm0_data       ),      
               .std__pe9__lane22_strm0_data_valid    ( std__pe9__lane22_strm0_data_valid ),      
               .std__pe9__lane22_strm0_data_mask     ( std__pe9__lane22_strm0_data_mask  ),      

               .pe9__std__lane22_strm1_ready         ( pe9__std__lane22_strm1_ready      ),      
               .std__pe9__lane22_strm1_cntl          ( std__pe9__lane22_strm1_cntl       ),      
               .std__pe9__lane22_strm1_data          ( std__pe9__lane22_strm1_data       ),      
               .std__pe9__lane22_strm1_data_valid    ( std__pe9__lane22_strm1_data_valid ),      
               .std__pe9__lane22_strm1_data_mask     ( std__pe9__lane22_strm1_data_mask  ),      

               // PE 9, Lane 23                 
               .pe9__std__lane23_strm0_ready         ( pe9__std__lane23_strm0_ready      ),      
               .std__pe9__lane23_strm0_cntl          ( std__pe9__lane23_strm0_cntl       ),      
               .std__pe9__lane23_strm0_data          ( std__pe9__lane23_strm0_data       ),      
               .std__pe9__lane23_strm0_data_valid    ( std__pe9__lane23_strm0_data_valid ),      
               .std__pe9__lane23_strm0_data_mask     ( std__pe9__lane23_strm0_data_mask  ),      

               .pe9__std__lane23_strm1_ready         ( pe9__std__lane23_strm1_ready      ),      
               .std__pe9__lane23_strm1_cntl          ( std__pe9__lane23_strm1_cntl       ),      
               .std__pe9__lane23_strm1_data          ( std__pe9__lane23_strm1_data       ),      
               .std__pe9__lane23_strm1_data_valid    ( std__pe9__lane23_strm1_data_valid ),      
               .std__pe9__lane23_strm1_data_mask     ( std__pe9__lane23_strm1_data_mask  ),      

               // PE 9, Lane 24                 
               .pe9__std__lane24_strm0_ready         ( pe9__std__lane24_strm0_ready      ),      
               .std__pe9__lane24_strm0_cntl          ( std__pe9__lane24_strm0_cntl       ),      
               .std__pe9__lane24_strm0_data          ( std__pe9__lane24_strm0_data       ),      
               .std__pe9__lane24_strm0_data_valid    ( std__pe9__lane24_strm0_data_valid ),      
               .std__pe9__lane24_strm0_data_mask     ( std__pe9__lane24_strm0_data_mask  ),      

               .pe9__std__lane24_strm1_ready         ( pe9__std__lane24_strm1_ready      ),      
               .std__pe9__lane24_strm1_cntl          ( std__pe9__lane24_strm1_cntl       ),      
               .std__pe9__lane24_strm1_data          ( std__pe9__lane24_strm1_data       ),      
               .std__pe9__lane24_strm1_data_valid    ( std__pe9__lane24_strm1_data_valid ),      
               .std__pe9__lane24_strm1_data_mask     ( std__pe9__lane24_strm1_data_mask  ),      

               // PE 9, Lane 25                 
               .pe9__std__lane25_strm0_ready         ( pe9__std__lane25_strm0_ready      ),      
               .std__pe9__lane25_strm0_cntl          ( std__pe9__lane25_strm0_cntl       ),      
               .std__pe9__lane25_strm0_data          ( std__pe9__lane25_strm0_data       ),      
               .std__pe9__lane25_strm0_data_valid    ( std__pe9__lane25_strm0_data_valid ),      
               .std__pe9__lane25_strm0_data_mask     ( std__pe9__lane25_strm0_data_mask  ),      

               .pe9__std__lane25_strm1_ready         ( pe9__std__lane25_strm1_ready      ),      
               .std__pe9__lane25_strm1_cntl          ( std__pe9__lane25_strm1_cntl       ),      
               .std__pe9__lane25_strm1_data          ( std__pe9__lane25_strm1_data       ),      
               .std__pe9__lane25_strm1_data_valid    ( std__pe9__lane25_strm1_data_valid ),      
               .std__pe9__lane25_strm1_data_mask     ( std__pe9__lane25_strm1_data_mask  ),      

               // PE 9, Lane 26                 
               .pe9__std__lane26_strm0_ready         ( pe9__std__lane26_strm0_ready      ),      
               .std__pe9__lane26_strm0_cntl          ( std__pe9__lane26_strm0_cntl       ),      
               .std__pe9__lane26_strm0_data          ( std__pe9__lane26_strm0_data       ),      
               .std__pe9__lane26_strm0_data_valid    ( std__pe9__lane26_strm0_data_valid ),      
               .std__pe9__lane26_strm0_data_mask     ( std__pe9__lane26_strm0_data_mask  ),      

               .pe9__std__lane26_strm1_ready         ( pe9__std__lane26_strm1_ready      ),      
               .std__pe9__lane26_strm1_cntl          ( std__pe9__lane26_strm1_cntl       ),      
               .std__pe9__lane26_strm1_data          ( std__pe9__lane26_strm1_data       ),      
               .std__pe9__lane26_strm1_data_valid    ( std__pe9__lane26_strm1_data_valid ),      
               .std__pe9__lane26_strm1_data_mask     ( std__pe9__lane26_strm1_data_mask  ),      

               // PE 9, Lane 27                 
               .pe9__std__lane27_strm0_ready         ( pe9__std__lane27_strm0_ready      ),      
               .std__pe9__lane27_strm0_cntl          ( std__pe9__lane27_strm0_cntl       ),      
               .std__pe9__lane27_strm0_data          ( std__pe9__lane27_strm0_data       ),      
               .std__pe9__lane27_strm0_data_valid    ( std__pe9__lane27_strm0_data_valid ),      
               .std__pe9__lane27_strm0_data_mask     ( std__pe9__lane27_strm0_data_mask  ),      

               .pe9__std__lane27_strm1_ready         ( pe9__std__lane27_strm1_ready      ),      
               .std__pe9__lane27_strm1_cntl          ( std__pe9__lane27_strm1_cntl       ),      
               .std__pe9__lane27_strm1_data          ( std__pe9__lane27_strm1_data       ),      
               .std__pe9__lane27_strm1_data_valid    ( std__pe9__lane27_strm1_data_valid ),      
               .std__pe9__lane27_strm1_data_mask     ( std__pe9__lane27_strm1_data_mask  ),      

               // PE 9, Lane 28                 
               .pe9__std__lane28_strm0_ready         ( pe9__std__lane28_strm0_ready      ),      
               .std__pe9__lane28_strm0_cntl          ( std__pe9__lane28_strm0_cntl       ),      
               .std__pe9__lane28_strm0_data          ( std__pe9__lane28_strm0_data       ),      
               .std__pe9__lane28_strm0_data_valid    ( std__pe9__lane28_strm0_data_valid ),      
               .std__pe9__lane28_strm0_data_mask     ( std__pe9__lane28_strm0_data_mask  ),      

               .pe9__std__lane28_strm1_ready         ( pe9__std__lane28_strm1_ready      ),      
               .std__pe9__lane28_strm1_cntl          ( std__pe9__lane28_strm1_cntl       ),      
               .std__pe9__lane28_strm1_data          ( std__pe9__lane28_strm1_data       ),      
               .std__pe9__lane28_strm1_data_valid    ( std__pe9__lane28_strm1_data_valid ),      
               .std__pe9__lane28_strm1_data_mask     ( std__pe9__lane28_strm1_data_mask  ),      

               // PE 9, Lane 29                 
               .pe9__std__lane29_strm0_ready         ( pe9__std__lane29_strm0_ready      ),      
               .std__pe9__lane29_strm0_cntl          ( std__pe9__lane29_strm0_cntl       ),      
               .std__pe9__lane29_strm0_data          ( std__pe9__lane29_strm0_data       ),      
               .std__pe9__lane29_strm0_data_valid    ( std__pe9__lane29_strm0_data_valid ),      
               .std__pe9__lane29_strm0_data_mask     ( std__pe9__lane29_strm0_data_mask  ),      

               .pe9__std__lane29_strm1_ready         ( pe9__std__lane29_strm1_ready      ),      
               .std__pe9__lane29_strm1_cntl          ( std__pe9__lane29_strm1_cntl       ),      
               .std__pe9__lane29_strm1_data          ( std__pe9__lane29_strm1_data       ),      
               .std__pe9__lane29_strm1_data_valid    ( std__pe9__lane29_strm1_data_valid ),      
               .std__pe9__lane29_strm1_data_mask     ( std__pe9__lane29_strm1_data_mask  ),      

               // PE 9, Lane 30                 
               .pe9__std__lane30_strm0_ready         ( pe9__std__lane30_strm0_ready      ),      
               .std__pe9__lane30_strm0_cntl          ( std__pe9__lane30_strm0_cntl       ),      
               .std__pe9__lane30_strm0_data          ( std__pe9__lane30_strm0_data       ),      
               .std__pe9__lane30_strm0_data_valid    ( std__pe9__lane30_strm0_data_valid ),      
               .std__pe9__lane30_strm0_data_mask     ( std__pe9__lane30_strm0_data_mask  ),      

               .pe9__std__lane30_strm1_ready         ( pe9__std__lane30_strm1_ready      ),      
               .std__pe9__lane30_strm1_cntl          ( std__pe9__lane30_strm1_cntl       ),      
               .std__pe9__lane30_strm1_data          ( std__pe9__lane30_strm1_data       ),      
               .std__pe9__lane30_strm1_data_valid    ( std__pe9__lane30_strm1_data_valid ),      
               .std__pe9__lane30_strm1_data_mask     ( std__pe9__lane30_strm1_data_mask  ),      

               // PE 9, Lane 31                 
               .pe9__std__lane31_strm0_ready         ( pe9__std__lane31_strm0_ready      ),      
               .std__pe9__lane31_strm0_cntl          ( std__pe9__lane31_strm0_cntl       ),      
               .std__pe9__lane31_strm0_data          ( std__pe9__lane31_strm0_data       ),      
               .std__pe9__lane31_strm0_data_valid    ( std__pe9__lane31_strm0_data_valid ),      
               .std__pe9__lane31_strm0_data_mask     ( std__pe9__lane31_strm0_data_mask  ),      

               .pe9__std__lane31_strm1_ready         ( pe9__std__lane31_strm1_ready      ),      
               .std__pe9__lane31_strm1_cntl          ( std__pe9__lane31_strm1_cntl       ),      
               .std__pe9__lane31_strm1_data          ( std__pe9__lane31_strm1_data       ),      
               .std__pe9__lane31_strm1_data_valid    ( std__pe9__lane31_strm1_data_valid ),      
               .std__pe9__lane31_strm1_data_mask     ( std__pe9__lane31_strm1_data_mask  ),      

               // PE 10, Lane 0                 
               .pe10__std__lane0_strm0_ready         ( pe10__std__lane0_strm0_ready      ),      
               .std__pe10__lane0_strm0_cntl          ( std__pe10__lane0_strm0_cntl       ),      
               .std__pe10__lane0_strm0_data          ( std__pe10__lane0_strm0_data       ),      
               .std__pe10__lane0_strm0_data_valid    ( std__pe10__lane0_strm0_data_valid ),      
               .std__pe10__lane0_strm0_data_mask     ( std__pe10__lane0_strm0_data_mask  ),      

               .pe10__std__lane0_strm1_ready         ( pe10__std__lane0_strm1_ready      ),      
               .std__pe10__lane0_strm1_cntl          ( std__pe10__lane0_strm1_cntl       ),      
               .std__pe10__lane0_strm1_data          ( std__pe10__lane0_strm1_data       ),      
               .std__pe10__lane0_strm1_data_valid    ( std__pe10__lane0_strm1_data_valid ),      
               .std__pe10__lane0_strm1_data_mask     ( std__pe10__lane0_strm1_data_mask  ),      

               // PE 10, Lane 1                 
               .pe10__std__lane1_strm0_ready         ( pe10__std__lane1_strm0_ready      ),      
               .std__pe10__lane1_strm0_cntl          ( std__pe10__lane1_strm0_cntl       ),      
               .std__pe10__lane1_strm0_data          ( std__pe10__lane1_strm0_data       ),      
               .std__pe10__lane1_strm0_data_valid    ( std__pe10__lane1_strm0_data_valid ),      
               .std__pe10__lane1_strm0_data_mask     ( std__pe10__lane1_strm0_data_mask  ),      

               .pe10__std__lane1_strm1_ready         ( pe10__std__lane1_strm1_ready      ),      
               .std__pe10__lane1_strm1_cntl          ( std__pe10__lane1_strm1_cntl       ),      
               .std__pe10__lane1_strm1_data          ( std__pe10__lane1_strm1_data       ),      
               .std__pe10__lane1_strm1_data_valid    ( std__pe10__lane1_strm1_data_valid ),      
               .std__pe10__lane1_strm1_data_mask     ( std__pe10__lane1_strm1_data_mask  ),      

               // PE 10, Lane 2                 
               .pe10__std__lane2_strm0_ready         ( pe10__std__lane2_strm0_ready      ),      
               .std__pe10__lane2_strm0_cntl          ( std__pe10__lane2_strm0_cntl       ),      
               .std__pe10__lane2_strm0_data          ( std__pe10__lane2_strm0_data       ),      
               .std__pe10__lane2_strm0_data_valid    ( std__pe10__lane2_strm0_data_valid ),      
               .std__pe10__lane2_strm0_data_mask     ( std__pe10__lane2_strm0_data_mask  ),      

               .pe10__std__lane2_strm1_ready         ( pe10__std__lane2_strm1_ready      ),      
               .std__pe10__lane2_strm1_cntl          ( std__pe10__lane2_strm1_cntl       ),      
               .std__pe10__lane2_strm1_data          ( std__pe10__lane2_strm1_data       ),      
               .std__pe10__lane2_strm1_data_valid    ( std__pe10__lane2_strm1_data_valid ),      
               .std__pe10__lane2_strm1_data_mask     ( std__pe10__lane2_strm1_data_mask  ),      

               // PE 10, Lane 3                 
               .pe10__std__lane3_strm0_ready         ( pe10__std__lane3_strm0_ready      ),      
               .std__pe10__lane3_strm0_cntl          ( std__pe10__lane3_strm0_cntl       ),      
               .std__pe10__lane3_strm0_data          ( std__pe10__lane3_strm0_data       ),      
               .std__pe10__lane3_strm0_data_valid    ( std__pe10__lane3_strm0_data_valid ),      
               .std__pe10__lane3_strm0_data_mask     ( std__pe10__lane3_strm0_data_mask  ),      

               .pe10__std__lane3_strm1_ready         ( pe10__std__lane3_strm1_ready      ),      
               .std__pe10__lane3_strm1_cntl          ( std__pe10__lane3_strm1_cntl       ),      
               .std__pe10__lane3_strm1_data          ( std__pe10__lane3_strm1_data       ),      
               .std__pe10__lane3_strm1_data_valid    ( std__pe10__lane3_strm1_data_valid ),      
               .std__pe10__lane3_strm1_data_mask     ( std__pe10__lane3_strm1_data_mask  ),      

               // PE 10, Lane 4                 
               .pe10__std__lane4_strm0_ready         ( pe10__std__lane4_strm0_ready      ),      
               .std__pe10__lane4_strm0_cntl          ( std__pe10__lane4_strm0_cntl       ),      
               .std__pe10__lane4_strm0_data          ( std__pe10__lane4_strm0_data       ),      
               .std__pe10__lane4_strm0_data_valid    ( std__pe10__lane4_strm0_data_valid ),      
               .std__pe10__lane4_strm0_data_mask     ( std__pe10__lane4_strm0_data_mask  ),      

               .pe10__std__lane4_strm1_ready         ( pe10__std__lane4_strm1_ready      ),      
               .std__pe10__lane4_strm1_cntl          ( std__pe10__lane4_strm1_cntl       ),      
               .std__pe10__lane4_strm1_data          ( std__pe10__lane4_strm1_data       ),      
               .std__pe10__lane4_strm1_data_valid    ( std__pe10__lane4_strm1_data_valid ),      
               .std__pe10__lane4_strm1_data_mask     ( std__pe10__lane4_strm1_data_mask  ),      

               // PE 10, Lane 5                 
               .pe10__std__lane5_strm0_ready         ( pe10__std__lane5_strm0_ready      ),      
               .std__pe10__lane5_strm0_cntl          ( std__pe10__lane5_strm0_cntl       ),      
               .std__pe10__lane5_strm0_data          ( std__pe10__lane5_strm0_data       ),      
               .std__pe10__lane5_strm0_data_valid    ( std__pe10__lane5_strm0_data_valid ),      
               .std__pe10__lane5_strm0_data_mask     ( std__pe10__lane5_strm0_data_mask  ),      

               .pe10__std__lane5_strm1_ready         ( pe10__std__lane5_strm1_ready      ),      
               .std__pe10__lane5_strm1_cntl          ( std__pe10__lane5_strm1_cntl       ),      
               .std__pe10__lane5_strm1_data          ( std__pe10__lane5_strm1_data       ),      
               .std__pe10__lane5_strm1_data_valid    ( std__pe10__lane5_strm1_data_valid ),      
               .std__pe10__lane5_strm1_data_mask     ( std__pe10__lane5_strm1_data_mask  ),      

               // PE 10, Lane 6                 
               .pe10__std__lane6_strm0_ready         ( pe10__std__lane6_strm0_ready      ),      
               .std__pe10__lane6_strm0_cntl          ( std__pe10__lane6_strm0_cntl       ),      
               .std__pe10__lane6_strm0_data          ( std__pe10__lane6_strm0_data       ),      
               .std__pe10__lane6_strm0_data_valid    ( std__pe10__lane6_strm0_data_valid ),      
               .std__pe10__lane6_strm0_data_mask     ( std__pe10__lane6_strm0_data_mask  ),      

               .pe10__std__lane6_strm1_ready         ( pe10__std__lane6_strm1_ready      ),      
               .std__pe10__lane6_strm1_cntl          ( std__pe10__lane6_strm1_cntl       ),      
               .std__pe10__lane6_strm1_data          ( std__pe10__lane6_strm1_data       ),      
               .std__pe10__lane6_strm1_data_valid    ( std__pe10__lane6_strm1_data_valid ),      
               .std__pe10__lane6_strm1_data_mask     ( std__pe10__lane6_strm1_data_mask  ),      

               // PE 10, Lane 7                 
               .pe10__std__lane7_strm0_ready         ( pe10__std__lane7_strm0_ready      ),      
               .std__pe10__lane7_strm0_cntl          ( std__pe10__lane7_strm0_cntl       ),      
               .std__pe10__lane7_strm0_data          ( std__pe10__lane7_strm0_data       ),      
               .std__pe10__lane7_strm0_data_valid    ( std__pe10__lane7_strm0_data_valid ),      
               .std__pe10__lane7_strm0_data_mask     ( std__pe10__lane7_strm0_data_mask  ),      

               .pe10__std__lane7_strm1_ready         ( pe10__std__lane7_strm1_ready      ),      
               .std__pe10__lane7_strm1_cntl          ( std__pe10__lane7_strm1_cntl       ),      
               .std__pe10__lane7_strm1_data          ( std__pe10__lane7_strm1_data       ),      
               .std__pe10__lane7_strm1_data_valid    ( std__pe10__lane7_strm1_data_valid ),      
               .std__pe10__lane7_strm1_data_mask     ( std__pe10__lane7_strm1_data_mask  ),      

               // PE 10, Lane 8                 
               .pe10__std__lane8_strm0_ready         ( pe10__std__lane8_strm0_ready      ),      
               .std__pe10__lane8_strm0_cntl          ( std__pe10__lane8_strm0_cntl       ),      
               .std__pe10__lane8_strm0_data          ( std__pe10__lane8_strm0_data       ),      
               .std__pe10__lane8_strm0_data_valid    ( std__pe10__lane8_strm0_data_valid ),      
               .std__pe10__lane8_strm0_data_mask     ( std__pe10__lane8_strm0_data_mask  ),      

               .pe10__std__lane8_strm1_ready         ( pe10__std__lane8_strm1_ready      ),      
               .std__pe10__lane8_strm1_cntl          ( std__pe10__lane8_strm1_cntl       ),      
               .std__pe10__lane8_strm1_data          ( std__pe10__lane8_strm1_data       ),      
               .std__pe10__lane8_strm1_data_valid    ( std__pe10__lane8_strm1_data_valid ),      
               .std__pe10__lane8_strm1_data_mask     ( std__pe10__lane8_strm1_data_mask  ),      

               // PE 10, Lane 9                 
               .pe10__std__lane9_strm0_ready         ( pe10__std__lane9_strm0_ready      ),      
               .std__pe10__lane9_strm0_cntl          ( std__pe10__lane9_strm0_cntl       ),      
               .std__pe10__lane9_strm0_data          ( std__pe10__lane9_strm0_data       ),      
               .std__pe10__lane9_strm0_data_valid    ( std__pe10__lane9_strm0_data_valid ),      
               .std__pe10__lane9_strm0_data_mask     ( std__pe10__lane9_strm0_data_mask  ),      

               .pe10__std__lane9_strm1_ready         ( pe10__std__lane9_strm1_ready      ),      
               .std__pe10__lane9_strm1_cntl          ( std__pe10__lane9_strm1_cntl       ),      
               .std__pe10__lane9_strm1_data          ( std__pe10__lane9_strm1_data       ),      
               .std__pe10__lane9_strm1_data_valid    ( std__pe10__lane9_strm1_data_valid ),      
               .std__pe10__lane9_strm1_data_mask     ( std__pe10__lane9_strm1_data_mask  ),      

               // PE 10, Lane 10                 
               .pe10__std__lane10_strm0_ready         ( pe10__std__lane10_strm0_ready      ),      
               .std__pe10__lane10_strm0_cntl          ( std__pe10__lane10_strm0_cntl       ),      
               .std__pe10__lane10_strm0_data          ( std__pe10__lane10_strm0_data       ),      
               .std__pe10__lane10_strm0_data_valid    ( std__pe10__lane10_strm0_data_valid ),      
               .std__pe10__lane10_strm0_data_mask     ( std__pe10__lane10_strm0_data_mask  ),      

               .pe10__std__lane10_strm1_ready         ( pe10__std__lane10_strm1_ready      ),      
               .std__pe10__lane10_strm1_cntl          ( std__pe10__lane10_strm1_cntl       ),      
               .std__pe10__lane10_strm1_data          ( std__pe10__lane10_strm1_data       ),      
               .std__pe10__lane10_strm1_data_valid    ( std__pe10__lane10_strm1_data_valid ),      
               .std__pe10__lane10_strm1_data_mask     ( std__pe10__lane10_strm1_data_mask  ),      

               // PE 10, Lane 11                 
               .pe10__std__lane11_strm0_ready         ( pe10__std__lane11_strm0_ready      ),      
               .std__pe10__lane11_strm0_cntl          ( std__pe10__lane11_strm0_cntl       ),      
               .std__pe10__lane11_strm0_data          ( std__pe10__lane11_strm0_data       ),      
               .std__pe10__lane11_strm0_data_valid    ( std__pe10__lane11_strm0_data_valid ),      
               .std__pe10__lane11_strm0_data_mask     ( std__pe10__lane11_strm0_data_mask  ),      

               .pe10__std__lane11_strm1_ready         ( pe10__std__lane11_strm1_ready      ),      
               .std__pe10__lane11_strm1_cntl          ( std__pe10__lane11_strm1_cntl       ),      
               .std__pe10__lane11_strm1_data          ( std__pe10__lane11_strm1_data       ),      
               .std__pe10__lane11_strm1_data_valid    ( std__pe10__lane11_strm1_data_valid ),      
               .std__pe10__lane11_strm1_data_mask     ( std__pe10__lane11_strm1_data_mask  ),      

               // PE 10, Lane 12                 
               .pe10__std__lane12_strm0_ready         ( pe10__std__lane12_strm0_ready      ),      
               .std__pe10__lane12_strm0_cntl          ( std__pe10__lane12_strm0_cntl       ),      
               .std__pe10__lane12_strm0_data          ( std__pe10__lane12_strm0_data       ),      
               .std__pe10__lane12_strm0_data_valid    ( std__pe10__lane12_strm0_data_valid ),      
               .std__pe10__lane12_strm0_data_mask     ( std__pe10__lane12_strm0_data_mask  ),      

               .pe10__std__lane12_strm1_ready         ( pe10__std__lane12_strm1_ready      ),      
               .std__pe10__lane12_strm1_cntl          ( std__pe10__lane12_strm1_cntl       ),      
               .std__pe10__lane12_strm1_data          ( std__pe10__lane12_strm1_data       ),      
               .std__pe10__lane12_strm1_data_valid    ( std__pe10__lane12_strm1_data_valid ),      
               .std__pe10__lane12_strm1_data_mask     ( std__pe10__lane12_strm1_data_mask  ),      

               // PE 10, Lane 13                 
               .pe10__std__lane13_strm0_ready         ( pe10__std__lane13_strm0_ready      ),      
               .std__pe10__lane13_strm0_cntl          ( std__pe10__lane13_strm0_cntl       ),      
               .std__pe10__lane13_strm0_data          ( std__pe10__lane13_strm0_data       ),      
               .std__pe10__lane13_strm0_data_valid    ( std__pe10__lane13_strm0_data_valid ),      
               .std__pe10__lane13_strm0_data_mask     ( std__pe10__lane13_strm0_data_mask  ),      

               .pe10__std__lane13_strm1_ready         ( pe10__std__lane13_strm1_ready      ),      
               .std__pe10__lane13_strm1_cntl          ( std__pe10__lane13_strm1_cntl       ),      
               .std__pe10__lane13_strm1_data          ( std__pe10__lane13_strm1_data       ),      
               .std__pe10__lane13_strm1_data_valid    ( std__pe10__lane13_strm1_data_valid ),      
               .std__pe10__lane13_strm1_data_mask     ( std__pe10__lane13_strm1_data_mask  ),      

               // PE 10, Lane 14                 
               .pe10__std__lane14_strm0_ready         ( pe10__std__lane14_strm0_ready      ),      
               .std__pe10__lane14_strm0_cntl          ( std__pe10__lane14_strm0_cntl       ),      
               .std__pe10__lane14_strm0_data          ( std__pe10__lane14_strm0_data       ),      
               .std__pe10__lane14_strm0_data_valid    ( std__pe10__lane14_strm0_data_valid ),      
               .std__pe10__lane14_strm0_data_mask     ( std__pe10__lane14_strm0_data_mask  ),      

               .pe10__std__lane14_strm1_ready         ( pe10__std__lane14_strm1_ready      ),      
               .std__pe10__lane14_strm1_cntl          ( std__pe10__lane14_strm1_cntl       ),      
               .std__pe10__lane14_strm1_data          ( std__pe10__lane14_strm1_data       ),      
               .std__pe10__lane14_strm1_data_valid    ( std__pe10__lane14_strm1_data_valid ),      
               .std__pe10__lane14_strm1_data_mask     ( std__pe10__lane14_strm1_data_mask  ),      

               // PE 10, Lane 15                 
               .pe10__std__lane15_strm0_ready         ( pe10__std__lane15_strm0_ready      ),      
               .std__pe10__lane15_strm0_cntl          ( std__pe10__lane15_strm0_cntl       ),      
               .std__pe10__lane15_strm0_data          ( std__pe10__lane15_strm0_data       ),      
               .std__pe10__lane15_strm0_data_valid    ( std__pe10__lane15_strm0_data_valid ),      
               .std__pe10__lane15_strm0_data_mask     ( std__pe10__lane15_strm0_data_mask  ),      

               .pe10__std__lane15_strm1_ready         ( pe10__std__lane15_strm1_ready      ),      
               .std__pe10__lane15_strm1_cntl          ( std__pe10__lane15_strm1_cntl       ),      
               .std__pe10__lane15_strm1_data          ( std__pe10__lane15_strm1_data       ),      
               .std__pe10__lane15_strm1_data_valid    ( std__pe10__lane15_strm1_data_valid ),      
               .std__pe10__lane15_strm1_data_mask     ( std__pe10__lane15_strm1_data_mask  ),      

               // PE 10, Lane 16                 
               .pe10__std__lane16_strm0_ready         ( pe10__std__lane16_strm0_ready      ),      
               .std__pe10__lane16_strm0_cntl          ( std__pe10__lane16_strm0_cntl       ),      
               .std__pe10__lane16_strm0_data          ( std__pe10__lane16_strm0_data       ),      
               .std__pe10__lane16_strm0_data_valid    ( std__pe10__lane16_strm0_data_valid ),      
               .std__pe10__lane16_strm0_data_mask     ( std__pe10__lane16_strm0_data_mask  ),      

               .pe10__std__lane16_strm1_ready         ( pe10__std__lane16_strm1_ready      ),      
               .std__pe10__lane16_strm1_cntl          ( std__pe10__lane16_strm1_cntl       ),      
               .std__pe10__lane16_strm1_data          ( std__pe10__lane16_strm1_data       ),      
               .std__pe10__lane16_strm1_data_valid    ( std__pe10__lane16_strm1_data_valid ),      
               .std__pe10__lane16_strm1_data_mask     ( std__pe10__lane16_strm1_data_mask  ),      

               // PE 10, Lane 17                 
               .pe10__std__lane17_strm0_ready         ( pe10__std__lane17_strm0_ready      ),      
               .std__pe10__lane17_strm0_cntl          ( std__pe10__lane17_strm0_cntl       ),      
               .std__pe10__lane17_strm0_data          ( std__pe10__lane17_strm0_data       ),      
               .std__pe10__lane17_strm0_data_valid    ( std__pe10__lane17_strm0_data_valid ),      
               .std__pe10__lane17_strm0_data_mask     ( std__pe10__lane17_strm0_data_mask  ),      

               .pe10__std__lane17_strm1_ready         ( pe10__std__lane17_strm1_ready      ),      
               .std__pe10__lane17_strm1_cntl          ( std__pe10__lane17_strm1_cntl       ),      
               .std__pe10__lane17_strm1_data          ( std__pe10__lane17_strm1_data       ),      
               .std__pe10__lane17_strm1_data_valid    ( std__pe10__lane17_strm1_data_valid ),      
               .std__pe10__lane17_strm1_data_mask     ( std__pe10__lane17_strm1_data_mask  ),      

               // PE 10, Lane 18                 
               .pe10__std__lane18_strm0_ready         ( pe10__std__lane18_strm0_ready      ),      
               .std__pe10__lane18_strm0_cntl          ( std__pe10__lane18_strm0_cntl       ),      
               .std__pe10__lane18_strm0_data          ( std__pe10__lane18_strm0_data       ),      
               .std__pe10__lane18_strm0_data_valid    ( std__pe10__lane18_strm0_data_valid ),      
               .std__pe10__lane18_strm0_data_mask     ( std__pe10__lane18_strm0_data_mask  ),      

               .pe10__std__lane18_strm1_ready         ( pe10__std__lane18_strm1_ready      ),      
               .std__pe10__lane18_strm1_cntl          ( std__pe10__lane18_strm1_cntl       ),      
               .std__pe10__lane18_strm1_data          ( std__pe10__lane18_strm1_data       ),      
               .std__pe10__lane18_strm1_data_valid    ( std__pe10__lane18_strm1_data_valid ),      
               .std__pe10__lane18_strm1_data_mask     ( std__pe10__lane18_strm1_data_mask  ),      

               // PE 10, Lane 19                 
               .pe10__std__lane19_strm0_ready         ( pe10__std__lane19_strm0_ready      ),      
               .std__pe10__lane19_strm0_cntl          ( std__pe10__lane19_strm0_cntl       ),      
               .std__pe10__lane19_strm0_data          ( std__pe10__lane19_strm0_data       ),      
               .std__pe10__lane19_strm0_data_valid    ( std__pe10__lane19_strm0_data_valid ),      
               .std__pe10__lane19_strm0_data_mask     ( std__pe10__lane19_strm0_data_mask  ),      

               .pe10__std__lane19_strm1_ready         ( pe10__std__lane19_strm1_ready      ),      
               .std__pe10__lane19_strm1_cntl          ( std__pe10__lane19_strm1_cntl       ),      
               .std__pe10__lane19_strm1_data          ( std__pe10__lane19_strm1_data       ),      
               .std__pe10__lane19_strm1_data_valid    ( std__pe10__lane19_strm1_data_valid ),      
               .std__pe10__lane19_strm1_data_mask     ( std__pe10__lane19_strm1_data_mask  ),      

               // PE 10, Lane 20                 
               .pe10__std__lane20_strm0_ready         ( pe10__std__lane20_strm0_ready      ),      
               .std__pe10__lane20_strm0_cntl          ( std__pe10__lane20_strm0_cntl       ),      
               .std__pe10__lane20_strm0_data          ( std__pe10__lane20_strm0_data       ),      
               .std__pe10__lane20_strm0_data_valid    ( std__pe10__lane20_strm0_data_valid ),      
               .std__pe10__lane20_strm0_data_mask     ( std__pe10__lane20_strm0_data_mask  ),      

               .pe10__std__lane20_strm1_ready         ( pe10__std__lane20_strm1_ready      ),      
               .std__pe10__lane20_strm1_cntl          ( std__pe10__lane20_strm1_cntl       ),      
               .std__pe10__lane20_strm1_data          ( std__pe10__lane20_strm1_data       ),      
               .std__pe10__lane20_strm1_data_valid    ( std__pe10__lane20_strm1_data_valid ),      
               .std__pe10__lane20_strm1_data_mask     ( std__pe10__lane20_strm1_data_mask  ),      

               // PE 10, Lane 21                 
               .pe10__std__lane21_strm0_ready         ( pe10__std__lane21_strm0_ready      ),      
               .std__pe10__lane21_strm0_cntl          ( std__pe10__lane21_strm0_cntl       ),      
               .std__pe10__lane21_strm0_data          ( std__pe10__lane21_strm0_data       ),      
               .std__pe10__lane21_strm0_data_valid    ( std__pe10__lane21_strm0_data_valid ),      
               .std__pe10__lane21_strm0_data_mask     ( std__pe10__lane21_strm0_data_mask  ),      

               .pe10__std__lane21_strm1_ready         ( pe10__std__lane21_strm1_ready      ),      
               .std__pe10__lane21_strm1_cntl          ( std__pe10__lane21_strm1_cntl       ),      
               .std__pe10__lane21_strm1_data          ( std__pe10__lane21_strm1_data       ),      
               .std__pe10__lane21_strm1_data_valid    ( std__pe10__lane21_strm1_data_valid ),      
               .std__pe10__lane21_strm1_data_mask     ( std__pe10__lane21_strm1_data_mask  ),      

               // PE 10, Lane 22                 
               .pe10__std__lane22_strm0_ready         ( pe10__std__lane22_strm0_ready      ),      
               .std__pe10__lane22_strm0_cntl          ( std__pe10__lane22_strm0_cntl       ),      
               .std__pe10__lane22_strm0_data          ( std__pe10__lane22_strm0_data       ),      
               .std__pe10__lane22_strm0_data_valid    ( std__pe10__lane22_strm0_data_valid ),      
               .std__pe10__lane22_strm0_data_mask     ( std__pe10__lane22_strm0_data_mask  ),      

               .pe10__std__lane22_strm1_ready         ( pe10__std__lane22_strm1_ready      ),      
               .std__pe10__lane22_strm1_cntl          ( std__pe10__lane22_strm1_cntl       ),      
               .std__pe10__lane22_strm1_data          ( std__pe10__lane22_strm1_data       ),      
               .std__pe10__lane22_strm1_data_valid    ( std__pe10__lane22_strm1_data_valid ),      
               .std__pe10__lane22_strm1_data_mask     ( std__pe10__lane22_strm1_data_mask  ),      

               // PE 10, Lane 23                 
               .pe10__std__lane23_strm0_ready         ( pe10__std__lane23_strm0_ready      ),      
               .std__pe10__lane23_strm0_cntl          ( std__pe10__lane23_strm0_cntl       ),      
               .std__pe10__lane23_strm0_data          ( std__pe10__lane23_strm0_data       ),      
               .std__pe10__lane23_strm0_data_valid    ( std__pe10__lane23_strm0_data_valid ),      
               .std__pe10__lane23_strm0_data_mask     ( std__pe10__lane23_strm0_data_mask  ),      

               .pe10__std__lane23_strm1_ready         ( pe10__std__lane23_strm1_ready      ),      
               .std__pe10__lane23_strm1_cntl          ( std__pe10__lane23_strm1_cntl       ),      
               .std__pe10__lane23_strm1_data          ( std__pe10__lane23_strm1_data       ),      
               .std__pe10__lane23_strm1_data_valid    ( std__pe10__lane23_strm1_data_valid ),      
               .std__pe10__lane23_strm1_data_mask     ( std__pe10__lane23_strm1_data_mask  ),      

               // PE 10, Lane 24                 
               .pe10__std__lane24_strm0_ready         ( pe10__std__lane24_strm0_ready      ),      
               .std__pe10__lane24_strm0_cntl          ( std__pe10__lane24_strm0_cntl       ),      
               .std__pe10__lane24_strm0_data          ( std__pe10__lane24_strm0_data       ),      
               .std__pe10__lane24_strm0_data_valid    ( std__pe10__lane24_strm0_data_valid ),      
               .std__pe10__lane24_strm0_data_mask     ( std__pe10__lane24_strm0_data_mask  ),      

               .pe10__std__lane24_strm1_ready         ( pe10__std__lane24_strm1_ready      ),      
               .std__pe10__lane24_strm1_cntl          ( std__pe10__lane24_strm1_cntl       ),      
               .std__pe10__lane24_strm1_data          ( std__pe10__lane24_strm1_data       ),      
               .std__pe10__lane24_strm1_data_valid    ( std__pe10__lane24_strm1_data_valid ),      
               .std__pe10__lane24_strm1_data_mask     ( std__pe10__lane24_strm1_data_mask  ),      

               // PE 10, Lane 25                 
               .pe10__std__lane25_strm0_ready         ( pe10__std__lane25_strm0_ready      ),      
               .std__pe10__lane25_strm0_cntl          ( std__pe10__lane25_strm0_cntl       ),      
               .std__pe10__lane25_strm0_data          ( std__pe10__lane25_strm0_data       ),      
               .std__pe10__lane25_strm0_data_valid    ( std__pe10__lane25_strm0_data_valid ),      
               .std__pe10__lane25_strm0_data_mask     ( std__pe10__lane25_strm0_data_mask  ),      

               .pe10__std__lane25_strm1_ready         ( pe10__std__lane25_strm1_ready      ),      
               .std__pe10__lane25_strm1_cntl          ( std__pe10__lane25_strm1_cntl       ),      
               .std__pe10__lane25_strm1_data          ( std__pe10__lane25_strm1_data       ),      
               .std__pe10__lane25_strm1_data_valid    ( std__pe10__lane25_strm1_data_valid ),      
               .std__pe10__lane25_strm1_data_mask     ( std__pe10__lane25_strm1_data_mask  ),      

               // PE 10, Lane 26                 
               .pe10__std__lane26_strm0_ready         ( pe10__std__lane26_strm0_ready      ),      
               .std__pe10__lane26_strm0_cntl          ( std__pe10__lane26_strm0_cntl       ),      
               .std__pe10__lane26_strm0_data          ( std__pe10__lane26_strm0_data       ),      
               .std__pe10__lane26_strm0_data_valid    ( std__pe10__lane26_strm0_data_valid ),      
               .std__pe10__lane26_strm0_data_mask     ( std__pe10__lane26_strm0_data_mask  ),      

               .pe10__std__lane26_strm1_ready         ( pe10__std__lane26_strm1_ready      ),      
               .std__pe10__lane26_strm1_cntl          ( std__pe10__lane26_strm1_cntl       ),      
               .std__pe10__lane26_strm1_data          ( std__pe10__lane26_strm1_data       ),      
               .std__pe10__lane26_strm1_data_valid    ( std__pe10__lane26_strm1_data_valid ),      
               .std__pe10__lane26_strm1_data_mask     ( std__pe10__lane26_strm1_data_mask  ),      

               // PE 10, Lane 27                 
               .pe10__std__lane27_strm0_ready         ( pe10__std__lane27_strm0_ready      ),      
               .std__pe10__lane27_strm0_cntl          ( std__pe10__lane27_strm0_cntl       ),      
               .std__pe10__lane27_strm0_data          ( std__pe10__lane27_strm0_data       ),      
               .std__pe10__lane27_strm0_data_valid    ( std__pe10__lane27_strm0_data_valid ),      
               .std__pe10__lane27_strm0_data_mask     ( std__pe10__lane27_strm0_data_mask  ),      

               .pe10__std__lane27_strm1_ready         ( pe10__std__lane27_strm1_ready      ),      
               .std__pe10__lane27_strm1_cntl          ( std__pe10__lane27_strm1_cntl       ),      
               .std__pe10__lane27_strm1_data          ( std__pe10__lane27_strm1_data       ),      
               .std__pe10__lane27_strm1_data_valid    ( std__pe10__lane27_strm1_data_valid ),      
               .std__pe10__lane27_strm1_data_mask     ( std__pe10__lane27_strm1_data_mask  ),      

               // PE 10, Lane 28                 
               .pe10__std__lane28_strm0_ready         ( pe10__std__lane28_strm0_ready      ),      
               .std__pe10__lane28_strm0_cntl          ( std__pe10__lane28_strm0_cntl       ),      
               .std__pe10__lane28_strm0_data          ( std__pe10__lane28_strm0_data       ),      
               .std__pe10__lane28_strm0_data_valid    ( std__pe10__lane28_strm0_data_valid ),      
               .std__pe10__lane28_strm0_data_mask     ( std__pe10__lane28_strm0_data_mask  ),      

               .pe10__std__lane28_strm1_ready         ( pe10__std__lane28_strm1_ready      ),      
               .std__pe10__lane28_strm1_cntl          ( std__pe10__lane28_strm1_cntl       ),      
               .std__pe10__lane28_strm1_data          ( std__pe10__lane28_strm1_data       ),      
               .std__pe10__lane28_strm1_data_valid    ( std__pe10__lane28_strm1_data_valid ),      
               .std__pe10__lane28_strm1_data_mask     ( std__pe10__lane28_strm1_data_mask  ),      

               // PE 10, Lane 29                 
               .pe10__std__lane29_strm0_ready         ( pe10__std__lane29_strm0_ready      ),      
               .std__pe10__lane29_strm0_cntl          ( std__pe10__lane29_strm0_cntl       ),      
               .std__pe10__lane29_strm0_data          ( std__pe10__lane29_strm0_data       ),      
               .std__pe10__lane29_strm0_data_valid    ( std__pe10__lane29_strm0_data_valid ),      
               .std__pe10__lane29_strm0_data_mask     ( std__pe10__lane29_strm0_data_mask  ),      

               .pe10__std__lane29_strm1_ready         ( pe10__std__lane29_strm1_ready      ),      
               .std__pe10__lane29_strm1_cntl          ( std__pe10__lane29_strm1_cntl       ),      
               .std__pe10__lane29_strm1_data          ( std__pe10__lane29_strm1_data       ),      
               .std__pe10__lane29_strm1_data_valid    ( std__pe10__lane29_strm1_data_valid ),      
               .std__pe10__lane29_strm1_data_mask     ( std__pe10__lane29_strm1_data_mask  ),      

               // PE 10, Lane 30                 
               .pe10__std__lane30_strm0_ready         ( pe10__std__lane30_strm0_ready      ),      
               .std__pe10__lane30_strm0_cntl          ( std__pe10__lane30_strm0_cntl       ),      
               .std__pe10__lane30_strm0_data          ( std__pe10__lane30_strm0_data       ),      
               .std__pe10__lane30_strm0_data_valid    ( std__pe10__lane30_strm0_data_valid ),      
               .std__pe10__lane30_strm0_data_mask     ( std__pe10__lane30_strm0_data_mask  ),      

               .pe10__std__lane30_strm1_ready         ( pe10__std__lane30_strm1_ready      ),      
               .std__pe10__lane30_strm1_cntl          ( std__pe10__lane30_strm1_cntl       ),      
               .std__pe10__lane30_strm1_data          ( std__pe10__lane30_strm1_data       ),      
               .std__pe10__lane30_strm1_data_valid    ( std__pe10__lane30_strm1_data_valid ),      
               .std__pe10__lane30_strm1_data_mask     ( std__pe10__lane30_strm1_data_mask  ),      

               // PE 10, Lane 31                 
               .pe10__std__lane31_strm0_ready         ( pe10__std__lane31_strm0_ready      ),      
               .std__pe10__lane31_strm0_cntl          ( std__pe10__lane31_strm0_cntl       ),      
               .std__pe10__lane31_strm0_data          ( std__pe10__lane31_strm0_data       ),      
               .std__pe10__lane31_strm0_data_valid    ( std__pe10__lane31_strm0_data_valid ),      
               .std__pe10__lane31_strm0_data_mask     ( std__pe10__lane31_strm0_data_mask  ),      

               .pe10__std__lane31_strm1_ready         ( pe10__std__lane31_strm1_ready      ),      
               .std__pe10__lane31_strm1_cntl          ( std__pe10__lane31_strm1_cntl       ),      
               .std__pe10__lane31_strm1_data          ( std__pe10__lane31_strm1_data       ),      
               .std__pe10__lane31_strm1_data_valid    ( std__pe10__lane31_strm1_data_valid ),      
               .std__pe10__lane31_strm1_data_mask     ( std__pe10__lane31_strm1_data_mask  ),      

               // PE 11, Lane 0                 
               .pe11__std__lane0_strm0_ready         ( pe11__std__lane0_strm0_ready      ),      
               .std__pe11__lane0_strm0_cntl          ( std__pe11__lane0_strm0_cntl       ),      
               .std__pe11__lane0_strm0_data          ( std__pe11__lane0_strm0_data       ),      
               .std__pe11__lane0_strm0_data_valid    ( std__pe11__lane0_strm0_data_valid ),      
               .std__pe11__lane0_strm0_data_mask     ( std__pe11__lane0_strm0_data_mask  ),      

               .pe11__std__lane0_strm1_ready         ( pe11__std__lane0_strm1_ready      ),      
               .std__pe11__lane0_strm1_cntl          ( std__pe11__lane0_strm1_cntl       ),      
               .std__pe11__lane0_strm1_data          ( std__pe11__lane0_strm1_data       ),      
               .std__pe11__lane0_strm1_data_valid    ( std__pe11__lane0_strm1_data_valid ),      
               .std__pe11__lane0_strm1_data_mask     ( std__pe11__lane0_strm1_data_mask  ),      

               // PE 11, Lane 1                 
               .pe11__std__lane1_strm0_ready         ( pe11__std__lane1_strm0_ready      ),      
               .std__pe11__lane1_strm0_cntl          ( std__pe11__lane1_strm0_cntl       ),      
               .std__pe11__lane1_strm0_data          ( std__pe11__lane1_strm0_data       ),      
               .std__pe11__lane1_strm0_data_valid    ( std__pe11__lane1_strm0_data_valid ),      
               .std__pe11__lane1_strm0_data_mask     ( std__pe11__lane1_strm0_data_mask  ),      

               .pe11__std__lane1_strm1_ready         ( pe11__std__lane1_strm1_ready      ),      
               .std__pe11__lane1_strm1_cntl          ( std__pe11__lane1_strm1_cntl       ),      
               .std__pe11__lane1_strm1_data          ( std__pe11__lane1_strm1_data       ),      
               .std__pe11__lane1_strm1_data_valid    ( std__pe11__lane1_strm1_data_valid ),      
               .std__pe11__lane1_strm1_data_mask     ( std__pe11__lane1_strm1_data_mask  ),      

               // PE 11, Lane 2                 
               .pe11__std__lane2_strm0_ready         ( pe11__std__lane2_strm0_ready      ),      
               .std__pe11__lane2_strm0_cntl          ( std__pe11__lane2_strm0_cntl       ),      
               .std__pe11__lane2_strm0_data          ( std__pe11__lane2_strm0_data       ),      
               .std__pe11__lane2_strm0_data_valid    ( std__pe11__lane2_strm0_data_valid ),      
               .std__pe11__lane2_strm0_data_mask     ( std__pe11__lane2_strm0_data_mask  ),      

               .pe11__std__lane2_strm1_ready         ( pe11__std__lane2_strm1_ready      ),      
               .std__pe11__lane2_strm1_cntl          ( std__pe11__lane2_strm1_cntl       ),      
               .std__pe11__lane2_strm1_data          ( std__pe11__lane2_strm1_data       ),      
               .std__pe11__lane2_strm1_data_valid    ( std__pe11__lane2_strm1_data_valid ),      
               .std__pe11__lane2_strm1_data_mask     ( std__pe11__lane2_strm1_data_mask  ),      

               // PE 11, Lane 3                 
               .pe11__std__lane3_strm0_ready         ( pe11__std__lane3_strm0_ready      ),      
               .std__pe11__lane3_strm0_cntl          ( std__pe11__lane3_strm0_cntl       ),      
               .std__pe11__lane3_strm0_data          ( std__pe11__lane3_strm0_data       ),      
               .std__pe11__lane3_strm0_data_valid    ( std__pe11__lane3_strm0_data_valid ),      
               .std__pe11__lane3_strm0_data_mask     ( std__pe11__lane3_strm0_data_mask  ),      

               .pe11__std__lane3_strm1_ready         ( pe11__std__lane3_strm1_ready      ),      
               .std__pe11__lane3_strm1_cntl          ( std__pe11__lane3_strm1_cntl       ),      
               .std__pe11__lane3_strm1_data          ( std__pe11__lane3_strm1_data       ),      
               .std__pe11__lane3_strm1_data_valid    ( std__pe11__lane3_strm1_data_valid ),      
               .std__pe11__lane3_strm1_data_mask     ( std__pe11__lane3_strm1_data_mask  ),      

               // PE 11, Lane 4                 
               .pe11__std__lane4_strm0_ready         ( pe11__std__lane4_strm0_ready      ),      
               .std__pe11__lane4_strm0_cntl          ( std__pe11__lane4_strm0_cntl       ),      
               .std__pe11__lane4_strm0_data          ( std__pe11__lane4_strm0_data       ),      
               .std__pe11__lane4_strm0_data_valid    ( std__pe11__lane4_strm0_data_valid ),      
               .std__pe11__lane4_strm0_data_mask     ( std__pe11__lane4_strm0_data_mask  ),      

               .pe11__std__lane4_strm1_ready         ( pe11__std__lane4_strm1_ready      ),      
               .std__pe11__lane4_strm1_cntl          ( std__pe11__lane4_strm1_cntl       ),      
               .std__pe11__lane4_strm1_data          ( std__pe11__lane4_strm1_data       ),      
               .std__pe11__lane4_strm1_data_valid    ( std__pe11__lane4_strm1_data_valid ),      
               .std__pe11__lane4_strm1_data_mask     ( std__pe11__lane4_strm1_data_mask  ),      

               // PE 11, Lane 5                 
               .pe11__std__lane5_strm0_ready         ( pe11__std__lane5_strm0_ready      ),      
               .std__pe11__lane5_strm0_cntl          ( std__pe11__lane5_strm0_cntl       ),      
               .std__pe11__lane5_strm0_data          ( std__pe11__lane5_strm0_data       ),      
               .std__pe11__lane5_strm0_data_valid    ( std__pe11__lane5_strm0_data_valid ),      
               .std__pe11__lane5_strm0_data_mask     ( std__pe11__lane5_strm0_data_mask  ),      

               .pe11__std__lane5_strm1_ready         ( pe11__std__lane5_strm1_ready      ),      
               .std__pe11__lane5_strm1_cntl          ( std__pe11__lane5_strm1_cntl       ),      
               .std__pe11__lane5_strm1_data          ( std__pe11__lane5_strm1_data       ),      
               .std__pe11__lane5_strm1_data_valid    ( std__pe11__lane5_strm1_data_valid ),      
               .std__pe11__lane5_strm1_data_mask     ( std__pe11__lane5_strm1_data_mask  ),      

               // PE 11, Lane 6                 
               .pe11__std__lane6_strm0_ready         ( pe11__std__lane6_strm0_ready      ),      
               .std__pe11__lane6_strm0_cntl          ( std__pe11__lane6_strm0_cntl       ),      
               .std__pe11__lane6_strm0_data          ( std__pe11__lane6_strm0_data       ),      
               .std__pe11__lane6_strm0_data_valid    ( std__pe11__lane6_strm0_data_valid ),      
               .std__pe11__lane6_strm0_data_mask     ( std__pe11__lane6_strm0_data_mask  ),      

               .pe11__std__lane6_strm1_ready         ( pe11__std__lane6_strm1_ready      ),      
               .std__pe11__lane6_strm1_cntl          ( std__pe11__lane6_strm1_cntl       ),      
               .std__pe11__lane6_strm1_data          ( std__pe11__lane6_strm1_data       ),      
               .std__pe11__lane6_strm1_data_valid    ( std__pe11__lane6_strm1_data_valid ),      
               .std__pe11__lane6_strm1_data_mask     ( std__pe11__lane6_strm1_data_mask  ),      

               // PE 11, Lane 7                 
               .pe11__std__lane7_strm0_ready         ( pe11__std__lane7_strm0_ready      ),      
               .std__pe11__lane7_strm0_cntl          ( std__pe11__lane7_strm0_cntl       ),      
               .std__pe11__lane7_strm0_data          ( std__pe11__lane7_strm0_data       ),      
               .std__pe11__lane7_strm0_data_valid    ( std__pe11__lane7_strm0_data_valid ),      
               .std__pe11__lane7_strm0_data_mask     ( std__pe11__lane7_strm0_data_mask  ),      

               .pe11__std__lane7_strm1_ready         ( pe11__std__lane7_strm1_ready      ),      
               .std__pe11__lane7_strm1_cntl          ( std__pe11__lane7_strm1_cntl       ),      
               .std__pe11__lane7_strm1_data          ( std__pe11__lane7_strm1_data       ),      
               .std__pe11__lane7_strm1_data_valid    ( std__pe11__lane7_strm1_data_valid ),      
               .std__pe11__lane7_strm1_data_mask     ( std__pe11__lane7_strm1_data_mask  ),      

               // PE 11, Lane 8                 
               .pe11__std__lane8_strm0_ready         ( pe11__std__lane8_strm0_ready      ),      
               .std__pe11__lane8_strm0_cntl          ( std__pe11__lane8_strm0_cntl       ),      
               .std__pe11__lane8_strm0_data          ( std__pe11__lane8_strm0_data       ),      
               .std__pe11__lane8_strm0_data_valid    ( std__pe11__lane8_strm0_data_valid ),      
               .std__pe11__lane8_strm0_data_mask     ( std__pe11__lane8_strm0_data_mask  ),      

               .pe11__std__lane8_strm1_ready         ( pe11__std__lane8_strm1_ready      ),      
               .std__pe11__lane8_strm1_cntl          ( std__pe11__lane8_strm1_cntl       ),      
               .std__pe11__lane8_strm1_data          ( std__pe11__lane8_strm1_data       ),      
               .std__pe11__lane8_strm1_data_valid    ( std__pe11__lane8_strm1_data_valid ),      
               .std__pe11__lane8_strm1_data_mask     ( std__pe11__lane8_strm1_data_mask  ),      

               // PE 11, Lane 9                 
               .pe11__std__lane9_strm0_ready         ( pe11__std__lane9_strm0_ready      ),      
               .std__pe11__lane9_strm0_cntl          ( std__pe11__lane9_strm0_cntl       ),      
               .std__pe11__lane9_strm0_data          ( std__pe11__lane9_strm0_data       ),      
               .std__pe11__lane9_strm0_data_valid    ( std__pe11__lane9_strm0_data_valid ),      
               .std__pe11__lane9_strm0_data_mask     ( std__pe11__lane9_strm0_data_mask  ),      

               .pe11__std__lane9_strm1_ready         ( pe11__std__lane9_strm1_ready      ),      
               .std__pe11__lane9_strm1_cntl          ( std__pe11__lane9_strm1_cntl       ),      
               .std__pe11__lane9_strm1_data          ( std__pe11__lane9_strm1_data       ),      
               .std__pe11__lane9_strm1_data_valid    ( std__pe11__lane9_strm1_data_valid ),      
               .std__pe11__lane9_strm1_data_mask     ( std__pe11__lane9_strm1_data_mask  ),      

               // PE 11, Lane 10                 
               .pe11__std__lane10_strm0_ready         ( pe11__std__lane10_strm0_ready      ),      
               .std__pe11__lane10_strm0_cntl          ( std__pe11__lane10_strm0_cntl       ),      
               .std__pe11__lane10_strm0_data          ( std__pe11__lane10_strm0_data       ),      
               .std__pe11__lane10_strm0_data_valid    ( std__pe11__lane10_strm0_data_valid ),      
               .std__pe11__lane10_strm0_data_mask     ( std__pe11__lane10_strm0_data_mask  ),      

               .pe11__std__lane10_strm1_ready         ( pe11__std__lane10_strm1_ready      ),      
               .std__pe11__lane10_strm1_cntl          ( std__pe11__lane10_strm1_cntl       ),      
               .std__pe11__lane10_strm1_data          ( std__pe11__lane10_strm1_data       ),      
               .std__pe11__lane10_strm1_data_valid    ( std__pe11__lane10_strm1_data_valid ),      
               .std__pe11__lane10_strm1_data_mask     ( std__pe11__lane10_strm1_data_mask  ),      

               // PE 11, Lane 11                 
               .pe11__std__lane11_strm0_ready         ( pe11__std__lane11_strm0_ready      ),      
               .std__pe11__lane11_strm0_cntl          ( std__pe11__lane11_strm0_cntl       ),      
               .std__pe11__lane11_strm0_data          ( std__pe11__lane11_strm0_data       ),      
               .std__pe11__lane11_strm0_data_valid    ( std__pe11__lane11_strm0_data_valid ),      
               .std__pe11__lane11_strm0_data_mask     ( std__pe11__lane11_strm0_data_mask  ),      

               .pe11__std__lane11_strm1_ready         ( pe11__std__lane11_strm1_ready      ),      
               .std__pe11__lane11_strm1_cntl          ( std__pe11__lane11_strm1_cntl       ),      
               .std__pe11__lane11_strm1_data          ( std__pe11__lane11_strm1_data       ),      
               .std__pe11__lane11_strm1_data_valid    ( std__pe11__lane11_strm1_data_valid ),      
               .std__pe11__lane11_strm1_data_mask     ( std__pe11__lane11_strm1_data_mask  ),      

               // PE 11, Lane 12                 
               .pe11__std__lane12_strm0_ready         ( pe11__std__lane12_strm0_ready      ),      
               .std__pe11__lane12_strm0_cntl          ( std__pe11__lane12_strm0_cntl       ),      
               .std__pe11__lane12_strm0_data          ( std__pe11__lane12_strm0_data       ),      
               .std__pe11__lane12_strm0_data_valid    ( std__pe11__lane12_strm0_data_valid ),      
               .std__pe11__lane12_strm0_data_mask     ( std__pe11__lane12_strm0_data_mask  ),      

               .pe11__std__lane12_strm1_ready         ( pe11__std__lane12_strm1_ready      ),      
               .std__pe11__lane12_strm1_cntl          ( std__pe11__lane12_strm1_cntl       ),      
               .std__pe11__lane12_strm1_data          ( std__pe11__lane12_strm1_data       ),      
               .std__pe11__lane12_strm1_data_valid    ( std__pe11__lane12_strm1_data_valid ),      
               .std__pe11__lane12_strm1_data_mask     ( std__pe11__lane12_strm1_data_mask  ),      

               // PE 11, Lane 13                 
               .pe11__std__lane13_strm0_ready         ( pe11__std__lane13_strm0_ready      ),      
               .std__pe11__lane13_strm0_cntl          ( std__pe11__lane13_strm0_cntl       ),      
               .std__pe11__lane13_strm0_data          ( std__pe11__lane13_strm0_data       ),      
               .std__pe11__lane13_strm0_data_valid    ( std__pe11__lane13_strm0_data_valid ),      
               .std__pe11__lane13_strm0_data_mask     ( std__pe11__lane13_strm0_data_mask  ),      

               .pe11__std__lane13_strm1_ready         ( pe11__std__lane13_strm1_ready      ),      
               .std__pe11__lane13_strm1_cntl          ( std__pe11__lane13_strm1_cntl       ),      
               .std__pe11__lane13_strm1_data          ( std__pe11__lane13_strm1_data       ),      
               .std__pe11__lane13_strm1_data_valid    ( std__pe11__lane13_strm1_data_valid ),      
               .std__pe11__lane13_strm1_data_mask     ( std__pe11__lane13_strm1_data_mask  ),      

               // PE 11, Lane 14                 
               .pe11__std__lane14_strm0_ready         ( pe11__std__lane14_strm0_ready      ),      
               .std__pe11__lane14_strm0_cntl          ( std__pe11__lane14_strm0_cntl       ),      
               .std__pe11__lane14_strm0_data          ( std__pe11__lane14_strm0_data       ),      
               .std__pe11__lane14_strm0_data_valid    ( std__pe11__lane14_strm0_data_valid ),      
               .std__pe11__lane14_strm0_data_mask     ( std__pe11__lane14_strm0_data_mask  ),      

               .pe11__std__lane14_strm1_ready         ( pe11__std__lane14_strm1_ready      ),      
               .std__pe11__lane14_strm1_cntl          ( std__pe11__lane14_strm1_cntl       ),      
               .std__pe11__lane14_strm1_data          ( std__pe11__lane14_strm1_data       ),      
               .std__pe11__lane14_strm1_data_valid    ( std__pe11__lane14_strm1_data_valid ),      
               .std__pe11__lane14_strm1_data_mask     ( std__pe11__lane14_strm1_data_mask  ),      

               // PE 11, Lane 15                 
               .pe11__std__lane15_strm0_ready         ( pe11__std__lane15_strm0_ready      ),      
               .std__pe11__lane15_strm0_cntl          ( std__pe11__lane15_strm0_cntl       ),      
               .std__pe11__lane15_strm0_data          ( std__pe11__lane15_strm0_data       ),      
               .std__pe11__lane15_strm0_data_valid    ( std__pe11__lane15_strm0_data_valid ),      
               .std__pe11__lane15_strm0_data_mask     ( std__pe11__lane15_strm0_data_mask  ),      

               .pe11__std__lane15_strm1_ready         ( pe11__std__lane15_strm1_ready      ),      
               .std__pe11__lane15_strm1_cntl          ( std__pe11__lane15_strm1_cntl       ),      
               .std__pe11__lane15_strm1_data          ( std__pe11__lane15_strm1_data       ),      
               .std__pe11__lane15_strm1_data_valid    ( std__pe11__lane15_strm1_data_valid ),      
               .std__pe11__lane15_strm1_data_mask     ( std__pe11__lane15_strm1_data_mask  ),      

               // PE 11, Lane 16                 
               .pe11__std__lane16_strm0_ready         ( pe11__std__lane16_strm0_ready      ),      
               .std__pe11__lane16_strm0_cntl          ( std__pe11__lane16_strm0_cntl       ),      
               .std__pe11__lane16_strm0_data          ( std__pe11__lane16_strm0_data       ),      
               .std__pe11__lane16_strm0_data_valid    ( std__pe11__lane16_strm0_data_valid ),      
               .std__pe11__lane16_strm0_data_mask     ( std__pe11__lane16_strm0_data_mask  ),      

               .pe11__std__lane16_strm1_ready         ( pe11__std__lane16_strm1_ready      ),      
               .std__pe11__lane16_strm1_cntl          ( std__pe11__lane16_strm1_cntl       ),      
               .std__pe11__lane16_strm1_data          ( std__pe11__lane16_strm1_data       ),      
               .std__pe11__lane16_strm1_data_valid    ( std__pe11__lane16_strm1_data_valid ),      
               .std__pe11__lane16_strm1_data_mask     ( std__pe11__lane16_strm1_data_mask  ),      

               // PE 11, Lane 17                 
               .pe11__std__lane17_strm0_ready         ( pe11__std__lane17_strm0_ready      ),      
               .std__pe11__lane17_strm0_cntl          ( std__pe11__lane17_strm0_cntl       ),      
               .std__pe11__lane17_strm0_data          ( std__pe11__lane17_strm0_data       ),      
               .std__pe11__lane17_strm0_data_valid    ( std__pe11__lane17_strm0_data_valid ),      
               .std__pe11__lane17_strm0_data_mask     ( std__pe11__lane17_strm0_data_mask  ),      

               .pe11__std__lane17_strm1_ready         ( pe11__std__lane17_strm1_ready      ),      
               .std__pe11__lane17_strm1_cntl          ( std__pe11__lane17_strm1_cntl       ),      
               .std__pe11__lane17_strm1_data          ( std__pe11__lane17_strm1_data       ),      
               .std__pe11__lane17_strm1_data_valid    ( std__pe11__lane17_strm1_data_valid ),      
               .std__pe11__lane17_strm1_data_mask     ( std__pe11__lane17_strm1_data_mask  ),      

               // PE 11, Lane 18                 
               .pe11__std__lane18_strm0_ready         ( pe11__std__lane18_strm0_ready      ),      
               .std__pe11__lane18_strm0_cntl          ( std__pe11__lane18_strm0_cntl       ),      
               .std__pe11__lane18_strm0_data          ( std__pe11__lane18_strm0_data       ),      
               .std__pe11__lane18_strm0_data_valid    ( std__pe11__lane18_strm0_data_valid ),      
               .std__pe11__lane18_strm0_data_mask     ( std__pe11__lane18_strm0_data_mask  ),      

               .pe11__std__lane18_strm1_ready         ( pe11__std__lane18_strm1_ready      ),      
               .std__pe11__lane18_strm1_cntl          ( std__pe11__lane18_strm1_cntl       ),      
               .std__pe11__lane18_strm1_data          ( std__pe11__lane18_strm1_data       ),      
               .std__pe11__lane18_strm1_data_valid    ( std__pe11__lane18_strm1_data_valid ),      
               .std__pe11__lane18_strm1_data_mask     ( std__pe11__lane18_strm1_data_mask  ),      

               // PE 11, Lane 19                 
               .pe11__std__lane19_strm0_ready         ( pe11__std__lane19_strm0_ready      ),      
               .std__pe11__lane19_strm0_cntl          ( std__pe11__lane19_strm0_cntl       ),      
               .std__pe11__lane19_strm0_data          ( std__pe11__lane19_strm0_data       ),      
               .std__pe11__lane19_strm0_data_valid    ( std__pe11__lane19_strm0_data_valid ),      
               .std__pe11__lane19_strm0_data_mask     ( std__pe11__lane19_strm0_data_mask  ),      

               .pe11__std__lane19_strm1_ready         ( pe11__std__lane19_strm1_ready      ),      
               .std__pe11__lane19_strm1_cntl          ( std__pe11__lane19_strm1_cntl       ),      
               .std__pe11__lane19_strm1_data          ( std__pe11__lane19_strm1_data       ),      
               .std__pe11__lane19_strm1_data_valid    ( std__pe11__lane19_strm1_data_valid ),      
               .std__pe11__lane19_strm1_data_mask     ( std__pe11__lane19_strm1_data_mask  ),      

               // PE 11, Lane 20                 
               .pe11__std__lane20_strm0_ready         ( pe11__std__lane20_strm0_ready      ),      
               .std__pe11__lane20_strm0_cntl          ( std__pe11__lane20_strm0_cntl       ),      
               .std__pe11__lane20_strm0_data          ( std__pe11__lane20_strm0_data       ),      
               .std__pe11__lane20_strm0_data_valid    ( std__pe11__lane20_strm0_data_valid ),      
               .std__pe11__lane20_strm0_data_mask     ( std__pe11__lane20_strm0_data_mask  ),      

               .pe11__std__lane20_strm1_ready         ( pe11__std__lane20_strm1_ready      ),      
               .std__pe11__lane20_strm1_cntl          ( std__pe11__lane20_strm1_cntl       ),      
               .std__pe11__lane20_strm1_data          ( std__pe11__lane20_strm1_data       ),      
               .std__pe11__lane20_strm1_data_valid    ( std__pe11__lane20_strm1_data_valid ),      
               .std__pe11__lane20_strm1_data_mask     ( std__pe11__lane20_strm1_data_mask  ),      

               // PE 11, Lane 21                 
               .pe11__std__lane21_strm0_ready         ( pe11__std__lane21_strm0_ready      ),      
               .std__pe11__lane21_strm0_cntl          ( std__pe11__lane21_strm0_cntl       ),      
               .std__pe11__lane21_strm0_data          ( std__pe11__lane21_strm0_data       ),      
               .std__pe11__lane21_strm0_data_valid    ( std__pe11__lane21_strm0_data_valid ),      
               .std__pe11__lane21_strm0_data_mask     ( std__pe11__lane21_strm0_data_mask  ),      

               .pe11__std__lane21_strm1_ready         ( pe11__std__lane21_strm1_ready      ),      
               .std__pe11__lane21_strm1_cntl          ( std__pe11__lane21_strm1_cntl       ),      
               .std__pe11__lane21_strm1_data          ( std__pe11__lane21_strm1_data       ),      
               .std__pe11__lane21_strm1_data_valid    ( std__pe11__lane21_strm1_data_valid ),      
               .std__pe11__lane21_strm1_data_mask     ( std__pe11__lane21_strm1_data_mask  ),      

               // PE 11, Lane 22                 
               .pe11__std__lane22_strm0_ready         ( pe11__std__lane22_strm0_ready      ),      
               .std__pe11__lane22_strm0_cntl          ( std__pe11__lane22_strm0_cntl       ),      
               .std__pe11__lane22_strm0_data          ( std__pe11__lane22_strm0_data       ),      
               .std__pe11__lane22_strm0_data_valid    ( std__pe11__lane22_strm0_data_valid ),      
               .std__pe11__lane22_strm0_data_mask     ( std__pe11__lane22_strm0_data_mask  ),      

               .pe11__std__lane22_strm1_ready         ( pe11__std__lane22_strm1_ready      ),      
               .std__pe11__lane22_strm1_cntl          ( std__pe11__lane22_strm1_cntl       ),      
               .std__pe11__lane22_strm1_data          ( std__pe11__lane22_strm1_data       ),      
               .std__pe11__lane22_strm1_data_valid    ( std__pe11__lane22_strm1_data_valid ),      
               .std__pe11__lane22_strm1_data_mask     ( std__pe11__lane22_strm1_data_mask  ),      

               // PE 11, Lane 23                 
               .pe11__std__lane23_strm0_ready         ( pe11__std__lane23_strm0_ready      ),      
               .std__pe11__lane23_strm0_cntl          ( std__pe11__lane23_strm0_cntl       ),      
               .std__pe11__lane23_strm0_data          ( std__pe11__lane23_strm0_data       ),      
               .std__pe11__lane23_strm0_data_valid    ( std__pe11__lane23_strm0_data_valid ),      
               .std__pe11__lane23_strm0_data_mask     ( std__pe11__lane23_strm0_data_mask  ),      

               .pe11__std__lane23_strm1_ready         ( pe11__std__lane23_strm1_ready      ),      
               .std__pe11__lane23_strm1_cntl          ( std__pe11__lane23_strm1_cntl       ),      
               .std__pe11__lane23_strm1_data          ( std__pe11__lane23_strm1_data       ),      
               .std__pe11__lane23_strm1_data_valid    ( std__pe11__lane23_strm1_data_valid ),      
               .std__pe11__lane23_strm1_data_mask     ( std__pe11__lane23_strm1_data_mask  ),      

               // PE 11, Lane 24                 
               .pe11__std__lane24_strm0_ready         ( pe11__std__lane24_strm0_ready      ),      
               .std__pe11__lane24_strm0_cntl          ( std__pe11__lane24_strm0_cntl       ),      
               .std__pe11__lane24_strm0_data          ( std__pe11__lane24_strm0_data       ),      
               .std__pe11__lane24_strm0_data_valid    ( std__pe11__lane24_strm0_data_valid ),      
               .std__pe11__lane24_strm0_data_mask     ( std__pe11__lane24_strm0_data_mask  ),      

               .pe11__std__lane24_strm1_ready         ( pe11__std__lane24_strm1_ready      ),      
               .std__pe11__lane24_strm1_cntl          ( std__pe11__lane24_strm1_cntl       ),      
               .std__pe11__lane24_strm1_data          ( std__pe11__lane24_strm1_data       ),      
               .std__pe11__lane24_strm1_data_valid    ( std__pe11__lane24_strm1_data_valid ),      
               .std__pe11__lane24_strm1_data_mask     ( std__pe11__lane24_strm1_data_mask  ),      

               // PE 11, Lane 25                 
               .pe11__std__lane25_strm0_ready         ( pe11__std__lane25_strm0_ready      ),      
               .std__pe11__lane25_strm0_cntl          ( std__pe11__lane25_strm0_cntl       ),      
               .std__pe11__lane25_strm0_data          ( std__pe11__lane25_strm0_data       ),      
               .std__pe11__lane25_strm0_data_valid    ( std__pe11__lane25_strm0_data_valid ),      
               .std__pe11__lane25_strm0_data_mask     ( std__pe11__lane25_strm0_data_mask  ),      

               .pe11__std__lane25_strm1_ready         ( pe11__std__lane25_strm1_ready      ),      
               .std__pe11__lane25_strm1_cntl          ( std__pe11__lane25_strm1_cntl       ),      
               .std__pe11__lane25_strm1_data          ( std__pe11__lane25_strm1_data       ),      
               .std__pe11__lane25_strm1_data_valid    ( std__pe11__lane25_strm1_data_valid ),      
               .std__pe11__lane25_strm1_data_mask     ( std__pe11__lane25_strm1_data_mask  ),      

               // PE 11, Lane 26                 
               .pe11__std__lane26_strm0_ready         ( pe11__std__lane26_strm0_ready      ),      
               .std__pe11__lane26_strm0_cntl          ( std__pe11__lane26_strm0_cntl       ),      
               .std__pe11__lane26_strm0_data          ( std__pe11__lane26_strm0_data       ),      
               .std__pe11__lane26_strm0_data_valid    ( std__pe11__lane26_strm0_data_valid ),      
               .std__pe11__lane26_strm0_data_mask     ( std__pe11__lane26_strm0_data_mask  ),      

               .pe11__std__lane26_strm1_ready         ( pe11__std__lane26_strm1_ready      ),      
               .std__pe11__lane26_strm1_cntl          ( std__pe11__lane26_strm1_cntl       ),      
               .std__pe11__lane26_strm1_data          ( std__pe11__lane26_strm1_data       ),      
               .std__pe11__lane26_strm1_data_valid    ( std__pe11__lane26_strm1_data_valid ),      
               .std__pe11__lane26_strm1_data_mask     ( std__pe11__lane26_strm1_data_mask  ),      

               // PE 11, Lane 27                 
               .pe11__std__lane27_strm0_ready         ( pe11__std__lane27_strm0_ready      ),      
               .std__pe11__lane27_strm0_cntl          ( std__pe11__lane27_strm0_cntl       ),      
               .std__pe11__lane27_strm0_data          ( std__pe11__lane27_strm0_data       ),      
               .std__pe11__lane27_strm0_data_valid    ( std__pe11__lane27_strm0_data_valid ),      
               .std__pe11__lane27_strm0_data_mask     ( std__pe11__lane27_strm0_data_mask  ),      

               .pe11__std__lane27_strm1_ready         ( pe11__std__lane27_strm1_ready      ),      
               .std__pe11__lane27_strm1_cntl          ( std__pe11__lane27_strm1_cntl       ),      
               .std__pe11__lane27_strm1_data          ( std__pe11__lane27_strm1_data       ),      
               .std__pe11__lane27_strm1_data_valid    ( std__pe11__lane27_strm1_data_valid ),      
               .std__pe11__lane27_strm1_data_mask     ( std__pe11__lane27_strm1_data_mask  ),      

               // PE 11, Lane 28                 
               .pe11__std__lane28_strm0_ready         ( pe11__std__lane28_strm0_ready      ),      
               .std__pe11__lane28_strm0_cntl          ( std__pe11__lane28_strm0_cntl       ),      
               .std__pe11__lane28_strm0_data          ( std__pe11__lane28_strm0_data       ),      
               .std__pe11__lane28_strm0_data_valid    ( std__pe11__lane28_strm0_data_valid ),      
               .std__pe11__lane28_strm0_data_mask     ( std__pe11__lane28_strm0_data_mask  ),      

               .pe11__std__lane28_strm1_ready         ( pe11__std__lane28_strm1_ready      ),      
               .std__pe11__lane28_strm1_cntl          ( std__pe11__lane28_strm1_cntl       ),      
               .std__pe11__lane28_strm1_data          ( std__pe11__lane28_strm1_data       ),      
               .std__pe11__lane28_strm1_data_valid    ( std__pe11__lane28_strm1_data_valid ),      
               .std__pe11__lane28_strm1_data_mask     ( std__pe11__lane28_strm1_data_mask  ),      

               // PE 11, Lane 29                 
               .pe11__std__lane29_strm0_ready         ( pe11__std__lane29_strm0_ready      ),      
               .std__pe11__lane29_strm0_cntl          ( std__pe11__lane29_strm0_cntl       ),      
               .std__pe11__lane29_strm0_data          ( std__pe11__lane29_strm0_data       ),      
               .std__pe11__lane29_strm0_data_valid    ( std__pe11__lane29_strm0_data_valid ),      
               .std__pe11__lane29_strm0_data_mask     ( std__pe11__lane29_strm0_data_mask  ),      

               .pe11__std__lane29_strm1_ready         ( pe11__std__lane29_strm1_ready      ),      
               .std__pe11__lane29_strm1_cntl          ( std__pe11__lane29_strm1_cntl       ),      
               .std__pe11__lane29_strm1_data          ( std__pe11__lane29_strm1_data       ),      
               .std__pe11__lane29_strm1_data_valid    ( std__pe11__lane29_strm1_data_valid ),      
               .std__pe11__lane29_strm1_data_mask     ( std__pe11__lane29_strm1_data_mask  ),      

               // PE 11, Lane 30                 
               .pe11__std__lane30_strm0_ready         ( pe11__std__lane30_strm0_ready      ),      
               .std__pe11__lane30_strm0_cntl          ( std__pe11__lane30_strm0_cntl       ),      
               .std__pe11__lane30_strm0_data          ( std__pe11__lane30_strm0_data       ),      
               .std__pe11__lane30_strm0_data_valid    ( std__pe11__lane30_strm0_data_valid ),      
               .std__pe11__lane30_strm0_data_mask     ( std__pe11__lane30_strm0_data_mask  ),      

               .pe11__std__lane30_strm1_ready         ( pe11__std__lane30_strm1_ready      ),      
               .std__pe11__lane30_strm1_cntl          ( std__pe11__lane30_strm1_cntl       ),      
               .std__pe11__lane30_strm1_data          ( std__pe11__lane30_strm1_data       ),      
               .std__pe11__lane30_strm1_data_valid    ( std__pe11__lane30_strm1_data_valid ),      
               .std__pe11__lane30_strm1_data_mask     ( std__pe11__lane30_strm1_data_mask  ),      

               // PE 11, Lane 31                 
               .pe11__std__lane31_strm0_ready         ( pe11__std__lane31_strm0_ready      ),      
               .std__pe11__lane31_strm0_cntl          ( std__pe11__lane31_strm0_cntl       ),      
               .std__pe11__lane31_strm0_data          ( std__pe11__lane31_strm0_data       ),      
               .std__pe11__lane31_strm0_data_valid    ( std__pe11__lane31_strm0_data_valid ),      
               .std__pe11__lane31_strm0_data_mask     ( std__pe11__lane31_strm0_data_mask  ),      

               .pe11__std__lane31_strm1_ready         ( pe11__std__lane31_strm1_ready      ),      
               .std__pe11__lane31_strm1_cntl          ( std__pe11__lane31_strm1_cntl       ),      
               .std__pe11__lane31_strm1_data          ( std__pe11__lane31_strm1_data       ),      
               .std__pe11__lane31_strm1_data_valid    ( std__pe11__lane31_strm1_data_valid ),      
               .std__pe11__lane31_strm1_data_mask     ( std__pe11__lane31_strm1_data_mask  ),      

               // PE 12, Lane 0                 
               .pe12__std__lane0_strm0_ready         ( pe12__std__lane0_strm0_ready      ),      
               .std__pe12__lane0_strm0_cntl          ( std__pe12__lane0_strm0_cntl       ),      
               .std__pe12__lane0_strm0_data          ( std__pe12__lane0_strm0_data       ),      
               .std__pe12__lane0_strm0_data_valid    ( std__pe12__lane0_strm0_data_valid ),      
               .std__pe12__lane0_strm0_data_mask     ( std__pe12__lane0_strm0_data_mask  ),      

               .pe12__std__lane0_strm1_ready         ( pe12__std__lane0_strm1_ready      ),      
               .std__pe12__lane0_strm1_cntl          ( std__pe12__lane0_strm1_cntl       ),      
               .std__pe12__lane0_strm1_data          ( std__pe12__lane0_strm1_data       ),      
               .std__pe12__lane0_strm1_data_valid    ( std__pe12__lane0_strm1_data_valid ),      
               .std__pe12__lane0_strm1_data_mask     ( std__pe12__lane0_strm1_data_mask  ),      

               // PE 12, Lane 1                 
               .pe12__std__lane1_strm0_ready         ( pe12__std__lane1_strm0_ready      ),      
               .std__pe12__lane1_strm0_cntl          ( std__pe12__lane1_strm0_cntl       ),      
               .std__pe12__lane1_strm0_data          ( std__pe12__lane1_strm0_data       ),      
               .std__pe12__lane1_strm0_data_valid    ( std__pe12__lane1_strm0_data_valid ),      
               .std__pe12__lane1_strm0_data_mask     ( std__pe12__lane1_strm0_data_mask  ),      

               .pe12__std__lane1_strm1_ready         ( pe12__std__lane1_strm1_ready      ),      
               .std__pe12__lane1_strm1_cntl          ( std__pe12__lane1_strm1_cntl       ),      
               .std__pe12__lane1_strm1_data          ( std__pe12__lane1_strm1_data       ),      
               .std__pe12__lane1_strm1_data_valid    ( std__pe12__lane1_strm1_data_valid ),      
               .std__pe12__lane1_strm1_data_mask     ( std__pe12__lane1_strm1_data_mask  ),      

               // PE 12, Lane 2                 
               .pe12__std__lane2_strm0_ready         ( pe12__std__lane2_strm0_ready      ),      
               .std__pe12__lane2_strm0_cntl          ( std__pe12__lane2_strm0_cntl       ),      
               .std__pe12__lane2_strm0_data          ( std__pe12__lane2_strm0_data       ),      
               .std__pe12__lane2_strm0_data_valid    ( std__pe12__lane2_strm0_data_valid ),      
               .std__pe12__lane2_strm0_data_mask     ( std__pe12__lane2_strm0_data_mask  ),      

               .pe12__std__lane2_strm1_ready         ( pe12__std__lane2_strm1_ready      ),      
               .std__pe12__lane2_strm1_cntl          ( std__pe12__lane2_strm1_cntl       ),      
               .std__pe12__lane2_strm1_data          ( std__pe12__lane2_strm1_data       ),      
               .std__pe12__lane2_strm1_data_valid    ( std__pe12__lane2_strm1_data_valid ),      
               .std__pe12__lane2_strm1_data_mask     ( std__pe12__lane2_strm1_data_mask  ),      

               // PE 12, Lane 3                 
               .pe12__std__lane3_strm0_ready         ( pe12__std__lane3_strm0_ready      ),      
               .std__pe12__lane3_strm0_cntl          ( std__pe12__lane3_strm0_cntl       ),      
               .std__pe12__lane3_strm0_data          ( std__pe12__lane3_strm0_data       ),      
               .std__pe12__lane3_strm0_data_valid    ( std__pe12__lane3_strm0_data_valid ),      
               .std__pe12__lane3_strm0_data_mask     ( std__pe12__lane3_strm0_data_mask  ),      

               .pe12__std__lane3_strm1_ready         ( pe12__std__lane3_strm1_ready      ),      
               .std__pe12__lane3_strm1_cntl          ( std__pe12__lane3_strm1_cntl       ),      
               .std__pe12__lane3_strm1_data          ( std__pe12__lane3_strm1_data       ),      
               .std__pe12__lane3_strm1_data_valid    ( std__pe12__lane3_strm1_data_valid ),      
               .std__pe12__lane3_strm1_data_mask     ( std__pe12__lane3_strm1_data_mask  ),      

               // PE 12, Lane 4                 
               .pe12__std__lane4_strm0_ready         ( pe12__std__lane4_strm0_ready      ),      
               .std__pe12__lane4_strm0_cntl          ( std__pe12__lane4_strm0_cntl       ),      
               .std__pe12__lane4_strm0_data          ( std__pe12__lane4_strm0_data       ),      
               .std__pe12__lane4_strm0_data_valid    ( std__pe12__lane4_strm0_data_valid ),      
               .std__pe12__lane4_strm0_data_mask     ( std__pe12__lane4_strm0_data_mask  ),      

               .pe12__std__lane4_strm1_ready         ( pe12__std__lane4_strm1_ready      ),      
               .std__pe12__lane4_strm1_cntl          ( std__pe12__lane4_strm1_cntl       ),      
               .std__pe12__lane4_strm1_data          ( std__pe12__lane4_strm1_data       ),      
               .std__pe12__lane4_strm1_data_valid    ( std__pe12__lane4_strm1_data_valid ),      
               .std__pe12__lane4_strm1_data_mask     ( std__pe12__lane4_strm1_data_mask  ),      

               // PE 12, Lane 5                 
               .pe12__std__lane5_strm0_ready         ( pe12__std__lane5_strm0_ready      ),      
               .std__pe12__lane5_strm0_cntl          ( std__pe12__lane5_strm0_cntl       ),      
               .std__pe12__lane5_strm0_data          ( std__pe12__lane5_strm0_data       ),      
               .std__pe12__lane5_strm0_data_valid    ( std__pe12__lane5_strm0_data_valid ),      
               .std__pe12__lane5_strm0_data_mask     ( std__pe12__lane5_strm0_data_mask  ),      

               .pe12__std__lane5_strm1_ready         ( pe12__std__lane5_strm1_ready      ),      
               .std__pe12__lane5_strm1_cntl          ( std__pe12__lane5_strm1_cntl       ),      
               .std__pe12__lane5_strm1_data          ( std__pe12__lane5_strm1_data       ),      
               .std__pe12__lane5_strm1_data_valid    ( std__pe12__lane5_strm1_data_valid ),      
               .std__pe12__lane5_strm1_data_mask     ( std__pe12__lane5_strm1_data_mask  ),      

               // PE 12, Lane 6                 
               .pe12__std__lane6_strm0_ready         ( pe12__std__lane6_strm0_ready      ),      
               .std__pe12__lane6_strm0_cntl          ( std__pe12__lane6_strm0_cntl       ),      
               .std__pe12__lane6_strm0_data          ( std__pe12__lane6_strm0_data       ),      
               .std__pe12__lane6_strm0_data_valid    ( std__pe12__lane6_strm0_data_valid ),      
               .std__pe12__lane6_strm0_data_mask     ( std__pe12__lane6_strm0_data_mask  ),      

               .pe12__std__lane6_strm1_ready         ( pe12__std__lane6_strm1_ready      ),      
               .std__pe12__lane6_strm1_cntl          ( std__pe12__lane6_strm1_cntl       ),      
               .std__pe12__lane6_strm1_data          ( std__pe12__lane6_strm1_data       ),      
               .std__pe12__lane6_strm1_data_valid    ( std__pe12__lane6_strm1_data_valid ),      
               .std__pe12__lane6_strm1_data_mask     ( std__pe12__lane6_strm1_data_mask  ),      

               // PE 12, Lane 7                 
               .pe12__std__lane7_strm0_ready         ( pe12__std__lane7_strm0_ready      ),      
               .std__pe12__lane7_strm0_cntl          ( std__pe12__lane7_strm0_cntl       ),      
               .std__pe12__lane7_strm0_data          ( std__pe12__lane7_strm0_data       ),      
               .std__pe12__lane7_strm0_data_valid    ( std__pe12__lane7_strm0_data_valid ),      
               .std__pe12__lane7_strm0_data_mask     ( std__pe12__lane7_strm0_data_mask  ),      

               .pe12__std__lane7_strm1_ready         ( pe12__std__lane7_strm1_ready      ),      
               .std__pe12__lane7_strm1_cntl          ( std__pe12__lane7_strm1_cntl       ),      
               .std__pe12__lane7_strm1_data          ( std__pe12__lane7_strm1_data       ),      
               .std__pe12__lane7_strm1_data_valid    ( std__pe12__lane7_strm1_data_valid ),      
               .std__pe12__lane7_strm1_data_mask     ( std__pe12__lane7_strm1_data_mask  ),      

               // PE 12, Lane 8                 
               .pe12__std__lane8_strm0_ready         ( pe12__std__lane8_strm0_ready      ),      
               .std__pe12__lane8_strm0_cntl          ( std__pe12__lane8_strm0_cntl       ),      
               .std__pe12__lane8_strm0_data          ( std__pe12__lane8_strm0_data       ),      
               .std__pe12__lane8_strm0_data_valid    ( std__pe12__lane8_strm0_data_valid ),      
               .std__pe12__lane8_strm0_data_mask     ( std__pe12__lane8_strm0_data_mask  ),      

               .pe12__std__lane8_strm1_ready         ( pe12__std__lane8_strm1_ready      ),      
               .std__pe12__lane8_strm1_cntl          ( std__pe12__lane8_strm1_cntl       ),      
               .std__pe12__lane8_strm1_data          ( std__pe12__lane8_strm1_data       ),      
               .std__pe12__lane8_strm1_data_valid    ( std__pe12__lane8_strm1_data_valid ),      
               .std__pe12__lane8_strm1_data_mask     ( std__pe12__lane8_strm1_data_mask  ),      

               // PE 12, Lane 9                 
               .pe12__std__lane9_strm0_ready         ( pe12__std__lane9_strm0_ready      ),      
               .std__pe12__lane9_strm0_cntl          ( std__pe12__lane9_strm0_cntl       ),      
               .std__pe12__lane9_strm0_data          ( std__pe12__lane9_strm0_data       ),      
               .std__pe12__lane9_strm0_data_valid    ( std__pe12__lane9_strm0_data_valid ),      
               .std__pe12__lane9_strm0_data_mask     ( std__pe12__lane9_strm0_data_mask  ),      

               .pe12__std__lane9_strm1_ready         ( pe12__std__lane9_strm1_ready      ),      
               .std__pe12__lane9_strm1_cntl          ( std__pe12__lane9_strm1_cntl       ),      
               .std__pe12__lane9_strm1_data          ( std__pe12__lane9_strm1_data       ),      
               .std__pe12__lane9_strm1_data_valid    ( std__pe12__lane9_strm1_data_valid ),      
               .std__pe12__lane9_strm1_data_mask     ( std__pe12__lane9_strm1_data_mask  ),      

               // PE 12, Lane 10                 
               .pe12__std__lane10_strm0_ready         ( pe12__std__lane10_strm0_ready      ),      
               .std__pe12__lane10_strm0_cntl          ( std__pe12__lane10_strm0_cntl       ),      
               .std__pe12__lane10_strm0_data          ( std__pe12__lane10_strm0_data       ),      
               .std__pe12__lane10_strm0_data_valid    ( std__pe12__lane10_strm0_data_valid ),      
               .std__pe12__lane10_strm0_data_mask     ( std__pe12__lane10_strm0_data_mask  ),      

               .pe12__std__lane10_strm1_ready         ( pe12__std__lane10_strm1_ready      ),      
               .std__pe12__lane10_strm1_cntl          ( std__pe12__lane10_strm1_cntl       ),      
               .std__pe12__lane10_strm1_data          ( std__pe12__lane10_strm1_data       ),      
               .std__pe12__lane10_strm1_data_valid    ( std__pe12__lane10_strm1_data_valid ),      
               .std__pe12__lane10_strm1_data_mask     ( std__pe12__lane10_strm1_data_mask  ),      

               // PE 12, Lane 11                 
               .pe12__std__lane11_strm0_ready         ( pe12__std__lane11_strm0_ready      ),      
               .std__pe12__lane11_strm0_cntl          ( std__pe12__lane11_strm0_cntl       ),      
               .std__pe12__lane11_strm0_data          ( std__pe12__lane11_strm0_data       ),      
               .std__pe12__lane11_strm0_data_valid    ( std__pe12__lane11_strm0_data_valid ),      
               .std__pe12__lane11_strm0_data_mask     ( std__pe12__lane11_strm0_data_mask  ),      

               .pe12__std__lane11_strm1_ready         ( pe12__std__lane11_strm1_ready      ),      
               .std__pe12__lane11_strm1_cntl          ( std__pe12__lane11_strm1_cntl       ),      
               .std__pe12__lane11_strm1_data          ( std__pe12__lane11_strm1_data       ),      
               .std__pe12__lane11_strm1_data_valid    ( std__pe12__lane11_strm1_data_valid ),      
               .std__pe12__lane11_strm1_data_mask     ( std__pe12__lane11_strm1_data_mask  ),      

               // PE 12, Lane 12                 
               .pe12__std__lane12_strm0_ready         ( pe12__std__lane12_strm0_ready      ),      
               .std__pe12__lane12_strm0_cntl          ( std__pe12__lane12_strm0_cntl       ),      
               .std__pe12__lane12_strm0_data          ( std__pe12__lane12_strm0_data       ),      
               .std__pe12__lane12_strm0_data_valid    ( std__pe12__lane12_strm0_data_valid ),      
               .std__pe12__lane12_strm0_data_mask     ( std__pe12__lane12_strm0_data_mask  ),      

               .pe12__std__lane12_strm1_ready         ( pe12__std__lane12_strm1_ready      ),      
               .std__pe12__lane12_strm1_cntl          ( std__pe12__lane12_strm1_cntl       ),      
               .std__pe12__lane12_strm1_data          ( std__pe12__lane12_strm1_data       ),      
               .std__pe12__lane12_strm1_data_valid    ( std__pe12__lane12_strm1_data_valid ),      
               .std__pe12__lane12_strm1_data_mask     ( std__pe12__lane12_strm1_data_mask  ),      

               // PE 12, Lane 13                 
               .pe12__std__lane13_strm0_ready         ( pe12__std__lane13_strm0_ready      ),      
               .std__pe12__lane13_strm0_cntl          ( std__pe12__lane13_strm0_cntl       ),      
               .std__pe12__lane13_strm0_data          ( std__pe12__lane13_strm0_data       ),      
               .std__pe12__lane13_strm0_data_valid    ( std__pe12__lane13_strm0_data_valid ),      
               .std__pe12__lane13_strm0_data_mask     ( std__pe12__lane13_strm0_data_mask  ),      

               .pe12__std__lane13_strm1_ready         ( pe12__std__lane13_strm1_ready      ),      
               .std__pe12__lane13_strm1_cntl          ( std__pe12__lane13_strm1_cntl       ),      
               .std__pe12__lane13_strm1_data          ( std__pe12__lane13_strm1_data       ),      
               .std__pe12__lane13_strm1_data_valid    ( std__pe12__lane13_strm1_data_valid ),      
               .std__pe12__lane13_strm1_data_mask     ( std__pe12__lane13_strm1_data_mask  ),      

               // PE 12, Lane 14                 
               .pe12__std__lane14_strm0_ready         ( pe12__std__lane14_strm0_ready      ),      
               .std__pe12__lane14_strm0_cntl          ( std__pe12__lane14_strm0_cntl       ),      
               .std__pe12__lane14_strm0_data          ( std__pe12__lane14_strm0_data       ),      
               .std__pe12__lane14_strm0_data_valid    ( std__pe12__lane14_strm0_data_valid ),      
               .std__pe12__lane14_strm0_data_mask     ( std__pe12__lane14_strm0_data_mask  ),      

               .pe12__std__lane14_strm1_ready         ( pe12__std__lane14_strm1_ready      ),      
               .std__pe12__lane14_strm1_cntl          ( std__pe12__lane14_strm1_cntl       ),      
               .std__pe12__lane14_strm1_data          ( std__pe12__lane14_strm1_data       ),      
               .std__pe12__lane14_strm1_data_valid    ( std__pe12__lane14_strm1_data_valid ),      
               .std__pe12__lane14_strm1_data_mask     ( std__pe12__lane14_strm1_data_mask  ),      

               // PE 12, Lane 15                 
               .pe12__std__lane15_strm0_ready         ( pe12__std__lane15_strm0_ready      ),      
               .std__pe12__lane15_strm0_cntl          ( std__pe12__lane15_strm0_cntl       ),      
               .std__pe12__lane15_strm0_data          ( std__pe12__lane15_strm0_data       ),      
               .std__pe12__lane15_strm0_data_valid    ( std__pe12__lane15_strm0_data_valid ),      
               .std__pe12__lane15_strm0_data_mask     ( std__pe12__lane15_strm0_data_mask  ),      

               .pe12__std__lane15_strm1_ready         ( pe12__std__lane15_strm1_ready      ),      
               .std__pe12__lane15_strm1_cntl          ( std__pe12__lane15_strm1_cntl       ),      
               .std__pe12__lane15_strm1_data          ( std__pe12__lane15_strm1_data       ),      
               .std__pe12__lane15_strm1_data_valid    ( std__pe12__lane15_strm1_data_valid ),      
               .std__pe12__lane15_strm1_data_mask     ( std__pe12__lane15_strm1_data_mask  ),      

               // PE 12, Lane 16                 
               .pe12__std__lane16_strm0_ready         ( pe12__std__lane16_strm0_ready      ),      
               .std__pe12__lane16_strm0_cntl          ( std__pe12__lane16_strm0_cntl       ),      
               .std__pe12__lane16_strm0_data          ( std__pe12__lane16_strm0_data       ),      
               .std__pe12__lane16_strm0_data_valid    ( std__pe12__lane16_strm0_data_valid ),      
               .std__pe12__lane16_strm0_data_mask     ( std__pe12__lane16_strm0_data_mask  ),      

               .pe12__std__lane16_strm1_ready         ( pe12__std__lane16_strm1_ready      ),      
               .std__pe12__lane16_strm1_cntl          ( std__pe12__lane16_strm1_cntl       ),      
               .std__pe12__lane16_strm1_data          ( std__pe12__lane16_strm1_data       ),      
               .std__pe12__lane16_strm1_data_valid    ( std__pe12__lane16_strm1_data_valid ),      
               .std__pe12__lane16_strm1_data_mask     ( std__pe12__lane16_strm1_data_mask  ),      

               // PE 12, Lane 17                 
               .pe12__std__lane17_strm0_ready         ( pe12__std__lane17_strm0_ready      ),      
               .std__pe12__lane17_strm0_cntl          ( std__pe12__lane17_strm0_cntl       ),      
               .std__pe12__lane17_strm0_data          ( std__pe12__lane17_strm0_data       ),      
               .std__pe12__lane17_strm0_data_valid    ( std__pe12__lane17_strm0_data_valid ),      
               .std__pe12__lane17_strm0_data_mask     ( std__pe12__lane17_strm0_data_mask  ),      

               .pe12__std__lane17_strm1_ready         ( pe12__std__lane17_strm1_ready      ),      
               .std__pe12__lane17_strm1_cntl          ( std__pe12__lane17_strm1_cntl       ),      
               .std__pe12__lane17_strm1_data          ( std__pe12__lane17_strm1_data       ),      
               .std__pe12__lane17_strm1_data_valid    ( std__pe12__lane17_strm1_data_valid ),      
               .std__pe12__lane17_strm1_data_mask     ( std__pe12__lane17_strm1_data_mask  ),      

               // PE 12, Lane 18                 
               .pe12__std__lane18_strm0_ready         ( pe12__std__lane18_strm0_ready      ),      
               .std__pe12__lane18_strm0_cntl          ( std__pe12__lane18_strm0_cntl       ),      
               .std__pe12__lane18_strm0_data          ( std__pe12__lane18_strm0_data       ),      
               .std__pe12__lane18_strm0_data_valid    ( std__pe12__lane18_strm0_data_valid ),      
               .std__pe12__lane18_strm0_data_mask     ( std__pe12__lane18_strm0_data_mask  ),      

               .pe12__std__lane18_strm1_ready         ( pe12__std__lane18_strm1_ready      ),      
               .std__pe12__lane18_strm1_cntl          ( std__pe12__lane18_strm1_cntl       ),      
               .std__pe12__lane18_strm1_data          ( std__pe12__lane18_strm1_data       ),      
               .std__pe12__lane18_strm1_data_valid    ( std__pe12__lane18_strm1_data_valid ),      
               .std__pe12__lane18_strm1_data_mask     ( std__pe12__lane18_strm1_data_mask  ),      

               // PE 12, Lane 19                 
               .pe12__std__lane19_strm0_ready         ( pe12__std__lane19_strm0_ready      ),      
               .std__pe12__lane19_strm0_cntl          ( std__pe12__lane19_strm0_cntl       ),      
               .std__pe12__lane19_strm0_data          ( std__pe12__lane19_strm0_data       ),      
               .std__pe12__lane19_strm0_data_valid    ( std__pe12__lane19_strm0_data_valid ),      
               .std__pe12__lane19_strm0_data_mask     ( std__pe12__lane19_strm0_data_mask  ),      

               .pe12__std__lane19_strm1_ready         ( pe12__std__lane19_strm1_ready      ),      
               .std__pe12__lane19_strm1_cntl          ( std__pe12__lane19_strm1_cntl       ),      
               .std__pe12__lane19_strm1_data          ( std__pe12__lane19_strm1_data       ),      
               .std__pe12__lane19_strm1_data_valid    ( std__pe12__lane19_strm1_data_valid ),      
               .std__pe12__lane19_strm1_data_mask     ( std__pe12__lane19_strm1_data_mask  ),      

               // PE 12, Lane 20                 
               .pe12__std__lane20_strm0_ready         ( pe12__std__lane20_strm0_ready      ),      
               .std__pe12__lane20_strm0_cntl          ( std__pe12__lane20_strm0_cntl       ),      
               .std__pe12__lane20_strm0_data          ( std__pe12__lane20_strm0_data       ),      
               .std__pe12__lane20_strm0_data_valid    ( std__pe12__lane20_strm0_data_valid ),      
               .std__pe12__lane20_strm0_data_mask     ( std__pe12__lane20_strm0_data_mask  ),      

               .pe12__std__lane20_strm1_ready         ( pe12__std__lane20_strm1_ready      ),      
               .std__pe12__lane20_strm1_cntl          ( std__pe12__lane20_strm1_cntl       ),      
               .std__pe12__lane20_strm1_data          ( std__pe12__lane20_strm1_data       ),      
               .std__pe12__lane20_strm1_data_valid    ( std__pe12__lane20_strm1_data_valid ),      
               .std__pe12__lane20_strm1_data_mask     ( std__pe12__lane20_strm1_data_mask  ),      

               // PE 12, Lane 21                 
               .pe12__std__lane21_strm0_ready         ( pe12__std__lane21_strm0_ready      ),      
               .std__pe12__lane21_strm0_cntl          ( std__pe12__lane21_strm0_cntl       ),      
               .std__pe12__lane21_strm0_data          ( std__pe12__lane21_strm0_data       ),      
               .std__pe12__lane21_strm0_data_valid    ( std__pe12__lane21_strm0_data_valid ),      
               .std__pe12__lane21_strm0_data_mask     ( std__pe12__lane21_strm0_data_mask  ),      

               .pe12__std__lane21_strm1_ready         ( pe12__std__lane21_strm1_ready      ),      
               .std__pe12__lane21_strm1_cntl          ( std__pe12__lane21_strm1_cntl       ),      
               .std__pe12__lane21_strm1_data          ( std__pe12__lane21_strm1_data       ),      
               .std__pe12__lane21_strm1_data_valid    ( std__pe12__lane21_strm1_data_valid ),      
               .std__pe12__lane21_strm1_data_mask     ( std__pe12__lane21_strm1_data_mask  ),      

               // PE 12, Lane 22                 
               .pe12__std__lane22_strm0_ready         ( pe12__std__lane22_strm0_ready      ),      
               .std__pe12__lane22_strm0_cntl          ( std__pe12__lane22_strm0_cntl       ),      
               .std__pe12__lane22_strm0_data          ( std__pe12__lane22_strm0_data       ),      
               .std__pe12__lane22_strm0_data_valid    ( std__pe12__lane22_strm0_data_valid ),      
               .std__pe12__lane22_strm0_data_mask     ( std__pe12__lane22_strm0_data_mask  ),      

               .pe12__std__lane22_strm1_ready         ( pe12__std__lane22_strm1_ready      ),      
               .std__pe12__lane22_strm1_cntl          ( std__pe12__lane22_strm1_cntl       ),      
               .std__pe12__lane22_strm1_data          ( std__pe12__lane22_strm1_data       ),      
               .std__pe12__lane22_strm1_data_valid    ( std__pe12__lane22_strm1_data_valid ),      
               .std__pe12__lane22_strm1_data_mask     ( std__pe12__lane22_strm1_data_mask  ),      

               // PE 12, Lane 23                 
               .pe12__std__lane23_strm0_ready         ( pe12__std__lane23_strm0_ready      ),      
               .std__pe12__lane23_strm0_cntl          ( std__pe12__lane23_strm0_cntl       ),      
               .std__pe12__lane23_strm0_data          ( std__pe12__lane23_strm0_data       ),      
               .std__pe12__lane23_strm0_data_valid    ( std__pe12__lane23_strm0_data_valid ),      
               .std__pe12__lane23_strm0_data_mask     ( std__pe12__lane23_strm0_data_mask  ),      

               .pe12__std__lane23_strm1_ready         ( pe12__std__lane23_strm1_ready      ),      
               .std__pe12__lane23_strm1_cntl          ( std__pe12__lane23_strm1_cntl       ),      
               .std__pe12__lane23_strm1_data          ( std__pe12__lane23_strm1_data       ),      
               .std__pe12__lane23_strm1_data_valid    ( std__pe12__lane23_strm1_data_valid ),      
               .std__pe12__lane23_strm1_data_mask     ( std__pe12__lane23_strm1_data_mask  ),      

               // PE 12, Lane 24                 
               .pe12__std__lane24_strm0_ready         ( pe12__std__lane24_strm0_ready      ),      
               .std__pe12__lane24_strm0_cntl          ( std__pe12__lane24_strm0_cntl       ),      
               .std__pe12__lane24_strm0_data          ( std__pe12__lane24_strm0_data       ),      
               .std__pe12__lane24_strm0_data_valid    ( std__pe12__lane24_strm0_data_valid ),      
               .std__pe12__lane24_strm0_data_mask     ( std__pe12__lane24_strm0_data_mask  ),      

               .pe12__std__lane24_strm1_ready         ( pe12__std__lane24_strm1_ready      ),      
               .std__pe12__lane24_strm1_cntl          ( std__pe12__lane24_strm1_cntl       ),      
               .std__pe12__lane24_strm1_data          ( std__pe12__lane24_strm1_data       ),      
               .std__pe12__lane24_strm1_data_valid    ( std__pe12__lane24_strm1_data_valid ),      
               .std__pe12__lane24_strm1_data_mask     ( std__pe12__lane24_strm1_data_mask  ),      

               // PE 12, Lane 25                 
               .pe12__std__lane25_strm0_ready         ( pe12__std__lane25_strm0_ready      ),      
               .std__pe12__lane25_strm0_cntl          ( std__pe12__lane25_strm0_cntl       ),      
               .std__pe12__lane25_strm0_data          ( std__pe12__lane25_strm0_data       ),      
               .std__pe12__lane25_strm0_data_valid    ( std__pe12__lane25_strm0_data_valid ),      
               .std__pe12__lane25_strm0_data_mask     ( std__pe12__lane25_strm0_data_mask  ),      

               .pe12__std__lane25_strm1_ready         ( pe12__std__lane25_strm1_ready      ),      
               .std__pe12__lane25_strm1_cntl          ( std__pe12__lane25_strm1_cntl       ),      
               .std__pe12__lane25_strm1_data          ( std__pe12__lane25_strm1_data       ),      
               .std__pe12__lane25_strm1_data_valid    ( std__pe12__lane25_strm1_data_valid ),      
               .std__pe12__lane25_strm1_data_mask     ( std__pe12__lane25_strm1_data_mask  ),      

               // PE 12, Lane 26                 
               .pe12__std__lane26_strm0_ready         ( pe12__std__lane26_strm0_ready      ),      
               .std__pe12__lane26_strm0_cntl          ( std__pe12__lane26_strm0_cntl       ),      
               .std__pe12__lane26_strm0_data          ( std__pe12__lane26_strm0_data       ),      
               .std__pe12__lane26_strm0_data_valid    ( std__pe12__lane26_strm0_data_valid ),      
               .std__pe12__lane26_strm0_data_mask     ( std__pe12__lane26_strm0_data_mask  ),      

               .pe12__std__lane26_strm1_ready         ( pe12__std__lane26_strm1_ready      ),      
               .std__pe12__lane26_strm1_cntl          ( std__pe12__lane26_strm1_cntl       ),      
               .std__pe12__lane26_strm1_data          ( std__pe12__lane26_strm1_data       ),      
               .std__pe12__lane26_strm1_data_valid    ( std__pe12__lane26_strm1_data_valid ),      
               .std__pe12__lane26_strm1_data_mask     ( std__pe12__lane26_strm1_data_mask  ),      

               // PE 12, Lane 27                 
               .pe12__std__lane27_strm0_ready         ( pe12__std__lane27_strm0_ready      ),      
               .std__pe12__lane27_strm0_cntl          ( std__pe12__lane27_strm0_cntl       ),      
               .std__pe12__lane27_strm0_data          ( std__pe12__lane27_strm0_data       ),      
               .std__pe12__lane27_strm0_data_valid    ( std__pe12__lane27_strm0_data_valid ),      
               .std__pe12__lane27_strm0_data_mask     ( std__pe12__lane27_strm0_data_mask  ),      

               .pe12__std__lane27_strm1_ready         ( pe12__std__lane27_strm1_ready      ),      
               .std__pe12__lane27_strm1_cntl          ( std__pe12__lane27_strm1_cntl       ),      
               .std__pe12__lane27_strm1_data          ( std__pe12__lane27_strm1_data       ),      
               .std__pe12__lane27_strm1_data_valid    ( std__pe12__lane27_strm1_data_valid ),      
               .std__pe12__lane27_strm1_data_mask     ( std__pe12__lane27_strm1_data_mask  ),      

               // PE 12, Lane 28                 
               .pe12__std__lane28_strm0_ready         ( pe12__std__lane28_strm0_ready      ),      
               .std__pe12__lane28_strm0_cntl          ( std__pe12__lane28_strm0_cntl       ),      
               .std__pe12__lane28_strm0_data          ( std__pe12__lane28_strm0_data       ),      
               .std__pe12__lane28_strm0_data_valid    ( std__pe12__lane28_strm0_data_valid ),      
               .std__pe12__lane28_strm0_data_mask     ( std__pe12__lane28_strm0_data_mask  ),      

               .pe12__std__lane28_strm1_ready         ( pe12__std__lane28_strm1_ready      ),      
               .std__pe12__lane28_strm1_cntl          ( std__pe12__lane28_strm1_cntl       ),      
               .std__pe12__lane28_strm1_data          ( std__pe12__lane28_strm1_data       ),      
               .std__pe12__lane28_strm1_data_valid    ( std__pe12__lane28_strm1_data_valid ),      
               .std__pe12__lane28_strm1_data_mask     ( std__pe12__lane28_strm1_data_mask  ),      

               // PE 12, Lane 29                 
               .pe12__std__lane29_strm0_ready         ( pe12__std__lane29_strm0_ready      ),      
               .std__pe12__lane29_strm0_cntl          ( std__pe12__lane29_strm0_cntl       ),      
               .std__pe12__lane29_strm0_data          ( std__pe12__lane29_strm0_data       ),      
               .std__pe12__lane29_strm0_data_valid    ( std__pe12__lane29_strm0_data_valid ),      
               .std__pe12__lane29_strm0_data_mask     ( std__pe12__lane29_strm0_data_mask  ),      

               .pe12__std__lane29_strm1_ready         ( pe12__std__lane29_strm1_ready      ),      
               .std__pe12__lane29_strm1_cntl          ( std__pe12__lane29_strm1_cntl       ),      
               .std__pe12__lane29_strm1_data          ( std__pe12__lane29_strm1_data       ),      
               .std__pe12__lane29_strm1_data_valid    ( std__pe12__lane29_strm1_data_valid ),      
               .std__pe12__lane29_strm1_data_mask     ( std__pe12__lane29_strm1_data_mask  ),      

               // PE 12, Lane 30                 
               .pe12__std__lane30_strm0_ready         ( pe12__std__lane30_strm0_ready      ),      
               .std__pe12__lane30_strm0_cntl          ( std__pe12__lane30_strm0_cntl       ),      
               .std__pe12__lane30_strm0_data          ( std__pe12__lane30_strm0_data       ),      
               .std__pe12__lane30_strm0_data_valid    ( std__pe12__lane30_strm0_data_valid ),      
               .std__pe12__lane30_strm0_data_mask     ( std__pe12__lane30_strm0_data_mask  ),      

               .pe12__std__lane30_strm1_ready         ( pe12__std__lane30_strm1_ready      ),      
               .std__pe12__lane30_strm1_cntl          ( std__pe12__lane30_strm1_cntl       ),      
               .std__pe12__lane30_strm1_data          ( std__pe12__lane30_strm1_data       ),      
               .std__pe12__lane30_strm1_data_valid    ( std__pe12__lane30_strm1_data_valid ),      
               .std__pe12__lane30_strm1_data_mask     ( std__pe12__lane30_strm1_data_mask  ),      

               // PE 12, Lane 31                 
               .pe12__std__lane31_strm0_ready         ( pe12__std__lane31_strm0_ready      ),      
               .std__pe12__lane31_strm0_cntl          ( std__pe12__lane31_strm0_cntl       ),      
               .std__pe12__lane31_strm0_data          ( std__pe12__lane31_strm0_data       ),      
               .std__pe12__lane31_strm0_data_valid    ( std__pe12__lane31_strm0_data_valid ),      
               .std__pe12__lane31_strm0_data_mask     ( std__pe12__lane31_strm0_data_mask  ),      

               .pe12__std__lane31_strm1_ready         ( pe12__std__lane31_strm1_ready      ),      
               .std__pe12__lane31_strm1_cntl          ( std__pe12__lane31_strm1_cntl       ),      
               .std__pe12__lane31_strm1_data          ( std__pe12__lane31_strm1_data       ),      
               .std__pe12__lane31_strm1_data_valid    ( std__pe12__lane31_strm1_data_valid ),      
               .std__pe12__lane31_strm1_data_mask     ( std__pe12__lane31_strm1_data_mask  ),      

               // PE 13, Lane 0                 
               .pe13__std__lane0_strm0_ready         ( pe13__std__lane0_strm0_ready      ),      
               .std__pe13__lane0_strm0_cntl          ( std__pe13__lane0_strm0_cntl       ),      
               .std__pe13__lane0_strm0_data          ( std__pe13__lane0_strm0_data       ),      
               .std__pe13__lane0_strm0_data_valid    ( std__pe13__lane0_strm0_data_valid ),      
               .std__pe13__lane0_strm0_data_mask     ( std__pe13__lane0_strm0_data_mask  ),      

               .pe13__std__lane0_strm1_ready         ( pe13__std__lane0_strm1_ready      ),      
               .std__pe13__lane0_strm1_cntl          ( std__pe13__lane0_strm1_cntl       ),      
               .std__pe13__lane0_strm1_data          ( std__pe13__lane0_strm1_data       ),      
               .std__pe13__lane0_strm1_data_valid    ( std__pe13__lane0_strm1_data_valid ),      
               .std__pe13__lane0_strm1_data_mask     ( std__pe13__lane0_strm1_data_mask  ),      

               // PE 13, Lane 1                 
               .pe13__std__lane1_strm0_ready         ( pe13__std__lane1_strm0_ready      ),      
               .std__pe13__lane1_strm0_cntl          ( std__pe13__lane1_strm0_cntl       ),      
               .std__pe13__lane1_strm0_data          ( std__pe13__lane1_strm0_data       ),      
               .std__pe13__lane1_strm0_data_valid    ( std__pe13__lane1_strm0_data_valid ),      
               .std__pe13__lane1_strm0_data_mask     ( std__pe13__lane1_strm0_data_mask  ),      

               .pe13__std__lane1_strm1_ready         ( pe13__std__lane1_strm1_ready      ),      
               .std__pe13__lane1_strm1_cntl          ( std__pe13__lane1_strm1_cntl       ),      
               .std__pe13__lane1_strm1_data          ( std__pe13__lane1_strm1_data       ),      
               .std__pe13__lane1_strm1_data_valid    ( std__pe13__lane1_strm1_data_valid ),      
               .std__pe13__lane1_strm1_data_mask     ( std__pe13__lane1_strm1_data_mask  ),      

               // PE 13, Lane 2                 
               .pe13__std__lane2_strm0_ready         ( pe13__std__lane2_strm0_ready      ),      
               .std__pe13__lane2_strm0_cntl          ( std__pe13__lane2_strm0_cntl       ),      
               .std__pe13__lane2_strm0_data          ( std__pe13__lane2_strm0_data       ),      
               .std__pe13__lane2_strm0_data_valid    ( std__pe13__lane2_strm0_data_valid ),      
               .std__pe13__lane2_strm0_data_mask     ( std__pe13__lane2_strm0_data_mask  ),      

               .pe13__std__lane2_strm1_ready         ( pe13__std__lane2_strm1_ready      ),      
               .std__pe13__lane2_strm1_cntl          ( std__pe13__lane2_strm1_cntl       ),      
               .std__pe13__lane2_strm1_data          ( std__pe13__lane2_strm1_data       ),      
               .std__pe13__lane2_strm1_data_valid    ( std__pe13__lane2_strm1_data_valid ),      
               .std__pe13__lane2_strm1_data_mask     ( std__pe13__lane2_strm1_data_mask  ),      

               // PE 13, Lane 3                 
               .pe13__std__lane3_strm0_ready         ( pe13__std__lane3_strm0_ready      ),      
               .std__pe13__lane3_strm0_cntl          ( std__pe13__lane3_strm0_cntl       ),      
               .std__pe13__lane3_strm0_data          ( std__pe13__lane3_strm0_data       ),      
               .std__pe13__lane3_strm0_data_valid    ( std__pe13__lane3_strm0_data_valid ),      
               .std__pe13__lane3_strm0_data_mask     ( std__pe13__lane3_strm0_data_mask  ),      

               .pe13__std__lane3_strm1_ready         ( pe13__std__lane3_strm1_ready      ),      
               .std__pe13__lane3_strm1_cntl          ( std__pe13__lane3_strm1_cntl       ),      
               .std__pe13__lane3_strm1_data          ( std__pe13__lane3_strm1_data       ),      
               .std__pe13__lane3_strm1_data_valid    ( std__pe13__lane3_strm1_data_valid ),      
               .std__pe13__lane3_strm1_data_mask     ( std__pe13__lane3_strm1_data_mask  ),      

               // PE 13, Lane 4                 
               .pe13__std__lane4_strm0_ready         ( pe13__std__lane4_strm0_ready      ),      
               .std__pe13__lane4_strm0_cntl          ( std__pe13__lane4_strm0_cntl       ),      
               .std__pe13__lane4_strm0_data          ( std__pe13__lane4_strm0_data       ),      
               .std__pe13__lane4_strm0_data_valid    ( std__pe13__lane4_strm0_data_valid ),      
               .std__pe13__lane4_strm0_data_mask     ( std__pe13__lane4_strm0_data_mask  ),      

               .pe13__std__lane4_strm1_ready         ( pe13__std__lane4_strm1_ready      ),      
               .std__pe13__lane4_strm1_cntl          ( std__pe13__lane4_strm1_cntl       ),      
               .std__pe13__lane4_strm1_data          ( std__pe13__lane4_strm1_data       ),      
               .std__pe13__lane4_strm1_data_valid    ( std__pe13__lane4_strm1_data_valid ),      
               .std__pe13__lane4_strm1_data_mask     ( std__pe13__lane4_strm1_data_mask  ),      

               // PE 13, Lane 5                 
               .pe13__std__lane5_strm0_ready         ( pe13__std__lane5_strm0_ready      ),      
               .std__pe13__lane5_strm0_cntl          ( std__pe13__lane5_strm0_cntl       ),      
               .std__pe13__lane5_strm0_data          ( std__pe13__lane5_strm0_data       ),      
               .std__pe13__lane5_strm0_data_valid    ( std__pe13__lane5_strm0_data_valid ),      
               .std__pe13__lane5_strm0_data_mask     ( std__pe13__lane5_strm0_data_mask  ),      

               .pe13__std__lane5_strm1_ready         ( pe13__std__lane5_strm1_ready      ),      
               .std__pe13__lane5_strm1_cntl          ( std__pe13__lane5_strm1_cntl       ),      
               .std__pe13__lane5_strm1_data          ( std__pe13__lane5_strm1_data       ),      
               .std__pe13__lane5_strm1_data_valid    ( std__pe13__lane5_strm1_data_valid ),      
               .std__pe13__lane5_strm1_data_mask     ( std__pe13__lane5_strm1_data_mask  ),      

               // PE 13, Lane 6                 
               .pe13__std__lane6_strm0_ready         ( pe13__std__lane6_strm0_ready      ),      
               .std__pe13__lane6_strm0_cntl          ( std__pe13__lane6_strm0_cntl       ),      
               .std__pe13__lane6_strm0_data          ( std__pe13__lane6_strm0_data       ),      
               .std__pe13__lane6_strm0_data_valid    ( std__pe13__lane6_strm0_data_valid ),      
               .std__pe13__lane6_strm0_data_mask     ( std__pe13__lane6_strm0_data_mask  ),      

               .pe13__std__lane6_strm1_ready         ( pe13__std__lane6_strm1_ready      ),      
               .std__pe13__lane6_strm1_cntl          ( std__pe13__lane6_strm1_cntl       ),      
               .std__pe13__lane6_strm1_data          ( std__pe13__lane6_strm1_data       ),      
               .std__pe13__lane6_strm1_data_valid    ( std__pe13__lane6_strm1_data_valid ),      
               .std__pe13__lane6_strm1_data_mask     ( std__pe13__lane6_strm1_data_mask  ),      

               // PE 13, Lane 7                 
               .pe13__std__lane7_strm0_ready         ( pe13__std__lane7_strm0_ready      ),      
               .std__pe13__lane7_strm0_cntl          ( std__pe13__lane7_strm0_cntl       ),      
               .std__pe13__lane7_strm0_data          ( std__pe13__lane7_strm0_data       ),      
               .std__pe13__lane7_strm0_data_valid    ( std__pe13__lane7_strm0_data_valid ),      
               .std__pe13__lane7_strm0_data_mask     ( std__pe13__lane7_strm0_data_mask  ),      

               .pe13__std__lane7_strm1_ready         ( pe13__std__lane7_strm1_ready      ),      
               .std__pe13__lane7_strm1_cntl          ( std__pe13__lane7_strm1_cntl       ),      
               .std__pe13__lane7_strm1_data          ( std__pe13__lane7_strm1_data       ),      
               .std__pe13__lane7_strm1_data_valid    ( std__pe13__lane7_strm1_data_valid ),      
               .std__pe13__lane7_strm1_data_mask     ( std__pe13__lane7_strm1_data_mask  ),      

               // PE 13, Lane 8                 
               .pe13__std__lane8_strm0_ready         ( pe13__std__lane8_strm0_ready      ),      
               .std__pe13__lane8_strm0_cntl          ( std__pe13__lane8_strm0_cntl       ),      
               .std__pe13__lane8_strm0_data          ( std__pe13__lane8_strm0_data       ),      
               .std__pe13__lane8_strm0_data_valid    ( std__pe13__lane8_strm0_data_valid ),      
               .std__pe13__lane8_strm0_data_mask     ( std__pe13__lane8_strm0_data_mask  ),      

               .pe13__std__lane8_strm1_ready         ( pe13__std__lane8_strm1_ready      ),      
               .std__pe13__lane8_strm1_cntl          ( std__pe13__lane8_strm1_cntl       ),      
               .std__pe13__lane8_strm1_data          ( std__pe13__lane8_strm1_data       ),      
               .std__pe13__lane8_strm1_data_valid    ( std__pe13__lane8_strm1_data_valid ),      
               .std__pe13__lane8_strm1_data_mask     ( std__pe13__lane8_strm1_data_mask  ),      

               // PE 13, Lane 9                 
               .pe13__std__lane9_strm0_ready         ( pe13__std__lane9_strm0_ready      ),      
               .std__pe13__lane9_strm0_cntl          ( std__pe13__lane9_strm0_cntl       ),      
               .std__pe13__lane9_strm0_data          ( std__pe13__lane9_strm0_data       ),      
               .std__pe13__lane9_strm0_data_valid    ( std__pe13__lane9_strm0_data_valid ),      
               .std__pe13__lane9_strm0_data_mask     ( std__pe13__lane9_strm0_data_mask  ),      

               .pe13__std__lane9_strm1_ready         ( pe13__std__lane9_strm1_ready      ),      
               .std__pe13__lane9_strm1_cntl          ( std__pe13__lane9_strm1_cntl       ),      
               .std__pe13__lane9_strm1_data          ( std__pe13__lane9_strm1_data       ),      
               .std__pe13__lane9_strm1_data_valid    ( std__pe13__lane9_strm1_data_valid ),      
               .std__pe13__lane9_strm1_data_mask     ( std__pe13__lane9_strm1_data_mask  ),      

               // PE 13, Lane 10                 
               .pe13__std__lane10_strm0_ready         ( pe13__std__lane10_strm0_ready      ),      
               .std__pe13__lane10_strm0_cntl          ( std__pe13__lane10_strm0_cntl       ),      
               .std__pe13__lane10_strm0_data          ( std__pe13__lane10_strm0_data       ),      
               .std__pe13__lane10_strm0_data_valid    ( std__pe13__lane10_strm0_data_valid ),      
               .std__pe13__lane10_strm0_data_mask     ( std__pe13__lane10_strm0_data_mask  ),      

               .pe13__std__lane10_strm1_ready         ( pe13__std__lane10_strm1_ready      ),      
               .std__pe13__lane10_strm1_cntl          ( std__pe13__lane10_strm1_cntl       ),      
               .std__pe13__lane10_strm1_data          ( std__pe13__lane10_strm1_data       ),      
               .std__pe13__lane10_strm1_data_valid    ( std__pe13__lane10_strm1_data_valid ),      
               .std__pe13__lane10_strm1_data_mask     ( std__pe13__lane10_strm1_data_mask  ),      

               // PE 13, Lane 11                 
               .pe13__std__lane11_strm0_ready         ( pe13__std__lane11_strm0_ready      ),      
               .std__pe13__lane11_strm0_cntl          ( std__pe13__lane11_strm0_cntl       ),      
               .std__pe13__lane11_strm0_data          ( std__pe13__lane11_strm0_data       ),      
               .std__pe13__lane11_strm0_data_valid    ( std__pe13__lane11_strm0_data_valid ),      
               .std__pe13__lane11_strm0_data_mask     ( std__pe13__lane11_strm0_data_mask  ),      

               .pe13__std__lane11_strm1_ready         ( pe13__std__lane11_strm1_ready      ),      
               .std__pe13__lane11_strm1_cntl          ( std__pe13__lane11_strm1_cntl       ),      
               .std__pe13__lane11_strm1_data          ( std__pe13__lane11_strm1_data       ),      
               .std__pe13__lane11_strm1_data_valid    ( std__pe13__lane11_strm1_data_valid ),      
               .std__pe13__lane11_strm1_data_mask     ( std__pe13__lane11_strm1_data_mask  ),      

               // PE 13, Lane 12                 
               .pe13__std__lane12_strm0_ready         ( pe13__std__lane12_strm0_ready      ),      
               .std__pe13__lane12_strm0_cntl          ( std__pe13__lane12_strm0_cntl       ),      
               .std__pe13__lane12_strm0_data          ( std__pe13__lane12_strm0_data       ),      
               .std__pe13__lane12_strm0_data_valid    ( std__pe13__lane12_strm0_data_valid ),      
               .std__pe13__lane12_strm0_data_mask     ( std__pe13__lane12_strm0_data_mask  ),      

               .pe13__std__lane12_strm1_ready         ( pe13__std__lane12_strm1_ready      ),      
               .std__pe13__lane12_strm1_cntl          ( std__pe13__lane12_strm1_cntl       ),      
               .std__pe13__lane12_strm1_data          ( std__pe13__lane12_strm1_data       ),      
               .std__pe13__lane12_strm1_data_valid    ( std__pe13__lane12_strm1_data_valid ),      
               .std__pe13__lane12_strm1_data_mask     ( std__pe13__lane12_strm1_data_mask  ),      

               // PE 13, Lane 13                 
               .pe13__std__lane13_strm0_ready         ( pe13__std__lane13_strm0_ready      ),      
               .std__pe13__lane13_strm0_cntl          ( std__pe13__lane13_strm0_cntl       ),      
               .std__pe13__lane13_strm0_data          ( std__pe13__lane13_strm0_data       ),      
               .std__pe13__lane13_strm0_data_valid    ( std__pe13__lane13_strm0_data_valid ),      
               .std__pe13__lane13_strm0_data_mask     ( std__pe13__lane13_strm0_data_mask  ),      

               .pe13__std__lane13_strm1_ready         ( pe13__std__lane13_strm1_ready      ),      
               .std__pe13__lane13_strm1_cntl          ( std__pe13__lane13_strm1_cntl       ),      
               .std__pe13__lane13_strm1_data          ( std__pe13__lane13_strm1_data       ),      
               .std__pe13__lane13_strm1_data_valid    ( std__pe13__lane13_strm1_data_valid ),      
               .std__pe13__lane13_strm1_data_mask     ( std__pe13__lane13_strm1_data_mask  ),      

               // PE 13, Lane 14                 
               .pe13__std__lane14_strm0_ready         ( pe13__std__lane14_strm0_ready      ),      
               .std__pe13__lane14_strm0_cntl          ( std__pe13__lane14_strm0_cntl       ),      
               .std__pe13__lane14_strm0_data          ( std__pe13__lane14_strm0_data       ),      
               .std__pe13__lane14_strm0_data_valid    ( std__pe13__lane14_strm0_data_valid ),      
               .std__pe13__lane14_strm0_data_mask     ( std__pe13__lane14_strm0_data_mask  ),      

               .pe13__std__lane14_strm1_ready         ( pe13__std__lane14_strm1_ready      ),      
               .std__pe13__lane14_strm1_cntl          ( std__pe13__lane14_strm1_cntl       ),      
               .std__pe13__lane14_strm1_data          ( std__pe13__lane14_strm1_data       ),      
               .std__pe13__lane14_strm1_data_valid    ( std__pe13__lane14_strm1_data_valid ),      
               .std__pe13__lane14_strm1_data_mask     ( std__pe13__lane14_strm1_data_mask  ),      

               // PE 13, Lane 15                 
               .pe13__std__lane15_strm0_ready         ( pe13__std__lane15_strm0_ready      ),      
               .std__pe13__lane15_strm0_cntl          ( std__pe13__lane15_strm0_cntl       ),      
               .std__pe13__lane15_strm0_data          ( std__pe13__lane15_strm0_data       ),      
               .std__pe13__lane15_strm0_data_valid    ( std__pe13__lane15_strm0_data_valid ),      
               .std__pe13__lane15_strm0_data_mask     ( std__pe13__lane15_strm0_data_mask  ),      

               .pe13__std__lane15_strm1_ready         ( pe13__std__lane15_strm1_ready      ),      
               .std__pe13__lane15_strm1_cntl          ( std__pe13__lane15_strm1_cntl       ),      
               .std__pe13__lane15_strm1_data          ( std__pe13__lane15_strm1_data       ),      
               .std__pe13__lane15_strm1_data_valid    ( std__pe13__lane15_strm1_data_valid ),      
               .std__pe13__lane15_strm1_data_mask     ( std__pe13__lane15_strm1_data_mask  ),      

               // PE 13, Lane 16                 
               .pe13__std__lane16_strm0_ready         ( pe13__std__lane16_strm0_ready      ),      
               .std__pe13__lane16_strm0_cntl          ( std__pe13__lane16_strm0_cntl       ),      
               .std__pe13__lane16_strm0_data          ( std__pe13__lane16_strm0_data       ),      
               .std__pe13__lane16_strm0_data_valid    ( std__pe13__lane16_strm0_data_valid ),      
               .std__pe13__lane16_strm0_data_mask     ( std__pe13__lane16_strm0_data_mask  ),      

               .pe13__std__lane16_strm1_ready         ( pe13__std__lane16_strm1_ready      ),      
               .std__pe13__lane16_strm1_cntl          ( std__pe13__lane16_strm1_cntl       ),      
               .std__pe13__lane16_strm1_data          ( std__pe13__lane16_strm1_data       ),      
               .std__pe13__lane16_strm1_data_valid    ( std__pe13__lane16_strm1_data_valid ),      
               .std__pe13__lane16_strm1_data_mask     ( std__pe13__lane16_strm1_data_mask  ),      

               // PE 13, Lane 17                 
               .pe13__std__lane17_strm0_ready         ( pe13__std__lane17_strm0_ready      ),      
               .std__pe13__lane17_strm0_cntl          ( std__pe13__lane17_strm0_cntl       ),      
               .std__pe13__lane17_strm0_data          ( std__pe13__lane17_strm0_data       ),      
               .std__pe13__lane17_strm0_data_valid    ( std__pe13__lane17_strm0_data_valid ),      
               .std__pe13__lane17_strm0_data_mask     ( std__pe13__lane17_strm0_data_mask  ),      

               .pe13__std__lane17_strm1_ready         ( pe13__std__lane17_strm1_ready      ),      
               .std__pe13__lane17_strm1_cntl          ( std__pe13__lane17_strm1_cntl       ),      
               .std__pe13__lane17_strm1_data          ( std__pe13__lane17_strm1_data       ),      
               .std__pe13__lane17_strm1_data_valid    ( std__pe13__lane17_strm1_data_valid ),      
               .std__pe13__lane17_strm1_data_mask     ( std__pe13__lane17_strm1_data_mask  ),      

               // PE 13, Lane 18                 
               .pe13__std__lane18_strm0_ready         ( pe13__std__lane18_strm0_ready      ),      
               .std__pe13__lane18_strm0_cntl          ( std__pe13__lane18_strm0_cntl       ),      
               .std__pe13__lane18_strm0_data          ( std__pe13__lane18_strm0_data       ),      
               .std__pe13__lane18_strm0_data_valid    ( std__pe13__lane18_strm0_data_valid ),      
               .std__pe13__lane18_strm0_data_mask     ( std__pe13__lane18_strm0_data_mask  ),      

               .pe13__std__lane18_strm1_ready         ( pe13__std__lane18_strm1_ready      ),      
               .std__pe13__lane18_strm1_cntl          ( std__pe13__lane18_strm1_cntl       ),      
               .std__pe13__lane18_strm1_data          ( std__pe13__lane18_strm1_data       ),      
               .std__pe13__lane18_strm1_data_valid    ( std__pe13__lane18_strm1_data_valid ),      
               .std__pe13__lane18_strm1_data_mask     ( std__pe13__lane18_strm1_data_mask  ),      

               // PE 13, Lane 19                 
               .pe13__std__lane19_strm0_ready         ( pe13__std__lane19_strm0_ready      ),      
               .std__pe13__lane19_strm0_cntl          ( std__pe13__lane19_strm0_cntl       ),      
               .std__pe13__lane19_strm0_data          ( std__pe13__lane19_strm0_data       ),      
               .std__pe13__lane19_strm0_data_valid    ( std__pe13__lane19_strm0_data_valid ),      
               .std__pe13__lane19_strm0_data_mask     ( std__pe13__lane19_strm0_data_mask  ),      

               .pe13__std__lane19_strm1_ready         ( pe13__std__lane19_strm1_ready      ),      
               .std__pe13__lane19_strm1_cntl          ( std__pe13__lane19_strm1_cntl       ),      
               .std__pe13__lane19_strm1_data          ( std__pe13__lane19_strm1_data       ),      
               .std__pe13__lane19_strm1_data_valid    ( std__pe13__lane19_strm1_data_valid ),      
               .std__pe13__lane19_strm1_data_mask     ( std__pe13__lane19_strm1_data_mask  ),      

               // PE 13, Lane 20                 
               .pe13__std__lane20_strm0_ready         ( pe13__std__lane20_strm0_ready      ),      
               .std__pe13__lane20_strm0_cntl          ( std__pe13__lane20_strm0_cntl       ),      
               .std__pe13__lane20_strm0_data          ( std__pe13__lane20_strm0_data       ),      
               .std__pe13__lane20_strm0_data_valid    ( std__pe13__lane20_strm0_data_valid ),      
               .std__pe13__lane20_strm0_data_mask     ( std__pe13__lane20_strm0_data_mask  ),      

               .pe13__std__lane20_strm1_ready         ( pe13__std__lane20_strm1_ready      ),      
               .std__pe13__lane20_strm1_cntl          ( std__pe13__lane20_strm1_cntl       ),      
               .std__pe13__lane20_strm1_data          ( std__pe13__lane20_strm1_data       ),      
               .std__pe13__lane20_strm1_data_valid    ( std__pe13__lane20_strm1_data_valid ),      
               .std__pe13__lane20_strm1_data_mask     ( std__pe13__lane20_strm1_data_mask  ),      

               // PE 13, Lane 21                 
               .pe13__std__lane21_strm0_ready         ( pe13__std__lane21_strm0_ready      ),      
               .std__pe13__lane21_strm0_cntl          ( std__pe13__lane21_strm0_cntl       ),      
               .std__pe13__lane21_strm0_data          ( std__pe13__lane21_strm0_data       ),      
               .std__pe13__lane21_strm0_data_valid    ( std__pe13__lane21_strm0_data_valid ),      
               .std__pe13__lane21_strm0_data_mask     ( std__pe13__lane21_strm0_data_mask  ),      

               .pe13__std__lane21_strm1_ready         ( pe13__std__lane21_strm1_ready      ),      
               .std__pe13__lane21_strm1_cntl          ( std__pe13__lane21_strm1_cntl       ),      
               .std__pe13__lane21_strm1_data          ( std__pe13__lane21_strm1_data       ),      
               .std__pe13__lane21_strm1_data_valid    ( std__pe13__lane21_strm1_data_valid ),      
               .std__pe13__lane21_strm1_data_mask     ( std__pe13__lane21_strm1_data_mask  ),      

               // PE 13, Lane 22                 
               .pe13__std__lane22_strm0_ready         ( pe13__std__lane22_strm0_ready      ),      
               .std__pe13__lane22_strm0_cntl          ( std__pe13__lane22_strm0_cntl       ),      
               .std__pe13__lane22_strm0_data          ( std__pe13__lane22_strm0_data       ),      
               .std__pe13__lane22_strm0_data_valid    ( std__pe13__lane22_strm0_data_valid ),      
               .std__pe13__lane22_strm0_data_mask     ( std__pe13__lane22_strm0_data_mask  ),      

               .pe13__std__lane22_strm1_ready         ( pe13__std__lane22_strm1_ready      ),      
               .std__pe13__lane22_strm1_cntl          ( std__pe13__lane22_strm1_cntl       ),      
               .std__pe13__lane22_strm1_data          ( std__pe13__lane22_strm1_data       ),      
               .std__pe13__lane22_strm1_data_valid    ( std__pe13__lane22_strm1_data_valid ),      
               .std__pe13__lane22_strm1_data_mask     ( std__pe13__lane22_strm1_data_mask  ),      

               // PE 13, Lane 23                 
               .pe13__std__lane23_strm0_ready         ( pe13__std__lane23_strm0_ready      ),      
               .std__pe13__lane23_strm0_cntl          ( std__pe13__lane23_strm0_cntl       ),      
               .std__pe13__lane23_strm0_data          ( std__pe13__lane23_strm0_data       ),      
               .std__pe13__lane23_strm0_data_valid    ( std__pe13__lane23_strm0_data_valid ),      
               .std__pe13__lane23_strm0_data_mask     ( std__pe13__lane23_strm0_data_mask  ),      

               .pe13__std__lane23_strm1_ready         ( pe13__std__lane23_strm1_ready      ),      
               .std__pe13__lane23_strm1_cntl          ( std__pe13__lane23_strm1_cntl       ),      
               .std__pe13__lane23_strm1_data          ( std__pe13__lane23_strm1_data       ),      
               .std__pe13__lane23_strm1_data_valid    ( std__pe13__lane23_strm1_data_valid ),      
               .std__pe13__lane23_strm1_data_mask     ( std__pe13__lane23_strm1_data_mask  ),      

               // PE 13, Lane 24                 
               .pe13__std__lane24_strm0_ready         ( pe13__std__lane24_strm0_ready      ),      
               .std__pe13__lane24_strm0_cntl          ( std__pe13__lane24_strm0_cntl       ),      
               .std__pe13__lane24_strm0_data          ( std__pe13__lane24_strm0_data       ),      
               .std__pe13__lane24_strm0_data_valid    ( std__pe13__lane24_strm0_data_valid ),      
               .std__pe13__lane24_strm0_data_mask     ( std__pe13__lane24_strm0_data_mask  ),      

               .pe13__std__lane24_strm1_ready         ( pe13__std__lane24_strm1_ready      ),      
               .std__pe13__lane24_strm1_cntl          ( std__pe13__lane24_strm1_cntl       ),      
               .std__pe13__lane24_strm1_data          ( std__pe13__lane24_strm1_data       ),      
               .std__pe13__lane24_strm1_data_valid    ( std__pe13__lane24_strm1_data_valid ),      
               .std__pe13__lane24_strm1_data_mask     ( std__pe13__lane24_strm1_data_mask  ),      

               // PE 13, Lane 25                 
               .pe13__std__lane25_strm0_ready         ( pe13__std__lane25_strm0_ready      ),      
               .std__pe13__lane25_strm0_cntl          ( std__pe13__lane25_strm0_cntl       ),      
               .std__pe13__lane25_strm0_data          ( std__pe13__lane25_strm0_data       ),      
               .std__pe13__lane25_strm0_data_valid    ( std__pe13__lane25_strm0_data_valid ),      
               .std__pe13__lane25_strm0_data_mask     ( std__pe13__lane25_strm0_data_mask  ),      

               .pe13__std__lane25_strm1_ready         ( pe13__std__lane25_strm1_ready      ),      
               .std__pe13__lane25_strm1_cntl          ( std__pe13__lane25_strm1_cntl       ),      
               .std__pe13__lane25_strm1_data          ( std__pe13__lane25_strm1_data       ),      
               .std__pe13__lane25_strm1_data_valid    ( std__pe13__lane25_strm1_data_valid ),      
               .std__pe13__lane25_strm1_data_mask     ( std__pe13__lane25_strm1_data_mask  ),      

               // PE 13, Lane 26                 
               .pe13__std__lane26_strm0_ready         ( pe13__std__lane26_strm0_ready      ),      
               .std__pe13__lane26_strm0_cntl          ( std__pe13__lane26_strm0_cntl       ),      
               .std__pe13__lane26_strm0_data          ( std__pe13__lane26_strm0_data       ),      
               .std__pe13__lane26_strm0_data_valid    ( std__pe13__lane26_strm0_data_valid ),      
               .std__pe13__lane26_strm0_data_mask     ( std__pe13__lane26_strm0_data_mask  ),      

               .pe13__std__lane26_strm1_ready         ( pe13__std__lane26_strm1_ready      ),      
               .std__pe13__lane26_strm1_cntl          ( std__pe13__lane26_strm1_cntl       ),      
               .std__pe13__lane26_strm1_data          ( std__pe13__lane26_strm1_data       ),      
               .std__pe13__lane26_strm1_data_valid    ( std__pe13__lane26_strm1_data_valid ),      
               .std__pe13__lane26_strm1_data_mask     ( std__pe13__lane26_strm1_data_mask  ),      

               // PE 13, Lane 27                 
               .pe13__std__lane27_strm0_ready         ( pe13__std__lane27_strm0_ready      ),      
               .std__pe13__lane27_strm0_cntl          ( std__pe13__lane27_strm0_cntl       ),      
               .std__pe13__lane27_strm0_data          ( std__pe13__lane27_strm0_data       ),      
               .std__pe13__lane27_strm0_data_valid    ( std__pe13__lane27_strm0_data_valid ),      
               .std__pe13__lane27_strm0_data_mask     ( std__pe13__lane27_strm0_data_mask  ),      

               .pe13__std__lane27_strm1_ready         ( pe13__std__lane27_strm1_ready      ),      
               .std__pe13__lane27_strm1_cntl          ( std__pe13__lane27_strm1_cntl       ),      
               .std__pe13__lane27_strm1_data          ( std__pe13__lane27_strm1_data       ),      
               .std__pe13__lane27_strm1_data_valid    ( std__pe13__lane27_strm1_data_valid ),      
               .std__pe13__lane27_strm1_data_mask     ( std__pe13__lane27_strm1_data_mask  ),      

               // PE 13, Lane 28                 
               .pe13__std__lane28_strm0_ready         ( pe13__std__lane28_strm0_ready      ),      
               .std__pe13__lane28_strm0_cntl          ( std__pe13__lane28_strm0_cntl       ),      
               .std__pe13__lane28_strm0_data          ( std__pe13__lane28_strm0_data       ),      
               .std__pe13__lane28_strm0_data_valid    ( std__pe13__lane28_strm0_data_valid ),      
               .std__pe13__lane28_strm0_data_mask     ( std__pe13__lane28_strm0_data_mask  ),      

               .pe13__std__lane28_strm1_ready         ( pe13__std__lane28_strm1_ready      ),      
               .std__pe13__lane28_strm1_cntl          ( std__pe13__lane28_strm1_cntl       ),      
               .std__pe13__lane28_strm1_data          ( std__pe13__lane28_strm1_data       ),      
               .std__pe13__lane28_strm1_data_valid    ( std__pe13__lane28_strm1_data_valid ),      
               .std__pe13__lane28_strm1_data_mask     ( std__pe13__lane28_strm1_data_mask  ),      

               // PE 13, Lane 29                 
               .pe13__std__lane29_strm0_ready         ( pe13__std__lane29_strm0_ready      ),      
               .std__pe13__lane29_strm0_cntl          ( std__pe13__lane29_strm0_cntl       ),      
               .std__pe13__lane29_strm0_data          ( std__pe13__lane29_strm0_data       ),      
               .std__pe13__lane29_strm0_data_valid    ( std__pe13__lane29_strm0_data_valid ),      
               .std__pe13__lane29_strm0_data_mask     ( std__pe13__lane29_strm0_data_mask  ),      

               .pe13__std__lane29_strm1_ready         ( pe13__std__lane29_strm1_ready      ),      
               .std__pe13__lane29_strm1_cntl          ( std__pe13__lane29_strm1_cntl       ),      
               .std__pe13__lane29_strm1_data          ( std__pe13__lane29_strm1_data       ),      
               .std__pe13__lane29_strm1_data_valid    ( std__pe13__lane29_strm1_data_valid ),      
               .std__pe13__lane29_strm1_data_mask     ( std__pe13__lane29_strm1_data_mask  ),      

               // PE 13, Lane 30                 
               .pe13__std__lane30_strm0_ready         ( pe13__std__lane30_strm0_ready      ),      
               .std__pe13__lane30_strm0_cntl          ( std__pe13__lane30_strm0_cntl       ),      
               .std__pe13__lane30_strm0_data          ( std__pe13__lane30_strm0_data       ),      
               .std__pe13__lane30_strm0_data_valid    ( std__pe13__lane30_strm0_data_valid ),      
               .std__pe13__lane30_strm0_data_mask     ( std__pe13__lane30_strm0_data_mask  ),      

               .pe13__std__lane30_strm1_ready         ( pe13__std__lane30_strm1_ready      ),      
               .std__pe13__lane30_strm1_cntl          ( std__pe13__lane30_strm1_cntl       ),      
               .std__pe13__lane30_strm1_data          ( std__pe13__lane30_strm1_data       ),      
               .std__pe13__lane30_strm1_data_valid    ( std__pe13__lane30_strm1_data_valid ),      
               .std__pe13__lane30_strm1_data_mask     ( std__pe13__lane30_strm1_data_mask  ),      

               // PE 13, Lane 31                 
               .pe13__std__lane31_strm0_ready         ( pe13__std__lane31_strm0_ready      ),      
               .std__pe13__lane31_strm0_cntl          ( std__pe13__lane31_strm0_cntl       ),      
               .std__pe13__lane31_strm0_data          ( std__pe13__lane31_strm0_data       ),      
               .std__pe13__lane31_strm0_data_valid    ( std__pe13__lane31_strm0_data_valid ),      
               .std__pe13__lane31_strm0_data_mask     ( std__pe13__lane31_strm0_data_mask  ),      

               .pe13__std__lane31_strm1_ready         ( pe13__std__lane31_strm1_ready      ),      
               .std__pe13__lane31_strm1_cntl          ( std__pe13__lane31_strm1_cntl       ),      
               .std__pe13__lane31_strm1_data          ( std__pe13__lane31_strm1_data       ),      
               .std__pe13__lane31_strm1_data_valid    ( std__pe13__lane31_strm1_data_valid ),      
               .std__pe13__lane31_strm1_data_mask     ( std__pe13__lane31_strm1_data_mask  ),      

               // PE 14, Lane 0                 
               .pe14__std__lane0_strm0_ready         ( pe14__std__lane0_strm0_ready      ),      
               .std__pe14__lane0_strm0_cntl          ( std__pe14__lane0_strm0_cntl       ),      
               .std__pe14__lane0_strm0_data          ( std__pe14__lane0_strm0_data       ),      
               .std__pe14__lane0_strm0_data_valid    ( std__pe14__lane0_strm0_data_valid ),      
               .std__pe14__lane0_strm0_data_mask     ( std__pe14__lane0_strm0_data_mask  ),      

               .pe14__std__lane0_strm1_ready         ( pe14__std__lane0_strm1_ready      ),      
               .std__pe14__lane0_strm1_cntl          ( std__pe14__lane0_strm1_cntl       ),      
               .std__pe14__lane0_strm1_data          ( std__pe14__lane0_strm1_data       ),      
               .std__pe14__lane0_strm1_data_valid    ( std__pe14__lane0_strm1_data_valid ),      
               .std__pe14__lane0_strm1_data_mask     ( std__pe14__lane0_strm1_data_mask  ),      

               // PE 14, Lane 1                 
               .pe14__std__lane1_strm0_ready         ( pe14__std__lane1_strm0_ready      ),      
               .std__pe14__lane1_strm0_cntl          ( std__pe14__lane1_strm0_cntl       ),      
               .std__pe14__lane1_strm0_data          ( std__pe14__lane1_strm0_data       ),      
               .std__pe14__lane1_strm0_data_valid    ( std__pe14__lane1_strm0_data_valid ),      
               .std__pe14__lane1_strm0_data_mask     ( std__pe14__lane1_strm0_data_mask  ),      

               .pe14__std__lane1_strm1_ready         ( pe14__std__lane1_strm1_ready      ),      
               .std__pe14__lane1_strm1_cntl          ( std__pe14__lane1_strm1_cntl       ),      
               .std__pe14__lane1_strm1_data          ( std__pe14__lane1_strm1_data       ),      
               .std__pe14__lane1_strm1_data_valid    ( std__pe14__lane1_strm1_data_valid ),      
               .std__pe14__lane1_strm1_data_mask     ( std__pe14__lane1_strm1_data_mask  ),      

               // PE 14, Lane 2                 
               .pe14__std__lane2_strm0_ready         ( pe14__std__lane2_strm0_ready      ),      
               .std__pe14__lane2_strm0_cntl          ( std__pe14__lane2_strm0_cntl       ),      
               .std__pe14__lane2_strm0_data          ( std__pe14__lane2_strm0_data       ),      
               .std__pe14__lane2_strm0_data_valid    ( std__pe14__lane2_strm0_data_valid ),      
               .std__pe14__lane2_strm0_data_mask     ( std__pe14__lane2_strm0_data_mask  ),      

               .pe14__std__lane2_strm1_ready         ( pe14__std__lane2_strm1_ready      ),      
               .std__pe14__lane2_strm1_cntl          ( std__pe14__lane2_strm1_cntl       ),      
               .std__pe14__lane2_strm1_data          ( std__pe14__lane2_strm1_data       ),      
               .std__pe14__lane2_strm1_data_valid    ( std__pe14__lane2_strm1_data_valid ),      
               .std__pe14__lane2_strm1_data_mask     ( std__pe14__lane2_strm1_data_mask  ),      

               // PE 14, Lane 3                 
               .pe14__std__lane3_strm0_ready         ( pe14__std__lane3_strm0_ready      ),      
               .std__pe14__lane3_strm0_cntl          ( std__pe14__lane3_strm0_cntl       ),      
               .std__pe14__lane3_strm0_data          ( std__pe14__lane3_strm0_data       ),      
               .std__pe14__lane3_strm0_data_valid    ( std__pe14__lane3_strm0_data_valid ),      
               .std__pe14__lane3_strm0_data_mask     ( std__pe14__lane3_strm0_data_mask  ),      

               .pe14__std__lane3_strm1_ready         ( pe14__std__lane3_strm1_ready      ),      
               .std__pe14__lane3_strm1_cntl          ( std__pe14__lane3_strm1_cntl       ),      
               .std__pe14__lane3_strm1_data          ( std__pe14__lane3_strm1_data       ),      
               .std__pe14__lane3_strm1_data_valid    ( std__pe14__lane3_strm1_data_valid ),      
               .std__pe14__lane3_strm1_data_mask     ( std__pe14__lane3_strm1_data_mask  ),      

               // PE 14, Lane 4                 
               .pe14__std__lane4_strm0_ready         ( pe14__std__lane4_strm0_ready      ),      
               .std__pe14__lane4_strm0_cntl          ( std__pe14__lane4_strm0_cntl       ),      
               .std__pe14__lane4_strm0_data          ( std__pe14__lane4_strm0_data       ),      
               .std__pe14__lane4_strm0_data_valid    ( std__pe14__lane4_strm0_data_valid ),      
               .std__pe14__lane4_strm0_data_mask     ( std__pe14__lane4_strm0_data_mask  ),      

               .pe14__std__lane4_strm1_ready         ( pe14__std__lane4_strm1_ready      ),      
               .std__pe14__lane4_strm1_cntl          ( std__pe14__lane4_strm1_cntl       ),      
               .std__pe14__lane4_strm1_data          ( std__pe14__lane4_strm1_data       ),      
               .std__pe14__lane4_strm1_data_valid    ( std__pe14__lane4_strm1_data_valid ),      
               .std__pe14__lane4_strm1_data_mask     ( std__pe14__lane4_strm1_data_mask  ),      

               // PE 14, Lane 5                 
               .pe14__std__lane5_strm0_ready         ( pe14__std__lane5_strm0_ready      ),      
               .std__pe14__lane5_strm0_cntl          ( std__pe14__lane5_strm0_cntl       ),      
               .std__pe14__lane5_strm0_data          ( std__pe14__lane5_strm0_data       ),      
               .std__pe14__lane5_strm0_data_valid    ( std__pe14__lane5_strm0_data_valid ),      
               .std__pe14__lane5_strm0_data_mask     ( std__pe14__lane5_strm0_data_mask  ),      

               .pe14__std__lane5_strm1_ready         ( pe14__std__lane5_strm1_ready      ),      
               .std__pe14__lane5_strm1_cntl          ( std__pe14__lane5_strm1_cntl       ),      
               .std__pe14__lane5_strm1_data          ( std__pe14__lane5_strm1_data       ),      
               .std__pe14__lane5_strm1_data_valid    ( std__pe14__lane5_strm1_data_valid ),      
               .std__pe14__lane5_strm1_data_mask     ( std__pe14__lane5_strm1_data_mask  ),      

               // PE 14, Lane 6                 
               .pe14__std__lane6_strm0_ready         ( pe14__std__lane6_strm0_ready      ),      
               .std__pe14__lane6_strm0_cntl          ( std__pe14__lane6_strm0_cntl       ),      
               .std__pe14__lane6_strm0_data          ( std__pe14__lane6_strm0_data       ),      
               .std__pe14__lane6_strm0_data_valid    ( std__pe14__lane6_strm0_data_valid ),      
               .std__pe14__lane6_strm0_data_mask     ( std__pe14__lane6_strm0_data_mask  ),      

               .pe14__std__lane6_strm1_ready         ( pe14__std__lane6_strm1_ready      ),      
               .std__pe14__lane6_strm1_cntl          ( std__pe14__lane6_strm1_cntl       ),      
               .std__pe14__lane6_strm1_data          ( std__pe14__lane6_strm1_data       ),      
               .std__pe14__lane6_strm1_data_valid    ( std__pe14__lane6_strm1_data_valid ),      
               .std__pe14__lane6_strm1_data_mask     ( std__pe14__lane6_strm1_data_mask  ),      

               // PE 14, Lane 7                 
               .pe14__std__lane7_strm0_ready         ( pe14__std__lane7_strm0_ready      ),      
               .std__pe14__lane7_strm0_cntl          ( std__pe14__lane7_strm0_cntl       ),      
               .std__pe14__lane7_strm0_data          ( std__pe14__lane7_strm0_data       ),      
               .std__pe14__lane7_strm0_data_valid    ( std__pe14__lane7_strm0_data_valid ),      
               .std__pe14__lane7_strm0_data_mask     ( std__pe14__lane7_strm0_data_mask  ),      

               .pe14__std__lane7_strm1_ready         ( pe14__std__lane7_strm1_ready      ),      
               .std__pe14__lane7_strm1_cntl          ( std__pe14__lane7_strm1_cntl       ),      
               .std__pe14__lane7_strm1_data          ( std__pe14__lane7_strm1_data       ),      
               .std__pe14__lane7_strm1_data_valid    ( std__pe14__lane7_strm1_data_valid ),      
               .std__pe14__lane7_strm1_data_mask     ( std__pe14__lane7_strm1_data_mask  ),      

               // PE 14, Lane 8                 
               .pe14__std__lane8_strm0_ready         ( pe14__std__lane8_strm0_ready      ),      
               .std__pe14__lane8_strm0_cntl          ( std__pe14__lane8_strm0_cntl       ),      
               .std__pe14__lane8_strm0_data          ( std__pe14__lane8_strm0_data       ),      
               .std__pe14__lane8_strm0_data_valid    ( std__pe14__lane8_strm0_data_valid ),      
               .std__pe14__lane8_strm0_data_mask     ( std__pe14__lane8_strm0_data_mask  ),      

               .pe14__std__lane8_strm1_ready         ( pe14__std__lane8_strm1_ready      ),      
               .std__pe14__lane8_strm1_cntl          ( std__pe14__lane8_strm1_cntl       ),      
               .std__pe14__lane8_strm1_data          ( std__pe14__lane8_strm1_data       ),      
               .std__pe14__lane8_strm1_data_valid    ( std__pe14__lane8_strm1_data_valid ),      
               .std__pe14__lane8_strm1_data_mask     ( std__pe14__lane8_strm1_data_mask  ),      

               // PE 14, Lane 9                 
               .pe14__std__lane9_strm0_ready         ( pe14__std__lane9_strm0_ready      ),      
               .std__pe14__lane9_strm0_cntl          ( std__pe14__lane9_strm0_cntl       ),      
               .std__pe14__lane9_strm0_data          ( std__pe14__lane9_strm0_data       ),      
               .std__pe14__lane9_strm0_data_valid    ( std__pe14__lane9_strm0_data_valid ),      
               .std__pe14__lane9_strm0_data_mask     ( std__pe14__lane9_strm0_data_mask  ),      

               .pe14__std__lane9_strm1_ready         ( pe14__std__lane9_strm1_ready      ),      
               .std__pe14__lane9_strm1_cntl          ( std__pe14__lane9_strm1_cntl       ),      
               .std__pe14__lane9_strm1_data          ( std__pe14__lane9_strm1_data       ),      
               .std__pe14__lane9_strm1_data_valid    ( std__pe14__lane9_strm1_data_valid ),      
               .std__pe14__lane9_strm1_data_mask     ( std__pe14__lane9_strm1_data_mask  ),      

               // PE 14, Lane 10                 
               .pe14__std__lane10_strm0_ready         ( pe14__std__lane10_strm0_ready      ),      
               .std__pe14__lane10_strm0_cntl          ( std__pe14__lane10_strm0_cntl       ),      
               .std__pe14__lane10_strm0_data          ( std__pe14__lane10_strm0_data       ),      
               .std__pe14__lane10_strm0_data_valid    ( std__pe14__lane10_strm0_data_valid ),      
               .std__pe14__lane10_strm0_data_mask     ( std__pe14__lane10_strm0_data_mask  ),      

               .pe14__std__lane10_strm1_ready         ( pe14__std__lane10_strm1_ready      ),      
               .std__pe14__lane10_strm1_cntl          ( std__pe14__lane10_strm1_cntl       ),      
               .std__pe14__lane10_strm1_data          ( std__pe14__lane10_strm1_data       ),      
               .std__pe14__lane10_strm1_data_valid    ( std__pe14__lane10_strm1_data_valid ),      
               .std__pe14__lane10_strm1_data_mask     ( std__pe14__lane10_strm1_data_mask  ),      

               // PE 14, Lane 11                 
               .pe14__std__lane11_strm0_ready         ( pe14__std__lane11_strm0_ready      ),      
               .std__pe14__lane11_strm0_cntl          ( std__pe14__lane11_strm0_cntl       ),      
               .std__pe14__lane11_strm0_data          ( std__pe14__lane11_strm0_data       ),      
               .std__pe14__lane11_strm0_data_valid    ( std__pe14__lane11_strm0_data_valid ),      
               .std__pe14__lane11_strm0_data_mask     ( std__pe14__lane11_strm0_data_mask  ),      

               .pe14__std__lane11_strm1_ready         ( pe14__std__lane11_strm1_ready      ),      
               .std__pe14__lane11_strm1_cntl          ( std__pe14__lane11_strm1_cntl       ),      
               .std__pe14__lane11_strm1_data          ( std__pe14__lane11_strm1_data       ),      
               .std__pe14__lane11_strm1_data_valid    ( std__pe14__lane11_strm1_data_valid ),      
               .std__pe14__lane11_strm1_data_mask     ( std__pe14__lane11_strm1_data_mask  ),      

               // PE 14, Lane 12                 
               .pe14__std__lane12_strm0_ready         ( pe14__std__lane12_strm0_ready      ),      
               .std__pe14__lane12_strm0_cntl          ( std__pe14__lane12_strm0_cntl       ),      
               .std__pe14__lane12_strm0_data          ( std__pe14__lane12_strm0_data       ),      
               .std__pe14__lane12_strm0_data_valid    ( std__pe14__lane12_strm0_data_valid ),      
               .std__pe14__lane12_strm0_data_mask     ( std__pe14__lane12_strm0_data_mask  ),      

               .pe14__std__lane12_strm1_ready         ( pe14__std__lane12_strm1_ready      ),      
               .std__pe14__lane12_strm1_cntl          ( std__pe14__lane12_strm1_cntl       ),      
               .std__pe14__lane12_strm1_data          ( std__pe14__lane12_strm1_data       ),      
               .std__pe14__lane12_strm1_data_valid    ( std__pe14__lane12_strm1_data_valid ),      
               .std__pe14__lane12_strm1_data_mask     ( std__pe14__lane12_strm1_data_mask  ),      

               // PE 14, Lane 13                 
               .pe14__std__lane13_strm0_ready         ( pe14__std__lane13_strm0_ready      ),      
               .std__pe14__lane13_strm0_cntl          ( std__pe14__lane13_strm0_cntl       ),      
               .std__pe14__lane13_strm0_data          ( std__pe14__lane13_strm0_data       ),      
               .std__pe14__lane13_strm0_data_valid    ( std__pe14__lane13_strm0_data_valid ),      
               .std__pe14__lane13_strm0_data_mask     ( std__pe14__lane13_strm0_data_mask  ),      

               .pe14__std__lane13_strm1_ready         ( pe14__std__lane13_strm1_ready      ),      
               .std__pe14__lane13_strm1_cntl          ( std__pe14__lane13_strm1_cntl       ),      
               .std__pe14__lane13_strm1_data          ( std__pe14__lane13_strm1_data       ),      
               .std__pe14__lane13_strm1_data_valid    ( std__pe14__lane13_strm1_data_valid ),      
               .std__pe14__lane13_strm1_data_mask     ( std__pe14__lane13_strm1_data_mask  ),      

               // PE 14, Lane 14                 
               .pe14__std__lane14_strm0_ready         ( pe14__std__lane14_strm0_ready      ),      
               .std__pe14__lane14_strm0_cntl          ( std__pe14__lane14_strm0_cntl       ),      
               .std__pe14__lane14_strm0_data          ( std__pe14__lane14_strm0_data       ),      
               .std__pe14__lane14_strm0_data_valid    ( std__pe14__lane14_strm0_data_valid ),      
               .std__pe14__lane14_strm0_data_mask     ( std__pe14__lane14_strm0_data_mask  ),      

               .pe14__std__lane14_strm1_ready         ( pe14__std__lane14_strm1_ready      ),      
               .std__pe14__lane14_strm1_cntl          ( std__pe14__lane14_strm1_cntl       ),      
               .std__pe14__lane14_strm1_data          ( std__pe14__lane14_strm1_data       ),      
               .std__pe14__lane14_strm1_data_valid    ( std__pe14__lane14_strm1_data_valid ),      
               .std__pe14__lane14_strm1_data_mask     ( std__pe14__lane14_strm1_data_mask  ),      

               // PE 14, Lane 15                 
               .pe14__std__lane15_strm0_ready         ( pe14__std__lane15_strm0_ready      ),      
               .std__pe14__lane15_strm0_cntl          ( std__pe14__lane15_strm0_cntl       ),      
               .std__pe14__lane15_strm0_data          ( std__pe14__lane15_strm0_data       ),      
               .std__pe14__lane15_strm0_data_valid    ( std__pe14__lane15_strm0_data_valid ),      
               .std__pe14__lane15_strm0_data_mask     ( std__pe14__lane15_strm0_data_mask  ),      

               .pe14__std__lane15_strm1_ready         ( pe14__std__lane15_strm1_ready      ),      
               .std__pe14__lane15_strm1_cntl          ( std__pe14__lane15_strm1_cntl       ),      
               .std__pe14__lane15_strm1_data          ( std__pe14__lane15_strm1_data       ),      
               .std__pe14__lane15_strm1_data_valid    ( std__pe14__lane15_strm1_data_valid ),      
               .std__pe14__lane15_strm1_data_mask     ( std__pe14__lane15_strm1_data_mask  ),      

               // PE 14, Lane 16                 
               .pe14__std__lane16_strm0_ready         ( pe14__std__lane16_strm0_ready      ),      
               .std__pe14__lane16_strm0_cntl          ( std__pe14__lane16_strm0_cntl       ),      
               .std__pe14__lane16_strm0_data          ( std__pe14__lane16_strm0_data       ),      
               .std__pe14__lane16_strm0_data_valid    ( std__pe14__lane16_strm0_data_valid ),      
               .std__pe14__lane16_strm0_data_mask     ( std__pe14__lane16_strm0_data_mask  ),      

               .pe14__std__lane16_strm1_ready         ( pe14__std__lane16_strm1_ready      ),      
               .std__pe14__lane16_strm1_cntl          ( std__pe14__lane16_strm1_cntl       ),      
               .std__pe14__lane16_strm1_data          ( std__pe14__lane16_strm1_data       ),      
               .std__pe14__lane16_strm1_data_valid    ( std__pe14__lane16_strm1_data_valid ),      
               .std__pe14__lane16_strm1_data_mask     ( std__pe14__lane16_strm1_data_mask  ),      

               // PE 14, Lane 17                 
               .pe14__std__lane17_strm0_ready         ( pe14__std__lane17_strm0_ready      ),      
               .std__pe14__lane17_strm0_cntl          ( std__pe14__lane17_strm0_cntl       ),      
               .std__pe14__lane17_strm0_data          ( std__pe14__lane17_strm0_data       ),      
               .std__pe14__lane17_strm0_data_valid    ( std__pe14__lane17_strm0_data_valid ),      
               .std__pe14__lane17_strm0_data_mask     ( std__pe14__lane17_strm0_data_mask  ),      

               .pe14__std__lane17_strm1_ready         ( pe14__std__lane17_strm1_ready      ),      
               .std__pe14__lane17_strm1_cntl          ( std__pe14__lane17_strm1_cntl       ),      
               .std__pe14__lane17_strm1_data          ( std__pe14__lane17_strm1_data       ),      
               .std__pe14__lane17_strm1_data_valid    ( std__pe14__lane17_strm1_data_valid ),      
               .std__pe14__lane17_strm1_data_mask     ( std__pe14__lane17_strm1_data_mask  ),      

               // PE 14, Lane 18                 
               .pe14__std__lane18_strm0_ready         ( pe14__std__lane18_strm0_ready      ),      
               .std__pe14__lane18_strm0_cntl          ( std__pe14__lane18_strm0_cntl       ),      
               .std__pe14__lane18_strm0_data          ( std__pe14__lane18_strm0_data       ),      
               .std__pe14__lane18_strm0_data_valid    ( std__pe14__lane18_strm0_data_valid ),      
               .std__pe14__lane18_strm0_data_mask     ( std__pe14__lane18_strm0_data_mask  ),      

               .pe14__std__lane18_strm1_ready         ( pe14__std__lane18_strm1_ready      ),      
               .std__pe14__lane18_strm1_cntl          ( std__pe14__lane18_strm1_cntl       ),      
               .std__pe14__lane18_strm1_data          ( std__pe14__lane18_strm1_data       ),      
               .std__pe14__lane18_strm1_data_valid    ( std__pe14__lane18_strm1_data_valid ),      
               .std__pe14__lane18_strm1_data_mask     ( std__pe14__lane18_strm1_data_mask  ),      

               // PE 14, Lane 19                 
               .pe14__std__lane19_strm0_ready         ( pe14__std__lane19_strm0_ready      ),      
               .std__pe14__lane19_strm0_cntl          ( std__pe14__lane19_strm0_cntl       ),      
               .std__pe14__lane19_strm0_data          ( std__pe14__lane19_strm0_data       ),      
               .std__pe14__lane19_strm0_data_valid    ( std__pe14__lane19_strm0_data_valid ),      
               .std__pe14__lane19_strm0_data_mask     ( std__pe14__lane19_strm0_data_mask  ),      

               .pe14__std__lane19_strm1_ready         ( pe14__std__lane19_strm1_ready      ),      
               .std__pe14__lane19_strm1_cntl          ( std__pe14__lane19_strm1_cntl       ),      
               .std__pe14__lane19_strm1_data          ( std__pe14__lane19_strm1_data       ),      
               .std__pe14__lane19_strm1_data_valid    ( std__pe14__lane19_strm1_data_valid ),      
               .std__pe14__lane19_strm1_data_mask     ( std__pe14__lane19_strm1_data_mask  ),      

               // PE 14, Lane 20                 
               .pe14__std__lane20_strm0_ready         ( pe14__std__lane20_strm0_ready      ),      
               .std__pe14__lane20_strm0_cntl          ( std__pe14__lane20_strm0_cntl       ),      
               .std__pe14__lane20_strm0_data          ( std__pe14__lane20_strm0_data       ),      
               .std__pe14__lane20_strm0_data_valid    ( std__pe14__lane20_strm0_data_valid ),      
               .std__pe14__lane20_strm0_data_mask     ( std__pe14__lane20_strm0_data_mask  ),      

               .pe14__std__lane20_strm1_ready         ( pe14__std__lane20_strm1_ready      ),      
               .std__pe14__lane20_strm1_cntl          ( std__pe14__lane20_strm1_cntl       ),      
               .std__pe14__lane20_strm1_data          ( std__pe14__lane20_strm1_data       ),      
               .std__pe14__lane20_strm1_data_valid    ( std__pe14__lane20_strm1_data_valid ),      
               .std__pe14__lane20_strm1_data_mask     ( std__pe14__lane20_strm1_data_mask  ),      

               // PE 14, Lane 21                 
               .pe14__std__lane21_strm0_ready         ( pe14__std__lane21_strm0_ready      ),      
               .std__pe14__lane21_strm0_cntl          ( std__pe14__lane21_strm0_cntl       ),      
               .std__pe14__lane21_strm0_data          ( std__pe14__lane21_strm0_data       ),      
               .std__pe14__lane21_strm0_data_valid    ( std__pe14__lane21_strm0_data_valid ),      
               .std__pe14__lane21_strm0_data_mask     ( std__pe14__lane21_strm0_data_mask  ),      

               .pe14__std__lane21_strm1_ready         ( pe14__std__lane21_strm1_ready      ),      
               .std__pe14__lane21_strm1_cntl          ( std__pe14__lane21_strm1_cntl       ),      
               .std__pe14__lane21_strm1_data          ( std__pe14__lane21_strm1_data       ),      
               .std__pe14__lane21_strm1_data_valid    ( std__pe14__lane21_strm1_data_valid ),      
               .std__pe14__lane21_strm1_data_mask     ( std__pe14__lane21_strm1_data_mask  ),      

               // PE 14, Lane 22                 
               .pe14__std__lane22_strm0_ready         ( pe14__std__lane22_strm0_ready      ),      
               .std__pe14__lane22_strm0_cntl          ( std__pe14__lane22_strm0_cntl       ),      
               .std__pe14__lane22_strm0_data          ( std__pe14__lane22_strm0_data       ),      
               .std__pe14__lane22_strm0_data_valid    ( std__pe14__lane22_strm0_data_valid ),      
               .std__pe14__lane22_strm0_data_mask     ( std__pe14__lane22_strm0_data_mask  ),      

               .pe14__std__lane22_strm1_ready         ( pe14__std__lane22_strm1_ready      ),      
               .std__pe14__lane22_strm1_cntl          ( std__pe14__lane22_strm1_cntl       ),      
               .std__pe14__lane22_strm1_data          ( std__pe14__lane22_strm1_data       ),      
               .std__pe14__lane22_strm1_data_valid    ( std__pe14__lane22_strm1_data_valid ),      
               .std__pe14__lane22_strm1_data_mask     ( std__pe14__lane22_strm1_data_mask  ),      

               // PE 14, Lane 23                 
               .pe14__std__lane23_strm0_ready         ( pe14__std__lane23_strm0_ready      ),      
               .std__pe14__lane23_strm0_cntl          ( std__pe14__lane23_strm0_cntl       ),      
               .std__pe14__lane23_strm0_data          ( std__pe14__lane23_strm0_data       ),      
               .std__pe14__lane23_strm0_data_valid    ( std__pe14__lane23_strm0_data_valid ),      
               .std__pe14__lane23_strm0_data_mask     ( std__pe14__lane23_strm0_data_mask  ),      

               .pe14__std__lane23_strm1_ready         ( pe14__std__lane23_strm1_ready      ),      
               .std__pe14__lane23_strm1_cntl          ( std__pe14__lane23_strm1_cntl       ),      
               .std__pe14__lane23_strm1_data          ( std__pe14__lane23_strm1_data       ),      
               .std__pe14__lane23_strm1_data_valid    ( std__pe14__lane23_strm1_data_valid ),      
               .std__pe14__lane23_strm1_data_mask     ( std__pe14__lane23_strm1_data_mask  ),      

               // PE 14, Lane 24                 
               .pe14__std__lane24_strm0_ready         ( pe14__std__lane24_strm0_ready      ),      
               .std__pe14__lane24_strm0_cntl          ( std__pe14__lane24_strm0_cntl       ),      
               .std__pe14__lane24_strm0_data          ( std__pe14__lane24_strm0_data       ),      
               .std__pe14__lane24_strm0_data_valid    ( std__pe14__lane24_strm0_data_valid ),      
               .std__pe14__lane24_strm0_data_mask     ( std__pe14__lane24_strm0_data_mask  ),      

               .pe14__std__lane24_strm1_ready         ( pe14__std__lane24_strm1_ready      ),      
               .std__pe14__lane24_strm1_cntl          ( std__pe14__lane24_strm1_cntl       ),      
               .std__pe14__lane24_strm1_data          ( std__pe14__lane24_strm1_data       ),      
               .std__pe14__lane24_strm1_data_valid    ( std__pe14__lane24_strm1_data_valid ),      
               .std__pe14__lane24_strm1_data_mask     ( std__pe14__lane24_strm1_data_mask  ),      

               // PE 14, Lane 25                 
               .pe14__std__lane25_strm0_ready         ( pe14__std__lane25_strm0_ready      ),      
               .std__pe14__lane25_strm0_cntl          ( std__pe14__lane25_strm0_cntl       ),      
               .std__pe14__lane25_strm0_data          ( std__pe14__lane25_strm0_data       ),      
               .std__pe14__lane25_strm0_data_valid    ( std__pe14__lane25_strm0_data_valid ),      
               .std__pe14__lane25_strm0_data_mask     ( std__pe14__lane25_strm0_data_mask  ),      

               .pe14__std__lane25_strm1_ready         ( pe14__std__lane25_strm1_ready      ),      
               .std__pe14__lane25_strm1_cntl          ( std__pe14__lane25_strm1_cntl       ),      
               .std__pe14__lane25_strm1_data          ( std__pe14__lane25_strm1_data       ),      
               .std__pe14__lane25_strm1_data_valid    ( std__pe14__lane25_strm1_data_valid ),      
               .std__pe14__lane25_strm1_data_mask     ( std__pe14__lane25_strm1_data_mask  ),      

               // PE 14, Lane 26                 
               .pe14__std__lane26_strm0_ready         ( pe14__std__lane26_strm0_ready      ),      
               .std__pe14__lane26_strm0_cntl          ( std__pe14__lane26_strm0_cntl       ),      
               .std__pe14__lane26_strm0_data          ( std__pe14__lane26_strm0_data       ),      
               .std__pe14__lane26_strm0_data_valid    ( std__pe14__lane26_strm0_data_valid ),      
               .std__pe14__lane26_strm0_data_mask     ( std__pe14__lane26_strm0_data_mask  ),      

               .pe14__std__lane26_strm1_ready         ( pe14__std__lane26_strm1_ready      ),      
               .std__pe14__lane26_strm1_cntl          ( std__pe14__lane26_strm1_cntl       ),      
               .std__pe14__lane26_strm1_data          ( std__pe14__lane26_strm1_data       ),      
               .std__pe14__lane26_strm1_data_valid    ( std__pe14__lane26_strm1_data_valid ),      
               .std__pe14__lane26_strm1_data_mask     ( std__pe14__lane26_strm1_data_mask  ),      

               // PE 14, Lane 27                 
               .pe14__std__lane27_strm0_ready         ( pe14__std__lane27_strm0_ready      ),      
               .std__pe14__lane27_strm0_cntl          ( std__pe14__lane27_strm0_cntl       ),      
               .std__pe14__lane27_strm0_data          ( std__pe14__lane27_strm0_data       ),      
               .std__pe14__lane27_strm0_data_valid    ( std__pe14__lane27_strm0_data_valid ),      
               .std__pe14__lane27_strm0_data_mask     ( std__pe14__lane27_strm0_data_mask  ),      

               .pe14__std__lane27_strm1_ready         ( pe14__std__lane27_strm1_ready      ),      
               .std__pe14__lane27_strm1_cntl          ( std__pe14__lane27_strm1_cntl       ),      
               .std__pe14__lane27_strm1_data          ( std__pe14__lane27_strm1_data       ),      
               .std__pe14__lane27_strm1_data_valid    ( std__pe14__lane27_strm1_data_valid ),      
               .std__pe14__lane27_strm1_data_mask     ( std__pe14__lane27_strm1_data_mask  ),      

               // PE 14, Lane 28                 
               .pe14__std__lane28_strm0_ready         ( pe14__std__lane28_strm0_ready      ),      
               .std__pe14__lane28_strm0_cntl          ( std__pe14__lane28_strm0_cntl       ),      
               .std__pe14__lane28_strm0_data          ( std__pe14__lane28_strm0_data       ),      
               .std__pe14__lane28_strm0_data_valid    ( std__pe14__lane28_strm0_data_valid ),      
               .std__pe14__lane28_strm0_data_mask     ( std__pe14__lane28_strm0_data_mask  ),      

               .pe14__std__lane28_strm1_ready         ( pe14__std__lane28_strm1_ready      ),      
               .std__pe14__lane28_strm1_cntl          ( std__pe14__lane28_strm1_cntl       ),      
               .std__pe14__lane28_strm1_data          ( std__pe14__lane28_strm1_data       ),      
               .std__pe14__lane28_strm1_data_valid    ( std__pe14__lane28_strm1_data_valid ),      
               .std__pe14__lane28_strm1_data_mask     ( std__pe14__lane28_strm1_data_mask  ),      

               // PE 14, Lane 29                 
               .pe14__std__lane29_strm0_ready         ( pe14__std__lane29_strm0_ready      ),      
               .std__pe14__lane29_strm0_cntl          ( std__pe14__lane29_strm0_cntl       ),      
               .std__pe14__lane29_strm0_data          ( std__pe14__lane29_strm0_data       ),      
               .std__pe14__lane29_strm0_data_valid    ( std__pe14__lane29_strm0_data_valid ),      
               .std__pe14__lane29_strm0_data_mask     ( std__pe14__lane29_strm0_data_mask  ),      

               .pe14__std__lane29_strm1_ready         ( pe14__std__lane29_strm1_ready      ),      
               .std__pe14__lane29_strm1_cntl          ( std__pe14__lane29_strm1_cntl       ),      
               .std__pe14__lane29_strm1_data          ( std__pe14__lane29_strm1_data       ),      
               .std__pe14__lane29_strm1_data_valid    ( std__pe14__lane29_strm1_data_valid ),      
               .std__pe14__lane29_strm1_data_mask     ( std__pe14__lane29_strm1_data_mask  ),      

               // PE 14, Lane 30                 
               .pe14__std__lane30_strm0_ready         ( pe14__std__lane30_strm0_ready      ),      
               .std__pe14__lane30_strm0_cntl          ( std__pe14__lane30_strm0_cntl       ),      
               .std__pe14__lane30_strm0_data          ( std__pe14__lane30_strm0_data       ),      
               .std__pe14__lane30_strm0_data_valid    ( std__pe14__lane30_strm0_data_valid ),      
               .std__pe14__lane30_strm0_data_mask     ( std__pe14__lane30_strm0_data_mask  ),      

               .pe14__std__lane30_strm1_ready         ( pe14__std__lane30_strm1_ready      ),      
               .std__pe14__lane30_strm1_cntl          ( std__pe14__lane30_strm1_cntl       ),      
               .std__pe14__lane30_strm1_data          ( std__pe14__lane30_strm1_data       ),      
               .std__pe14__lane30_strm1_data_valid    ( std__pe14__lane30_strm1_data_valid ),      
               .std__pe14__lane30_strm1_data_mask     ( std__pe14__lane30_strm1_data_mask  ),      

               // PE 14, Lane 31                 
               .pe14__std__lane31_strm0_ready         ( pe14__std__lane31_strm0_ready      ),      
               .std__pe14__lane31_strm0_cntl          ( std__pe14__lane31_strm0_cntl       ),      
               .std__pe14__lane31_strm0_data          ( std__pe14__lane31_strm0_data       ),      
               .std__pe14__lane31_strm0_data_valid    ( std__pe14__lane31_strm0_data_valid ),      
               .std__pe14__lane31_strm0_data_mask     ( std__pe14__lane31_strm0_data_mask  ),      

               .pe14__std__lane31_strm1_ready         ( pe14__std__lane31_strm1_ready      ),      
               .std__pe14__lane31_strm1_cntl          ( std__pe14__lane31_strm1_cntl       ),      
               .std__pe14__lane31_strm1_data          ( std__pe14__lane31_strm1_data       ),      
               .std__pe14__lane31_strm1_data_valid    ( std__pe14__lane31_strm1_data_valid ),      
               .std__pe14__lane31_strm1_data_mask     ( std__pe14__lane31_strm1_data_mask  ),      

               // PE 15, Lane 0                 
               .pe15__std__lane0_strm0_ready         ( pe15__std__lane0_strm0_ready      ),      
               .std__pe15__lane0_strm0_cntl          ( std__pe15__lane0_strm0_cntl       ),      
               .std__pe15__lane0_strm0_data          ( std__pe15__lane0_strm0_data       ),      
               .std__pe15__lane0_strm0_data_valid    ( std__pe15__lane0_strm0_data_valid ),      
               .std__pe15__lane0_strm0_data_mask     ( std__pe15__lane0_strm0_data_mask  ),      

               .pe15__std__lane0_strm1_ready         ( pe15__std__lane0_strm1_ready      ),      
               .std__pe15__lane0_strm1_cntl          ( std__pe15__lane0_strm1_cntl       ),      
               .std__pe15__lane0_strm1_data          ( std__pe15__lane0_strm1_data       ),      
               .std__pe15__lane0_strm1_data_valid    ( std__pe15__lane0_strm1_data_valid ),      
               .std__pe15__lane0_strm1_data_mask     ( std__pe15__lane0_strm1_data_mask  ),      

               // PE 15, Lane 1                 
               .pe15__std__lane1_strm0_ready         ( pe15__std__lane1_strm0_ready      ),      
               .std__pe15__lane1_strm0_cntl          ( std__pe15__lane1_strm0_cntl       ),      
               .std__pe15__lane1_strm0_data          ( std__pe15__lane1_strm0_data       ),      
               .std__pe15__lane1_strm0_data_valid    ( std__pe15__lane1_strm0_data_valid ),      
               .std__pe15__lane1_strm0_data_mask     ( std__pe15__lane1_strm0_data_mask  ),      

               .pe15__std__lane1_strm1_ready         ( pe15__std__lane1_strm1_ready      ),      
               .std__pe15__lane1_strm1_cntl          ( std__pe15__lane1_strm1_cntl       ),      
               .std__pe15__lane1_strm1_data          ( std__pe15__lane1_strm1_data       ),      
               .std__pe15__lane1_strm1_data_valid    ( std__pe15__lane1_strm1_data_valid ),      
               .std__pe15__lane1_strm1_data_mask     ( std__pe15__lane1_strm1_data_mask  ),      

               // PE 15, Lane 2                 
               .pe15__std__lane2_strm0_ready         ( pe15__std__lane2_strm0_ready      ),      
               .std__pe15__lane2_strm0_cntl          ( std__pe15__lane2_strm0_cntl       ),      
               .std__pe15__lane2_strm0_data          ( std__pe15__lane2_strm0_data       ),      
               .std__pe15__lane2_strm0_data_valid    ( std__pe15__lane2_strm0_data_valid ),      
               .std__pe15__lane2_strm0_data_mask     ( std__pe15__lane2_strm0_data_mask  ),      

               .pe15__std__lane2_strm1_ready         ( pe15__std__lane2_strm1_ready      ),      
               .std__pe15__lane2_strm1_cntl          ( std__pe15__lane2_strm1_cntl       ),      
               .std__pe15__lane2_strm1_data          ( std__pe15__lane2_strm1_data       ),      
               .std__pe15__lane2_strm1_data_valid    ( std__pe15__lane2_strm1_data_valid ),      
               .std__pe15__lane2_strm1_data_mask     ( std__pe15__lane2_strm1_data_mask  ),      

               // PE 15, Lane 3                 
               .pe15__std__lane3_strm0_ready         ( pe15__std__lane3_strm0_ready      ),      
               .std__pe15__lane3_strm0_cntl          ( std__pe15__lane3_strm0_cntl       ),      
               .std__pe15__lane3_strm0_data          ( std__pe15__lane3_strm0_data       ),      
               .std__pe15__lane3_strm0_data_valid    ( std__pe15__lane3_strm0_data_valid ),      
               .std__pe15__lane3_strm0_data_mask     ( std__pe15__lane3_strm0_data_mask  ),      

               .pe15__std__lane3_strm1_ready         ( pe15__std__lane3_strm1_ready      ),      
               .std__pe15__lane3_strm1_cntl          ( std__pe15__lane3_strm1_cntl       ),      
               .std__pe15__lane3_strm1_data          ( std__pe15__lane3_strm1_data       ),      
               .std__pe15__lane3_strm1_data_valid    ( std__pe15__lane3_strm1_data_valid ),      
               .std__pe15__lane3_strm1_data_mask     ( std__pe15__lane3_strm1_data_mask  ),      

               // PE 15, Lane 4                 
               .pe15__std__lane4_strm0_ready         ( pe15__std__lane4_strm0_ready      ),      
               .std__pe15__lane4_strm0_cntl          ( std__pe15__lane4_strm0_cntl       ),      
               .std__pe15__lane4_strm0_data          ( std__pe15__lane4_strm0_data       ),      
               .std__pe15__lane4_strm0_data_valid    ( std__pe15__lane4_strm0_data_valid ),      
               .std__pe15__lane4_strm0_data_mask     ( std__pe15__lane4_strm0_data_mask  ),      

               .pe15__std__lane4_strm1_ready         ( pe15__std__lane4_strm1_ready      ),      
               .std__pe15__lane4_strm1_cntl          ( std__pe15__lane4_strm1_cntl       ),      
               .std__pe15__lane4_strm1_data          ( std__pe15__lane4_strm1_data       ),      
               .std__pe15__lane4_strm1_data_valid    ( std__pe15__lane4_strm1_data_valid ),      
               .std__pe15__lane4_strm1_data_mask     ( std__pe15__lane4_strm1_data_mask  ),      

               // PE 15, Lane 5                 
               .pe15__std__lane5_strm0_ready         ( pe15__std__lane5_strm0_ready      ),      
               .std__pe15__lane5_strm0_cntl          ( std__pe15__lane5_strm0_cntl       ),      
               .std__pe15__lane5_strm0_data          ( std__pe15__lane5_strm0_data       ),      
               .std__pe15__lane5_strm0_data_valid    ( std__pe15__lane5_strm0_data_valid ),      
               .std__pe15__lane5_strm0_data_mask     ( std__pe15__lane5_strm0_data_mask  ),      

               .pe15__std__lane5_strm1_ready         ( pe15__std__lane5_strm1_ready      ),      
               .std__pe15__lane5_strm1_cntl          ( std__pe15__lane5_strm1_cntl       ),      
               .std__pe15__lane5_strm1_data          ( std__pe15__lane5_strm1_data       ),      
               .std__pe15__lane5_strm1_data_valid    ( std__pe15__lane5_strm1_data_valid ),      
               .std__pe15__lane5_strm1_data_mask     ( std__pe15__lane5_strm1_data_mask  ),      

               // PE 15, Lane 6                 
               .pe15__std__lane6_strm0_ready         ( pe15__std__lane6_strm0_ready      ),      
               .std__pe15__lane6_strm0_cntl          ( std__pe15__lane6_strm0_cntl       ),      
               .std__pe15__lane6_strm0_data          ( std__pe15__lane6_strm0_data       ),      
               .std__pe15__lane6_strm0_data_valid    ( std__pe15__lane6_strm0_data_valid ),      
               .std__pe15__lane6_strm0_data_mask     ( std__pe15__lane6_strm0_data_mask  ),      

               .pe15__std__lane6_strm1_ready         ( pe15__std__lane6_strm1_ready      ),      
               .std__pe15__lane6_strm1_cntl          ( std__pe15__lane6_strm1_cntl       ),      
               .std__pe15__lane6_strm1_data          ( std__pe15__lane6_strm1_data       ),      
               .std__pe15__lane6_strm1_data_valid    ( std__pe15__lane6_strm1_data_valid ),      
               .std__pe15__lane6_strm1_data_mask     ( std__pe15__lane6_strm1_data_mask  ),      

               // PE 15, Lane 7                 
               .pe15__std__lane7_strm0_ready         ( pe15__std__lane7_strm0_ready      ),      
               .std__pe15__lane7_strm0_cntl          ( std__pe15__lane7_strm0_cntl       ),      
               .std__pe15__lane7_strm0_data          ( std__pe15__lane7_strm0_data       ),      
               .std__pe15__lane7_strm0_data_valid    ( std__pe15__lane7_strm0_data_valid ),      
               .std__pe15__lane7_strm0_data_mask     ( std__pe15__lane7_strm0_data_mask  ),      

               .pe15__std__lane7_strm1_ready         ( pe15__std__lane7_strm1_ready      ),      
               .std__pe15__lane7_strm1_cntl          ( std__pe15__lane7_strm1_cntl       ),      
               .std__pe15__lane7_strm1_data          ( std__pe15__lane7_strm1_data       ),      
               .std__pe15__lane7_strm1_data_valid    ( std__pe15__lane7_strm1_data_valid ),      
               .std__pe15__lane7_strm1_data_mask     ( std__pe15__lane7_strm1_data_mask  ),      

               // PE 15, Lane 8                 
               .pe15__std__lane8_strm0_ready         ( pe15__std__lane8_strm0_ready      ),      
               .std__pe15__lane8_strm0_cntl          ( std__pe15__lane8_strm0_cntl       ),      
               .std__pe15__lane8_strm0_data          ( std__pe15__lane8_strm0_data       ),      
               .std__pe15__lane8_strm0_data_valid    ( std__pe15__lane8_strm0_data_valid ),      
               .std__pe15__lane8_strm0_data_mask     ( std__pe15__lane8_strm0_data_mask  ),      

               .pe15__std__lane8_strm1_ready         ( pe15__std__lane8_strm1_ready      ),      
               .std__pe15__lane8_strm1_cntl          ( std__pe15__lane8_strm1_cntl       ),      
               .std__pe15__lane8_strm1_data          ( std__pe15__lane8_strm1_data       ),      
               .std__pe15__lane8_strm1_data_valid    ( std__pe15__lane8_strm1_data_valid ),      
               .std__pe15__lane8_strm1_data_mask     ( std__pe15__lane8_strm1_data_mask  ),      

               // PE 15, Lane 9                 
               .pe15__std__lane9_strm0_ready         ( pe15__std__lane9_strm0_ready      ),      
               .std__pe15__lane9_strm0_cntl          ( std__pe15__lane9_strm0_cntl       ),      
               .std__pe15__lane9_strm0_data          ( std__pe15__lane9_strm0_data       ),      
               .std__pe15__lane9_strm0_data_valid    ( std__pe15__lane9_strm0_data_valid ),      
               .std__pe15__lane9_strm0_data_mask     ( std__pe15__lane9_strm0_data_mask  ),      

               .pe15__std__lane9_strm1_ready         ( pe15__std__lane9_strm1_ready      ),      
               .std__pe15__lane9_strm1_cntl          ( std__pe15__lane9_strm1_cntl       ),      
               .std__pe15__lane9_strm1_data          ( std__pe15__lane9_strm1_data       ),      
               .std__pe15__lane9_strm1_data_valid    ( std__pe15__lane9_strm1_data_valid ),      
               .std__pe15__lane9_strm1_data_mask     ( std__pe15__lane9_strm1_data_mask  ),      

               // PE 15, Lane 10                 
               .pe15__std__lane10_strm0_ready         ( pe15__std__lane10_strm0_ready      ),      
               .std__pe15__lane10_strm0_cntl          ( std__pe15__lane10_strm0_cntl       ),      
               .std__pe15__lane10_strm0_data          ( std__pe15__lane10_strm0_data       ),      
               .std__pe15__lane10_strm0_data_valid    ( std__pe15__lane10_strm0_data_valid ),      
               .std__pe15__lane10_strm0_data_mask     ( std__pe15__lane10_strm0_data_mask  ),      

               .pe15__std__lane10_strm1_ready         ( pe15__std__lane10_strm1_ready      ),      
               .std__pe15__lane10_strm1_cntl          ( std__pe15__lane10_strm1_cntl       ),      
               .std__pe15__lane10_strm1_data          ( std__pe15__lane10_strm1_data       ),      
               .std__pe15__lane10_strm1_data_valid    ( std__pe15__lane10_strm1_data_valid ),      
               .std__pe15__lane10_strm1_data_mask     ( std__pe15__lane10_strm1_data_mask  ),      

               // PE 15, Lane 11                 
               .pe15__std__lane11_strm0_ready         ( pe15__std__lane11_strm0_ready      ),      
               .std__pe15__lane11_strm0_cntl          ( std__pe15__lane11_strm0_cntl       ),      
               .std__pe15__lane11_strm0_data          ( std__pe15__lane11_strm0_data       ),      
               .std__pe15__lane11_strm0_data_valid    ( std__pe15__lane11_strm0_data_valid ),      
               .std__pe15__lane11_strm0_data_mask     ( std__pe15__lane11_strm0_data_mask  ),      

               .pe15__std__lane11_strm1_ready         ( pe15__std__lane11_strm1_ready      ),      
               .std__pe15__lane11_strm1_cntl          ( std__pe15__lane11_strm1_cntl       ),      
               .std__pe15__lane11_strm1_data          ( std__pe15__lane11_strm1_data       ),      
               .std__pe15__lane11_strm1_data_valid    ( std__pe15__lane11_strm1_data_valid ),      
               .std__pe15__lane11_strm1_data_mask     ( std__pe15__lane11_strm1_data_mask  ),      

               // PE 15, Lane 12                 
               .pe15__std__lane12_strm0_ready         ( pe15__std__lane12_strm0_ready      ),      
               .std__pe15__lane12_strm0_cntl          ( std__pe15__lane12_strm0_cntl       ),      
               .std__pe15__lane12_strm0_data          ( std__pe15__lane12_strm0_data       ),      
               .std__pe15__lane12_strm0_data_valid    ( std__pe15__lane12_strm0_data_valid ),      
               .std__pe15__lane12_strm0_data_mask     ( std__pe15__lane12_strm0_data_mask  ),      

               .pe15__std__lane12_strm1_ready         ( pe15__std__lane12_strm1_ready      ),      
               .std__pe15__lane12_strm1_cntl          ( std__pe15__lane12_strm1_cntl       ),      
               .std__pe15__lane12_strm1_data          ( std__pe15__lane12_strm1_data       ),      
               .std__pe15__lane12_strm1_data_valid    ( std__pe15__lane12_strm1_data_valid ),      
               .std__pe15__lane12_strm1_data_mask     ( std__pe15__lane12_strm1_data_mask  ),      

               // PE 15, Lane 13                 
               .pe15__std__lane13_strm0_ready         ( pe15__std__lane13_strm0_ready      ),      
               .std__pe15__lane13_strm0_cntl          ( std__pe15__lane13_strm0_cntl       ),      
               .std__pe15__lane13_strm0_data          ( std__pe15__lane13_strm0_data       ),      
               .std__pe15__lane13_strm0_data_valid    ( std__pe15__lane13_strm0_data_valid ),      
               .std__pe15__lane13_strm0_data_mask     ( std__pe15__lane13_strm0_data_mask  ),      

               .pe15__std__lane13_strm1_ready         ( pe15__std__lane13_strm1_ready      ),      
               .std__pe15__lane13_strm1_cntl          ( std__pe15__lane13_strm1_cntl       ),      
               .std__pe15__lane13_strm1_data          ( std__pe15__lane13_strm1_data       ),      
               .std__pe15__lane13_strm1_data_valid    ( std__pe15__lane13_strm1_data_valid ),      
               .std__pe15__lane13_strm1_data_mask     ( std__pe15__lane13_strm1_data_mask  ),      

               // PE 15, Lane 14                 
               .pe15__std__lane14_strm0_ready         ( pe15__std__lane14_strm0_ready      ),      
               .std__pe15__lane14_strm0_cntl          ( std__pe15__lane14_strm0_cntl       ),      
               .std__pe15__lane14_strm0_data          ( std__pe15__lane14_strm0_data       ),      
               .std__pe15__lane14_strm0_data_valid    ( std__pe15__lane14_strm0_data_valid ),      
               .std__pe15__lane14_strm0_data_mask     ( std__pe15__lane14_strm0_data_mask  ),      

               .pe15__std__lane14_strm1_ready         ( pe15__std__lane14_strm1_ready      ),      
               .std__pe15__lane14_strm1_cntl          ( std__pe15__lane14_strm1_cntl       ),      
               .std__pe15__lane14_strm1_data          ( std__pe15__lane14_strm1_data       ),      
               .std__pe15__lane14_strm1_data_valid    ( std__pe15__lane14_strm1_data_valid ),      
               .std__pe15__lane14_strm1_data_mask     ( std__pe15__lane14_strm1_data_mask  ),      

               // PE 15, Lane 15                 
               .pe15__std__lane15_strm0_ready         ( pe15__std__lane15_strm0_ready      ),      
               .std__pe15__lane15_strm0_cntl          ( std__pe15__lane15_strm0_cntl       ),      
               .std__pe15__lane15_strm0_data          ( std__pe15__lane15_strm0_data       ),      
               .std__pe15__lane15_strm0_data_valid    ( std__pe15__lane15_strm0_data_valid ),      
               .std__pe15__lane15_strm0_data_mask     ( std__pe15__lane15_strm0_data_mask  ),      

               .pe15__std__lane15_strm1_ready         ( pe15__std__lane15_strm1_ready      ),      
               .std__pe15__lane15_strm1_cntl          ( std__pe15__lane15_strm1_cntl       ),      
               .std__pe15__lane15_strm1_data          ( std__pe15__lane15_strm1_data       ),      
               .std__pe15__lane15_strm1_data_valid    ( std__pe15__lane15_strm1_data_valid ),      
               .std__pe15__lane15_strm1_data_mask     ( std__pe15__lane15_strm1_data_mask  ),      

               // PE 15, Lane 16                 
               .pe15__std__lane16_strm0_ready         ( pe15__std__lane16_strm0_ready      ),      
               .std__pe15__lane16_strm0_cntl          ( std__pe15__lane16_strm0_cntl       ),      
               .std__pe15__lane16_strm0_data          ( std__pe15__lane16_strm0_data       ),      
               .std__pe15__lane16_strm0_data_valid    ( std__pe15__lane16_strm0_data_valid ),      
               .std__pe15__lane16_strm0_data_mask     ( std__pe15__lane16_strm0_data_mask  ),      

               .pe15__std__lane16_strm1_ready         ( pe15__std__lane16_strm1_ready      ),      
               .std__pe15__lane16_strm1_cntl          ( std__pe15__lane16_strm1_cntl       ),      
               .std__pe15__lane16_strm1_data          ( std__pe15__lane16_strm1_data       ),      
               .std__pe15__lane16_strm1_data_valid    ( std__pe15__lane16_strm1_data_valid ),      
               .std__pe15__lane16_strm1_data_mask     ( std__pe15__lane16_strm1_data_mask  ),      

               // PE 15, Lane 17                 
               .pe15__std__lane17_strm0_ready         ( pe15__std__lane17_strm0_ready      ),      
               .std__pe15__lane17_strm0_cntl          ( std__pe15__lane17_strm0_cntl       ),      
               .std__pe15__lane17_strm0_data          ( std__pe15__lane17_strm0_data       ),      
               .std__pe15__lane17_strm0_data_valid    ( std__pe15__lane17_strm0_data_valid ),      
               .std__pe15__lane17_strm0_data_mask     ( std__pe15__lane17_strm0_data_mask  ),      

               .pe15__std__lane17_strm1_ready         ( pe15__std__lane17_strm1_ready      ),      
               .std__pe15__lane17_strm1_cntl          ( std__pe15__lane17_strm1_cntl       ),      
               .std__pe15__lane17_strm1_data          ( std__pe15__lane17_strm1_data       ),      
               .std__pe15__lane17_strm1_data_valid    ( std__pe15__lane17_strm1_data_valid ),      
               .std__pe15__lane17_strm1_data_mask     ( std__pe15__lane17_strm1_data_mask  ),      

               // PE 15, Lane 18                 
               .pe15__std__lane18_strm0_ready         ( pe15__std__lane18_strm0_ready      ),      
               .std__pe15__lane18_strm0_cntl          ( std__pe15__lane18_strm0_cntl       ),      
               .std__pe15__lane18_strm0_data          ( std__pe15__lane18_strm0_data       ),      
               .std__pe15__lane18_strm0_data_valid    ( std__pe15__lane18_strm0_data_valid ),      
               .std__pe15__lane18_strm0_data_mask     ( std__pe15__lane18_strm0_data_mask  ),      

               .pe15__std__lane18_strm1_ready         ( pe15__std__lane18_strm1_ready      ),      
               .std__pe15__lane18_strm1_cntl          ( std__pe15__lane18_strm1_cntl       ),      
               .std__pe15__lane18_strm1_data          ( std__pe15__lane18_strm1_data       ),      
               .std__pe15__lane18_strm1_data_valid    ( std__pe15__lane18_strm1_data_valid ),      
               .std__pe15__lane18_strm1_data_mask     ( std__pe15__lane18_strm1_data_mask  ),      

               // PE 15, Lane 19                 
               .pe15__std__lane19_strm0_ready         ( pe15__std__lane19_strm0_ready      ),      
               .std__pe15__lane19_strm0_cntl          ( std__pe15__lane19_strm0_cntl       ),      
               .std__pe15__lane19_strm0_data          ( std__pe15__lane19_strm0_data       ),      
               .std__pe15__lane19_strm0_data_valid    ( std__pe15__lane19_strm0_data_valid ),      
               .std__pe15__lane19_strm0_data_mask     ( std__pe15__lane19_strm0_data_mask  ),      

               .pe15__std__lane19_strm1_ready         ( pe15__std__lane19_strm1_ready      ),      
               .std__pe15__lane19_strm1_cntl          ( std__pe15__lane19_strm1_cntl       ),      
               .std__pe15__lane19_strm1_data          ( std__pe15__lane19_strm1_data       ),      
               .std__pe15__lane19_strm1_data_valid    ( std__pe15__lane19_strm1_data_valid ),      
               .std__pe15__lane19_strm1_data_mask     ( std__pe15__lane19_strm1_data_mask  ),      

               // PE 15, Lane 20                 
               .pe15__std__lane20_strm0_ready         ( pe15__std__lane20_strm0_ready      ),      
               .std__pe15__lane20_strm0_cntl          ( std__pe15__lane20_strm0_cntl       ),      
               .std__pe15__lane20_strm0_data          ( std__pe15__lane20_strm0_data       ),      
               .std__pe15__lane20_strm0_data_valid    ( std__pe15__lane20_strm0_data_valid ),      
               .std__pe15__lane20_strm0_data_mask     ( std__pe15__lane20_strm0_data_mask  ),      

               .pe15__std__lane20_strm1_ready         ( pe15__std__lane20_strm1_ready      ),      
               .std__pe15__lane20_strm1_cntl          ( std__pe15__lane20_strm1_cntl       ),      
               .std__pe15__lane20_strm1_data          ( std__pe15__lane20_strm1_data       ),      
               .std__pe15__lane20_strm1_data_valid    ( std__pe15__lane20_strm1_data_valid ),      
               .std__pe15__lane20_strm1_data_mask     ( std__pe15__lane20_strm1_data_mask  ),      

               // PE 15, Lane 21                 
               .pe15__std__lane21_strm0_ready         ( pe15__std__lane21_strm0_ready      ),      
               .std__pe15__lane21_strm0_cntl          ( std__pe15__lane21_strm0_cntl       ),      
               .std__pe15__lane21_strm0_data          ( std__pe15__lane21_strm0_data       ),      
               .std__pe15__lane21_strm0_data_valid    ( std__pe15__lane21_strm0_data_valid ),      
               .std__pe15__lane21_strm0_data_mask     ( std__pe15__lane21_strm0_data_mask  ),      

               .pe15__std__lane21_strm1_ready         ( pe15__std__lane21_strm1_ready      ),      
               .std__pe15__lane21_strm1_cntl          ( std__pe15__lane21_strm1_cntl       ),      
               .std__pe15__lane21_strm1_data          ( std__pe15__lane21_strm1_data       ),      
               .std__pe15__lane21_strm1_data_valid    ( std__pe15__lane21_strm1_data_valid ),      
               .std__pe15__lane21_strm1_data_mask     ( std__pe15__lane21_strm1_data_mask  ),      

               // PE 15, Lane 22                 
               .pe15__std__lane22_strm0_ready         ( pe15__std__lane22_strm0_ready      ),      
               .std__pe15__lane22_strm0_cntl          ( std__pe15__lane22_strm0_cntl       ),      
               .std__pe15__lane22_strm0_data          ( std__pe15__lane22_strm0_data       ),      
               .std__pe15__lane22_strm0_data_valid    ( std__pe15__lane22_strm0_data_valid ),      
               .std__pe15__lane22_strm0_data_mask     ( std__pe15__lane22_strm0_data_mask  ),      

               .pe15__std__lane22_strm1_ready         ( pe15__std__lane22_strm1_ready      ),      
               .std__pe15__lane22_strm1_cntl          ( std__pe15__lane22_strm1_cntl       ),      
               .std__pe15__lane22_strm1_data          ( std__pe15__lane22_strm1_data       ),      
               .std__pe15__lane22_strm1_data_valid    ( std__pe15__lane22_strm1_data_valid ),      
               .std__pe15__lane22_strm1_data_mask     ( std__pe15__lane22_strm1_data_mask  ),      

               // PE 15, Lane 23                 
               .pe15__std__lane23_strm0_ready         ( pe15__std__lane23_strm0_ready      ),      
               .std__pe15__lane23_strm0_cntl          ( std__pe15__lane23_strm0_cntl       ),      
               .std__pe15__lane23_strm0_data          ( std__pe15__lane23_strm0_data       ),      
               .std__pe15__lane23_strm0_data_valid    ( std__pe15__lane23_strm0_data_valid ),      
               .std__pe15__lane23_strm0_data_mask     ( std__pe15__lane23_strm0_data_mask  ),      

               .pe15__std__lane23_strm1_ready         ( pe15__std__lane23_strm1_ready      ),      
               .std__pe15__lane23_strm1_cntl          ( std__pe15__lane23_strm1_cntl       ),      
               .std__pe15__lane23_strm1_data          ( std__pe15__lane23_strm1_data       ),      
               .std__pe15__lane23_strm1_data_valid    ( std__pe15__lane23_strm1_data_valid ),      
               .std__pe15__lane23_strm1_data_mask     ( std__pe15__lane23_strm1_data_mask  ),      

               // PE 15, Lane 24                 
               .pe15__std__lane24_strm0_ready         ( pe15__std__lane24_strm0_ready      ),      
               .std__pe15__lane24_strm0_cntl          ( std__pe15__lane24_strm0_cntl       ),      
               .std__pe15__lane24_strm0_data          ( std__pe15__lane24_strm0_data       ),      
               .std__pe15__lane24_strm0_data_valid    ( std__pe15__lane24_strm0_data_valid ),      
               .std__pe15__lane24_strm0_data_mask     ( std__pe15__lane24_strm0_data_mask  ),      

               .pe15__std__lane24_strm1_ready         ( pe15__std__lane24_strm1_ready      ),      
               .std__pe15__lane24_strm1_cntl          ( std__pe15__lane24_strm1_cntl       ),      
               .std__pe15__lane24_strm1_data          ( std__pe15__lane24_strm1_data       ),      
               .std__pe15__lane24_strm1_data_valid    ( std__pe15__lane24_strm1_data_valid ),      
               .std__pe15__lane24_strm1_data_mask     ( std__pe15__lane24_strm1_data_mask  ),      

               // PE 15, Lane 25                 
               .pe15__std__lane25_strm0_ready         ( pe15__std__lane25_strm0_ready      ),      
               .std__pe15__lane25_strm0_cntl          ( std__pe15__lane25_strm0_cntl       ),      
               .std__pe15__lane25_strm0_data          ( std__pe15__lane25_strm0_data       ),      
               .std__pe15__lane25_strm0_data_valid    ( std__pe15__lane25_strm0_data_valid ),      
               .std__pe15__lane25_strm0_data_mask     ( std__pe15__lane25_strm0_data_mask  ),      

               .pe15__std__lane25_strm1_ready         ( pe15__std__lane25_strm1_ready      ),      
               .std__pe15__lane25_strm1_cntl          ( std__pe15__lane25_strm1_cntl       ),      
               .std__pe15__lane25_strm1_data          ( std__pe15__lane25_strm1_data       ),      
               .std__pe15__lane25_strm1_data_valid    ( std__pe15__lane25_strm1_data_valid ),      
               .std__pe15__lane25_strm1_data_mask     ( std__pe15__lane25_strm1_data_mask  ),      

               // PE 15, Lane 26                 
               .pe15__std__lane26_strm0_ready         ( pe15__std__lane26_strm0_ready      ),      
               .std__pe15__lane26_strm0_cntl          ( std__pe15__lane26_strm0_cntl       ),      
               .std__pe15__lane26_strm0_data          ( std__pe15__lane26_strm0_data       ),      
               .std__pe15__lane26_strm0_data_valid    ( std__pe15__lane26_strm0_data_valid ),      
               .std__pe15__lane26_strm0_data_mask     ( std__pe15__lane26_strm0_data_mask  ),      

               .pe15__std__lane26_strm1_ready         ( pe15__std__lane26_strm1_ready      ),      
               .std__pe15__lane26_strm1_cntl          ( std__pe15__lane26_strm1_cntl       ),      
               .std__pe15__lane26_strm1_data          ( std__pe15__lane26_strm1_data       ),      
               .std__pe15__lane26_strm1_data_valid    ( std__pe15__lane26_strm1_data_valid ),      
               .std__pe15__lane26_strm1_data_mask     ( std__pe15__lane26_strm1_data_mask  ),      

               // PE 15, Lane 27                 
               .pe15__std__lane27_strm0_ready         ( pe15__std__lane27_strm0_ready      ),      
               .std__pe15__lane27_strm0_cntl          ( std__pe15__lane27_strm0_cntl       ),      
               .std__pe15__lane27_strm0_data          ( std__pe15__lane27_strm0_data       ),      
               .std__pe15__lane27_strm0_data_valid    ( std__pe15__lane27_strm0_data_valid ),      
               .std__pe15__lane27_strm0_data_mask     ( std__pe15__lane27_strm0_data_mask  ),      

               .pe15__std__lane27_strm1_ready         ( pe15__std__lane27_strm1_ready      ),      
               .std__pe15__lane27_strm1_cntl          ( std__pe15__lane27_strm1_cntl       ),      
               .std__pe15__lane27_strm1_data          ( std__pe15__lane27_strm1_data       ),      
               .std__pe15__lane27_strm1_data_valid    ( std__pe15__lane27_strm1_data_valid ),      
               .std__pe15__lane27_strm1_data_mask     ( std__pe15__lane27_strm1_data_mask  ),      

               // PE 15, Lane 28                 
               .pe15__std__lane28_strm0_ready         ( pe15__std__lane28_strm0_ready      ),      
               .std__pe15__lane28_strm0_cntl          ( std__pe15__lane28_strm0_cntl       ),      
               .std__pe15__lane28_strm0_data          ( std__pe15__lane28_strm0_data       ),      
               .std__pe15__lane28_strm0_data_valid    ( std__pe15__lane28_strm0_data_valid ),      
               .std__pe15__lane28_strm0_data_mask     ( std__pe15__lane28_strm0_data_mask  ),      

               .pe15__std__lane28_strm1_ready         ( pe15__std__lane28_strm1_ready      ),      
               .std__pe15__lane28_strm1_cntl          ( std__pe15__lane28_strm1_cntl       ),      
               .std__pe15__lane28_strm1_data          ( std__pe15__lane28_strm1_data       ),      
               .std__pe15__lane28_strm1_data_valid    ( std__pe15__lane28_strm1_data_valid ),      
               .std__pe15__lane28_strm1_data_mask     ( std__pe15__lane28_strm1_data_mask  ),      

               // PE 15, Lane 29                 
               .pe15__std__lane29_strm0_ready         ( pe15__std__lane29_strm0_ready      ),      
               .std__pe15__lane29_strm0_cntl          ( std__pe15__lane29_strm0_cntl       ),      
               .std__pe15__lane29_strm0_data          ( std__pe15__lane29_strm0_data       ),      
               .std__pe15__lane29_strm0_data_valid    ( std__pe15__lane29_strm0_data_valid ),      
               .std__pe15__lane29_strm0_data_mask     ( std__pe15__lane29_strm0_data_mask  ),      

               .pe15__std__lane29_strm1_ready         ( pe15__std__lane29_strm1_ready      ),      
               .std__pe15__lane29_strm1_cntl          ( std__pe15__lane29_strm1_cntl       ),      
               .std__pe15__lane29_strm1_data          ( std__pe15__lane29_strm1_data       ),      
               .std__pe15__lane29_strm1_data_valid    ( std__pe15__lane29_strm1_data_valid ),      
               .std__pe15__lane29_strm1_data_mask     ( std__pe15__lane29_strm1_data_mask  ),      

               // PE 15, Lane 30                 
               .pe15__std__lane30_strm0_ready         ( pe15__std__lane30_strm0_ready      ),      
               .std__pe15__lane30_strm0_cntl          ( std__pe15__lane30_strm0_cntl       ),      
               .std__pe15__lane30_strm0_data          ( std__pe15__lane30_strm0_data       ),      
               .std__pe15__lane30_strm0_data_valid    ( std__pe15__lane30_strm0_data_valid ),      
               .std__pe15__lane30_strm0_data_mask     ( std__pe15__lane30_strm0_data_mask  ),      

               .pe15__std__lane30_strm1_ready         ( pe15__std__lane30_strm1_ready      ),      
               .std__pe15__lane30_strm1_cntl          ( std__pe15__lane30_strm1_cntl       ),      
               .std__pe15__lane30_strm1_data          ( std__pe15__lane30_strm1_data       ),      
               .std__pe15__lane30_strm1_data_valid    ( std__pe15__lane30_strm1_data_valid ),      
               .std__pe15__lane30_strm1_data_mask     ( std__pe15__lane30_strm1_data_mask  ),      

               // PE 15, Lane 31                 
               .pe15__std__lane31_strm0_ready         ( pe15__std__lane31_strm0_ready      ),      
               .std__pe15__lane31_strm0_cntl          ( std__pe15__lane31_strm0_cntl       ),      
               .std__pe15__lane31_strm0_data          ( std__pe15__lane31_strm0_data       ),      
               .std__pe15__lane31_strm0_data_valid    ( std__pe15__lane31_strm0_data_valid ),      
               .std__pe15__lane31_strm0_data_mask     ( std__pe15__lane31_strm0_data_mask  ),      

               .pe15__std__lane31_strm1_ready         ( pe15__std__lane31_strm1_ready      ),      
               .std__pe15__lane31_strm1_cntl          ( std__pe15__lane31_strm1_cntl       ),      
               .std__pe15__lane31_strm1_data          ( std__pe15__lane31_strm1_data       ),      
               .std__pe15__lane31_strm1_data_valid    ( std__pe15__lane31_strm1_data_valid ),      
               .std__pe15__lane31_strm1_data_mask     ( std__pe15__lane31_strm1_data_mask  ),      

               // PE 16, Lane 0                 
               .pe16__std__lane0_strm0_ready         ( pe16__std__lane0_strm0_ready      ),      
               .std__pe16__lane0_strm0_cntl          ( std__pe16__lane0_strm0_cntl       ),      
               .std__pe16__lane0_strm0_data          ( std__pe16__lane0_strm0_data       ),      
               .std__pe16__lane0_strm0_data_valid    ( std__pe16__lane0_strm0_data_valid ),      
               .std__pe16__lane0_strm0_data_mask     ( std__pe16__lane0_strm0_data_mask  ),      

               .pe16__std__lane0_strm1_ready         ( pe16__std__lane0_strm1_ready      ),      
               .std__pe16__lane0_strm1_cntl          ( std__pe16__lane0_strm1_cntl       ),      
               .std__pe16__lane0_strm1_data          ( std__pe16__lane0_strm1_data       ),      
               .std__pe16__lane0_strm1_data_valid    ( std__pe16__lane0_strm1_data_valid ),      
               .std__pe16__lane0_strm1_data_mask     ( std__pe16__lane0_strm1_data_mask  ),      

               // PE 16, Lane 1                 
               .pe16__std__lane1_strm0_ready         ( pe16__std__lane1_strm0_ready      ),      
               .std__pe16__lane1_strm0_cntl          ( std__pe16__lane1_strm0_cntl       ),      
               .std__pe16__lane1_strm0_data          ( std__pe16__lane1_strm0_data       ),      
               .std__pe16__lane1_strm0_data_valid    ( std__pe16__lane1_strm0_data_valid ),      
               .std__pe16__lane1_strm0_data_mask     ( std__pe16__lane1_strm0_data_mask  ),      

               .pe16__std__lane1_strm1_ready         ( pe16__std__lane1_strm1_ready      ),      
               .std__pe16__lane1_strm1_cntl          ( std__pe16__lane1_strm1_cntl       ),      
               .std__pe16__lane1_strm1_data          ( std__pe16__lane1_strm1_data       ),      
               .std__pe16__lane1_strm1_data_valid    ( std__pe16__lane1_strm1_data_valid ),      
               .std__pe16__lane1_strm1_data_mask     ( std__pe16__lane1_strm1_data_mask  ),      

               // PE 16, Lane 2                 
               .pe16__std__lane2_strm0_ready         ( pe16__std__lane2_strm0_ready      ),      
               .std__pe16__lane2_strm0_cntl          ( std__pe16__lane2_strm0_cntl       ),      
               .std__pe16__lane2_strm0_data          ( std__pe16__lane2_strm0_data       ),      
               .std__pe16__lane2_strm0_data_valid    ( std__pe16__lane2_strm0_data_valid ),      
               .std__pe16__lane2_strm0_data_mask     ( std__pe16__lane2_strm0_data_mask  ),      

               .pe16__std__lane2_strm1_ready         ( pe16__std__lane2_strm1_ready      ),      
               .std__pe16__lane2_strm1_cntl          ( std__pe16__lane2_strm1_cntl       ),      
               .std__pe16__lane2_strm1_data          ( std__pe16__lane2_strm1_data       ),      
               .std__pe16__lane2_strm1_data_valid    ( std__pe16__lane2_strm1_data_valid ),      
               .std__pe16__lane2_strm1_data_mask     ( std__pe16__lane2_strm1_data_mask  ),      

               // PE 16, Lane 3                 
               .pe16__std__lane3_strm0_ready         ( pe16__std__lane3_strm0_ready      ),      
               .std__pe16__lane3_strm0_cntl          ( std__pe16__lane3_strm0_cntl       ),      
               .std__pe16__lane3_strm0_data          ( std__pe16__lane3_strm0_data       ),      
               .std__pe16__lane3_strm0_data_valid    ( std__pe16__lane3_strm0_data_valid ),      
               .std__pe16__lane3_strm0_data_mask     ( std__pe16__lane3_strm0_data_mask  ),      

               .pe16__std__lane3_strm1_ready         ( pe16__std__lane3_strm1_ready      ),      
               .std__pe16__lane3_strm1_cntl          ( std__pe16__lane3_strm1_cntl       ),      
               .std__pe16__lane3_strm1_data          ( std__pe16__lane3_strm1_data       ),      
               .std__pe16__lane3_strm1_data_valid    ( std__pe16__lane3_strm1_data_valid ),      
               .std__pe16__lane3_strm1_data_mask     ( std__pe16__lane3_strm1_data_mask  ),      

               // PE 16, Lane 4                 
               .pe16__std__lane4_strm0_ready         ( pe16__std__lane4_strm0_ready      ),      
               .std__pe16__lane4_strm0_cntl          ( std__pe16__lane4_strm0_cntl       ),      
               .std__pe16__lane4_strm0_data          ( std__pe16__lane4_strm0_data       ),      
               .std__pe16__lane4_strm0_data_valid    ( std__pe16__lane4_strm0_data_valid ),      
               .std__pe16__lane4_strm0_data_mask     ( std__pe16__lane4_strm0_data_mask  ),      

               .pe16__std__lane4_strm1_ready         ( pe16__std__lane4_strm1_ready      ),      
               .std__pe16__lane4_strm1_cntl          ( std__pe16__lane4_strm1_cntl       ),      
               .std__pe16__lane4_strm1_data          ( std__pe16__lane4_strm1_data       ),      
               .std__pe16__lane4_strm1_data_valid    ( std__pe16__lane4_strm1_data_valid ),      
               .std__pe16__lane4_strm1_data_mask     ( std__pe16__lane4_strm1_data_mask  ),      

               // PE 16, Lane 5                 
               .pe16__std__lane5_strm0_ready         ( pe16__std__lane5_strm0_ready      ),      
               .std__pe16__lane5_strm0_cntl          ( std__pe16__lane5_strm0_cntl       ),      
               .std__pe16__lane5_strm0_data          ( std__pe16__lane5_strm0_data       ),      
               .std__pe16__lane5_strm0_data_valid    ( std__pe16__lane5_strm0_data_valid ),      
               .std__pe16__lane5_strm0_data_mask     ( std__pe16__lane5_strm0_data_mask  ),      

               .pe16__std__lane5_strm1_ready         ( pe16__std__lane5_strm1_ready      ),      
               .std__pe16__lane5_strm1_cntl          ( std__pe16__lane5_strm1_cntl       ),      
               .std__pe16__lane5_strm1_data          ( std__pe16__lane5_strm1_data       ),      
               .std__pe16__lane5_strm1_data_valid    ( std__pe16__lane5_strm1_data_valid ),      
               .std__pe16__lane5_strm1_data_mask     ( std__pe16__lane5_strm1_data_mask  ),      

               // PE 16, Lane 6                 
               .pe16__std__lane6_strm0_ready         ( pe16__std__lane6_strm0_ready      ),      
               .std__pe16__lane6_strm0_cntl          ( std__pe16__lane6_strm0_cntl       ),      
               .std__pe16__lane6_strm0_data          ( std__pe16__lane6_strm0_data       ),      
               .std__pe16__lane6_strm0_data_valid    ( std__pe16__lane6_strm0_data_valid ),      
               .std__pe16__lane6_strm0_data_mask     ( std__pe16__lane6_strm0_data_mask  ),      

               .pe16__std__lane6_strm1_ready         ( pe16__std__lane6_strm1_ready      ),      
               .std__pe16__lane6_strm1_cntl          ( std__pe16__lane6_strm1_cntl       ),      
               .std__pe16__lane6_strm1_data          ( std__pe16__lane6_strm1_data       ),      
               .std__pe16__lane6_strm1_data_valid    ( std__pe16__lane6_strm1_data_valid ),      
               .std__pe16__lane6_strm1_data_mask     ( std__pe16__lane6_strm1_data_mask  ),      

               // PE 16, Lane 7                 
               .pe16__std__lane7_strm0_ready         ( pe16__std__lane7_strm0_ready      ),      
               .std__pe16__lane7_strm0_cntl          ( std__pe16__lane7_strm0_cntl       ),      
               .std__pe16__lane7_strm0_data          ( std__pe16__lane7_strm0_data       ),      
               .std__pe16__lane7_strm0_data_valid    ( std__pe16__lane7_strm0_data_valid ),      
               .std__pe16__lane7_strm0_data_mask     ( std__pe16__lane7_strm0_data_mask  ),      

               .pe16__std__lane7_strm1_ready         ( pe16__std__lane7_strm1_ready      ),      
               .std__pe16__lane7_strm1_cntl          ( std__pe16__lane7_strm1_cntl       ),      
               .std__pe16__lane7_strm1_data          ( std__pe16__lane7_strm1_data       ),      
               .std__pe16__lane7_strm1_data_valid    ( std__pe16__lane7_strm1_data_valid ),      
               .std__pe16__lane7_strm1_data_mask     ( std__pe16__lane7_strm1_data_mask  ),      

               // PE 16, Lane 8                 
               .pe16__std__lane8_strm0_ready         ( pe16__std__lane8_strm0_ready      ),      
               .std__pe16__lane8_strm0_cntl          ( std__pe16__lane8_strm0_cntl       ),      
               .std__pe16__lane8_strm0_data          ( std__pe16__lane8_strm0_data       ),      
               .std__pe16__lane8_strm0_data_valid    ( std__pe16__lane8_strm0_data_valid ),      
               .std__pe16__lane8_strm0_data_mask     ( std__pe16__lane8_strm0_data_mask  ),      

               .pe16__std__lane8_strm1_ready         ( pe16__std__lane8_strm1_ready      ),      
               .std__pe16__lane8_strm1_cntl          ( std__pe16__lane8_strm1_cntl       ),      
               .std__pe16__lane8_strm1_data          ( std__pe16__lane8_strm1_data       ),      
               .std__pe16__lane8_strm1_data_valid    ( std__pe16__lane8_strm1_data_valid ),      
               .std__pe16__lane8_strm1_data_mask     ( std__pe16__lane8_strm1_data_mask  ),      

               // PE 16, Lane 9                 
               .pe16__std__lane9_strm0_ready         ( pe16__std__lane9_strm0_ready      ),      
               .std__pe16__lane9_strm0_cntl          ( std__pe16__lane9_strm0_cntl       ),      
               .std__pe16__lane9_strm0_data          ( std__pe16__lane9_strm0_data       ),      
               .std__pe16__lane9_strm0_data_valid    ( std__pe16__lane9_strm0_data_valid ),      
               .std__pe16__lane9_strm0_data_mask     ( std__pe16__lane9_strm0_data_mask  ),      

               .pe16__std__lane9_strm1_ready         ( pe16__std__lane9_strm1_ready      ),      
               .std__pe16__lane9_strm1_cntl          ( std__pe16__lane9_strm1_cntl       ),      
               .std__pe16__lane9_strm1_data          ( std__pe16__lane9_strm1_data       ),      
               .std__pe16__lane9_strm1_data_valid    ( std__pe16__lane9_strm1_data_valid ),      
               .std__pe16__lane9_strm1_data_mask     ( std__pe16__lane9_strm1_data_mask  ),      

               // PE 16, Lane 10                 
               .pe16__std__lane10_strm0_ready         ( pe16__std__lane10_strm0_ready      ),      
               .std__pe16__lane10_strm0_cntl          ( std__pe16__lane10_strm0_cntl       ),      
               .std__pe16__lane10_strm0_data          ( std__pe16__lane10_strm0_data       ),      
               .std__pe16__lane10_strm0_data_valid    ( std__pe16__lane10_strm0_data_valid ),      
               .std__pe16__lane10_strm0_data_mask     ( std__pe16__lane10_strm0_data_mask  ),      

               .pe16__std__lane10_strm1_ready         ( pe16__std__lane10_strm1_ready      ),      
               .std__pe16__lane10_strm1_cntl          ( std__pe16__lane10_strm1_cntl       ),      
               .std__pe16__lane10_strm1_data          ( std__pe16__lane10_strm1_data       ),      
               .std__pe16__lane10_strm1_data_valid    ( std__pe16__lane10_strm1_data_valid ),      
               .std__pe16__lane10_strm1_data_mask     ( std__pe16__lane10_strm1_data_mask  ),      

               // PE 16, Lane 11                 
               .pe16__std__lane11_strm0_ready         ( pe16__std__lane11_strm0_ready      ),      
               .std__pe16__lane11_strm0_cntl          ( std__pe16__lane11_strm0_cntl       ),      
               .std__pe16__lane11_strm0_data          ( std__pe16__lane11_strm0_data       ),      
               .std__pe16__lane11_strm0_data_valid    ( std__pe16__lane11_strm0_data_valid ),      
               .std__pe16__lane11_strm0_data_mask     ( std__pe16__lane11_strm0_data_mask  ),      

               .pe16__std__lane11_strm1_ready         ( pe16__std__lane11_strm1_ready      ),      
               .std__pe16__lane11_strm1_cntl          ( std__pe16__lane11_strm1_cntl       ),      
               .std__pe16__lane11_strm1_data          ( std__pe16__lane11_strm1_data       ),      
               .std__pe16__lane11_strm1_data_valid    ( std__pe16__lane11_strm1_data_valid ),      
               .std__pe16__lane11_strm1_data_mask     ( std__pe16__lane11_strm1_data_mask  ),      

               // PE 16, Lane 12                 
               .pe16__std__lane12_strm0_ready         ( pe16__std__lane12_strm0_ready      ),      
               .std__pe16__lane12_strm0_cntl          ( std__pe16__lane12_strm0_cntl       ),      
               .std__pe16__lane12_strm0_data          ( std__pe16__lane12_strm0_data       ),      
               .std__pe16__lane12_strm0_data_valid    ( std__pe16__lane12_strm0_data_valid ),      
               .std__pe16__lane12_strm0_data_mask     ( std__pe16__lane12_strm0_data_mask  ),      

               .pe16__std__lane12_strm1_ready         ( pe16__std__lane12_strm1_ready      ),      
               .std__pe16__lane12_strm1_cntl          ( std__pe16__lane12_strm1_cntl       ),      
               .std__pe16__lane12_strm1_data          ( std__pe16__lane12_strm1_data       ),      
               .std__pe16__lane12_strm1_data_valid    ( std__pe16__lane12_strm1_data_valid ),      
               .std__pe16__lane12_strm1_data_mask     ( std__pe16__lane12_strm1_data_mask  ),      

               // PE 16, Lane 13                 
               .pe16__std__lane13_strm0_ready         ( pe16__std__lane13_strm0_ready      ),      
               .std__pe16__lane13_strm0_cntl          ( std__pe16__lane13_strm0_cntl       ),      
               .std__pe16__lane13_strm0_data          ( std__pe16__lane13_strm0_data       ),      
               .std__pe16__lane13_strm0_data_valid    ( std__pe16__lane13_strm0_data_valid ),      
               .std__pe16__lane13_strm0_data_mask     ( std__pe16__lane13_strm0_data_mask  ),      

               .pe16__std__lane13_strm1_ready         ( pe16__std__lane13_strm1_ready      ),      
               .std__pe16__lane13_strm1_cntl          ( std__pe16__lane13_strm1_cntl       ),      
               .std__pe16__lane13_strm1_data          ( std__pe16__lane13_strm1_data       ),      
               .std__pe16__lane13_strm1_data_valid    ( std__pe16__lane13_strm1_data_valid ),      
               .std__pe16__lane13_strm1_data_mask     ( std__pe16__lane13_strm1_data_mask  ),      

               // PE 16, Lane 14                 
               .pe16__std__lane14_strm0_ready         ( pe16__std__lane14_strm0_ready      ),      
               .std__pe16__lane14_strm0_cntl          ( std__pe16__lane14_strm0_cntl       ),      
               .std__pe16__lane14_strm0_data          ( std__pe16__lane14_strm0_data       ),      
               .std__pe16__lane14_strm0_data_valid    ( std__pe16__lane14_strm0_data_valid ),      
               .std__pe16__lane14_strm0_data_mask     ( std__pe16__lane14_strm0_data_mask  ),      

               .pe16__std__lane14_strm1_ready         ( pe16__std__lane14_strm1_ready      ),      
               .std__pe16__lane14_strm1_cntl          ( std__pe16__lane14_strm1_cntl       ),      
               .std__pe16__lane14_strm1_data          ( std__pe16__lane14_strm1_data       ),      
               .std__pe16__lane14_strm1_data_valid    ( std__pe16__lane14_strm1_data_valid ),      
               .std__pe16__lane14_strm1_data_mask     ( std__pe16__lane14_strm1_data_mask  ),      

               // PE 16, Lane 15                 
               .pe16__std__lane15_strm0_ready         ( pe16__std__lane15_strm0_ready      ),      
               .std__pe16__lane15_strm0_cntl          ( std__pe16__lane15_strm0_cntl       ),      
               .std__pe16__lane15_strm0_data          ( std__pe16__lane15_strm0_data       ),      
               .std__pe16__lane15_strm0_data_valid    ( std__pe16__lane15_strm0_data_valid ),      
               .std__pe16__lane15_strm0_data_mask     ( std__pe16__lane15_strm0_data_mask  ),      

               .pe16__std__lane15_strm1_ready         ( pe16__std__lane15_strm1_ready      ),      
               .std__pe16__lane15_strm1_cntl          ( std__pe16__lane15_strm1_cntl       ),      
               .std__pe16__lane15_strm1_data          ( std__pe16__lane15_strm1_data       ),      
               .std__pe16__lane15_strm1_data_valid    ( std__pe16__lane15_strm1_data_valid ),      
               .std__pe16__lane15_strm1_data_mask     ( std__pe16__lane15_strm1_data_mask  ),      

               // PE 16, Lane 16                 
               .pe16__std__lane16_strm0_ready         ( pe16__std__lane16_strm0_ready      ),      
               .std__pe16__lane16_strm0_cntl          ( std__pe16__lane16_strm0_cntl       ),      
               .std__pe16__lane16_strm0_data          ( std__pe16__lane16_strm0_data       ),      
               .std__pe16__lane16_strm0_data_valid    ( std__pe16__lane16_strm0_data_valid ),      
               .std__pe16__lane16_strm0_data_mask     ( std__pe16__lane16_strm0_data_mask  ),      

               .pe16__std__lane16_strm1_ready         ( pe16__std__lane16_strm1_ready      ),      
               .std__pe16__lane16_strm1_cntl          ( std__pe16__lane16_strm1_cntl       ),      
               .std__pe16__lane16_strm1_data          ( std__pe16__lane16_strm1_data       ),      
               .std__pe16__lane16_strm1_data_valid    ( std__pe16__lane16_strm1_data_valid ),      
               .std__pe16__lane16_strm1_data_mask     ( std__pe16__lane16_strm1_data_mask  ),      

               // PE 16, Lane 17                 
               .pe16__std__lane17_strm0_ready         ( pe16__std__lane17_strm0_ready      ),      
               .std__pe16__lane17_strm0_cntl          ( std__pe16__lane17_strm0_cntl       ),      
               .std__pe16__lane17_strm0_data          ( std__pe16__lane17_strm0_data       ),      
               .std__pe16__lane17_strm0_data_valid    ( std__pe16__lane17_strm0_data_valid ),      
               .std__pe16__lane17_strm0_data_mask     ( std__pe16__lane17_strm0_data_mask  ),      

               .pe16__std__lane17_strm1_ready         ( pe16__std__lane17_strm1_ready      ),      
               .std__pe16__lane17_strm1_cntl          ( std__pe16__lane17_strm1_cntl       ),      
               .std__pe16__lane17_strm1_data          ( std__pe16__lane17_strm1_data       ),      
               .std__pe16__lane17_strm1_data_valid    ( std__pe16__lane17_strm1_data_valid ),      
               .std__pe16__lane17_strm1_data_mask     ( std__pe16__lane17_strm1_data_mask  ),      

               // PE 16, Lane 18                 
               .pe16__std__lane18_strm0_ready         ( pe16__std__lane18_strm0_ready      ),      
               .std__pe16__lane18_strm0_cntl          ( std__pe16__lane18_strm0_cntl       ),      
               .std__pe16__lane18_strm0_data          ( std__pe16__lane18_strm0_data       ),      
               .std__pe16__lane18_strm0_data_valid    ( std__pe16__lane18_strm0_data_valid ),      
               .std__pe16__lane18_strm0_data_mask     ( std__pe16__lane18_strm0_data_mask  ),      

               .pe16__std__lane18_strm1_ready         ( pe16__std__lane18_strm1_ready      ),      
               .std__pe16__lane18_strm1_cntl          ( std__pe16__lane18_strm1_cntl       ),      
               .std__pe16__lane18_strm1_data          ( std__pe16__lane18_strm1_data       ),      
               .std__pe16__lane18_strm1_data_valid    ( std__pe16__lane18_strm1_data_valid ),      
               .std__pe16__lane18_strm1_data_mask     ( std__pe16__lane18_strm1_data_mask  ),      

               // PE 16, Lane 19                 
               .pe16__std__lane19_strm0_ready         ( pe16__std__lane19_strm0_ready      ),      
               .std__pe16__lane19_strm0_cntl          ( std__pe16__lane19_strm0_cntl       ),      
               .std__pe16__lane19_strm0_data          ( std__pe16__lane19_strm0_data       ),      
               .std__pe16__lane19_strm0_data_valid    ( std__pe16__lane19_strm0_data_valid ),      
               .std__pe16__lane19_strm0_data_mask     ( std__pe16__lane19_strm0_data_mask  ),      

               .pe16__std__lane19_strm1_ready         ( pe16__std__lane19_strm1_ready      ),      
               .std__pe16__lane19_strm1_cntl          ( std__pe16__lane19_strm1_cntl       ),      
               .std__pe16__lane19_strm1_data          ( std__pe16__lane19_strm1_data       ),      
               .std__pe16__lane19_strm1_data_valid    ( std__pe16__lane19_strm1_data_valid ),      
               .std__pe16__lane19_strm1_data_mask     ( std__pe16__lane19_strm1_data_mask  ),      

               // PE 16, Lane 20                 
               .pe16__std__lane20_strm0_ready         ( pe16__std__lane20_strm0_ready      ),      
               .std__pe16__lane20_strm0_cntl          ( std__pe16__lane20_strm0_cntl       ),      
               .std__pe16__lane20_strm0_data          ( std__pe16__lane20_strm0_data       ),      
               .std__pe16__lane20_strm0_data_valid    ( std__pe16__lane20_strm0_data_valid ),      
               .std__pe16__lane20_strm0_data_mask     ( std__pe16__lane20_strm0_data_mask  ),      

               .pe16__std__lane20_strm1_ready         ( pe16__std__lane20_strm1_ready      ),      
               .std__pe16__lane20_strm1_cntl          ( std__pe16__lane20_strm1_cntl       ),      
               .std__pe16__lane20_strm1_data          ( std__pe16__lane20_strm1_data       ),      
               .std__pe16__lane20_strm1_data_valid    ( std__pe16__lane20_strm1_data_valid ),      
               .std__pe16__lane20_strm1_data_mask     ( std__pe16__lane20_strm1_data_mask  ),      

               // PE 16, Lane 21                 
               .pe16__std__lane21_strm0_ready         ( pe16__std__lane21_strm0_ready      ),      
               .std__pe16__lane21_strm0_cntl          ( std__pe16__lane21_strm0_cntl       ),      
               .std__pe16__lane21_strm0_data          ( std__pe16__lane21_strm0_data       ),      
               .std__pe16__lane21_strm0_data_valid    ( std__pe16__lane21_strm0_data_valid ),      
               .std__pe16__lane21_strm0_data_mask     ( std__pe16__lane21_strm0_data_mask  ),      

               .pe16__std__lane21_strm1_ready         ( pe16__std__lane21_strm1_ready      ),      
               .std__pe16__lane21_strm1_cntl          ( std__pe16__lane21_strm1_cntl       ),      
               .std__pe16__lane21_strm1_data          ( std__pe16__lane21_strm1_data       ),      
               .std__pe16__lane21_strm1_data_valid    ( std__pe16__lane21_strm1_data_valid ),      
               .std__pe16__lane21_strm1_data_mask     ( std__pe16__lane21_strm1_data_mask  ),      

               // PE 16, Lane 22                 
               .pe16__std__lane22_strm0_ready         ( pe16__std__lane22_strm0_ready      ),      
               .std__pe16__lane22_strm0_cntl          ( std__pe16__lane22_strm0_cntl       ),      
               .std__pe16__lane22_strm0_data          ( std__pe16__lane22_strm0_data       ),      
               .std__pe16__lane22_strm0_data_valid    ( std__pe16__lane22_strm0_data_valid ),      
               .std__pe16__lane22_strm0_data_mask     ( std__pe16__lane22_strm0_data_mask  ),      

               .pe16__std__lane22_strm1_ready         ( pe16__std__lane22_strm1_ready      ),      
               .std__pe16__lane22_strm1_cntl          ( std__pe16__lane22_strm1_cntl       ),      
               .std__pe16__lane22_strm1_data          ( std__pe16__lane22_strm1_data       ),      
               .std__pe16__lane22_strm1_data_valid    ( std__pe16__lane22_strm1_data_valid ),      
               .std__pe16__lane22_strm1_data_mask     ( std__pe16__lane22_strm1_data_mask  ),      

               // PE 16, Lane 23                 
               .pe16__std__lane23_strm0_ready         ( pe16__std__lane23_strm0_ready      ),      
               .std__pe16__lane23_strm0_cntl          ( std__pe16__lane23_strm0_cntl       ),      
               .std__pe16__lane23_strm0_data          ( std__pe16__lane23_strm0_data       ),      
               .std__pe16__lane23_strm0_data_valid    ( std__pe16__lane23_strm0_data_valid ),      
               .std__pe16__lane23_strm0_data_mask     ( std__pe16__lane23_strm0_data_mask  ),      

               .pe16__std__lane23_strm1_ready         ( pe16__std__lane23_strm1_ready      ),      
               .std__pe16__lane23_strm1_cntl          ( std__pe16__lane23_strm1_cntl       ),      
               .std__pe16__lane23_strm1_data          ( std__pe16__lane23_strm1_data       ),      
               .std__pe16__lane23_strm1_data_valid    ( std__pe16__lane23_strm1_data_valid ),      
               .std__pe16__lane23_strm1_data_mask     ( std__pe16__lane23_strm1_data_mask  ),      

               // PE 16, Lane 24                 
               .pe16__std__lane24_strm0_ready         ( pe16__std__lane24_strm0_ready      ),      
               .std__pe16__lane24_strm0_cntl          ( std__pe16__lane24_strm0_cntl       ),      
               .std__pe16__lane24_strm0_data          ( std__pe16__lane24_strm0_data       ),      
               .std__pe16__lane24_strm0_data_valid    ( std__pe16__lane24_strm0_data_valid ),      
               .std__pe16__lane24_strm0_data_mask     ( std__pe16__lane24_strm0_data_mask  ),      

               .pe16__std__lane24_strm1_ready         ( pe16__std__lane24_strm1_ready      ),      
               .std__pe16__lane24_strm1_cntl          ( std__pe16__lane24_strm1_cntl       ),      
               .std__pe16__lane24_strm1_data          ( std__pe16__lane24_strm1_data       ),      
               .std__pe16__lane24_strm1_data_valid    ( std__pe16__lane24_strm1_data_valid ),      
               .std__pe16__lane24_strm1_data_mask     ( std__pe16__lane24_strm1_data_mask  ),      

               // PE 16, Lane 25                 
               .pe16__std__lane25_strm0_ready         ( pe16__std__lane25_strm0_ready      ),      
               .std__pe16__lane25_strm0_cntl          ( std__pe16__lane25_strm0_cntl       ),      
               .std__pe16__lane25_strm0_data          ( std__pe16__lane25_strm0_data       ),      
               .std__pe16__lane25_strm0_data_valid    ( std__pe16__lane25_strm0_data_valid ),      
               .std__pe16__lane25_strm0_data_mask     ( std__pe16__lane25_strm0_data_mask  ),      

               .pe16__std__lane25_strm1_ready         ( pe16__std__lane25_strm1_ready      ),      
               .std__pe16__lane25_strm1_cntl          ( std__pe16__lane25_strm1_cntl       ),      
               .std__pe16__lane25_strm1_data          ( std__pe16__lane25_strm1_data       ),      
               .std__pe16__lane25_strm1_data_valid    ( std__pe16__lane25_strm1_data_valid ),      
               .std__pe16__lane25_strm1_data_mask     ( std__pe16__lane25_strm1_data_mask  ),      

               // PE 16, Lane 26                 
               .pe16__std__lane26_strm0_ready         ( pe16__std__lane26_strm0_ready      ),      
               .std__pe16__lane26_strm0_cntl          ( std__pe16__lane26_strm0_cntl       ),      
               .std__pe16__lane26_strm0_data          ( std__pe16__lane26_strm0_data       ),      
               .std__pe16__lane26_strm0_data_valid    ( std__pe16__lane26_strm0_data_valid ),      
               .std__pe16__lane26_strm0_data_mask     ( std__pe16__lane26_strm0_data_mask  ),      

               .pe16__std__lane26_strm1_ready         ( pe16__std__lane26_strm1_ready      ),      
               .std__pe16__lane26_strm1_cntl          ( std__pe16__lane26_strm1_cntl       ),      
               .std__pe16__lane26_strm1_data          ( std__pe16__lane26_strm1_data       ),      
               .std__pe16__lane26_strm1_data_valid    ( std__pe16__lane26_strm1_data_valid ),      
               .std__pe16__lane26_strm1_data_mask     ( std__pe16__lane26_strm1_data_mask  ),      

               // PE 16, Lane 27                 
               .pe16__std__lane27_strm0_ready         ( pe16__std__lane27_strm0_ready      ),      
               .std__pe16__lane27_strm0_cntl          ( std__pe16__lane27_strm0_cntl       ),      
               .std__pe16__lane27_strm0_data          ( std__pe16__lane27_strm0_data       ),      
               .std__pe16__lane27_strm0_data_valid    ( std__pe16__lane27_strm0_data_valid ),      
               .std__pe16__lane27_strm0_data_mask     ( std__pe16__lane27_strm0_data_mask  ),      

               .pe16__std__lane27_strm1_ready         ( pe16__std__lane27_strm1_ready      ),      
               .std__pe16__lane27_strm1_cntl          ( std__pe16__lane27_strm1_cntl       ),      
               .std__pe16__lane27_strm1_data          ( std__pe16__lane27_strm1_data       ),      
               .std__pe16__lane27_strm1_data_valid    ( std__pe16__lane27_strm1_data_valid ),      
               .std__pe16__lane27_strm1_data_mask     ( std__pe16__lane27_strm1_data_mask  ),      

               // PE 16, Lane 28                 
               .pe16__std__lane28_strm0_ready         ( pe16__std__lane28_strm0_ready      ),      
               .std__pe16__lane28_strm0_cntl          ( std__pe16__lane28_strm0_cntl       ),      
               .std__pe16__lane28_strm0_data          ( std__pe16__lane28_strm0_data       ),      
               .std__pe16__lane28_strm0_data_valid    ( std__pe16__lane28_strm0_data_valid ),      
               .std__pe16__lane28_strm0_data_mask     ( std__pe16__lane28_strm0_data_mask  ),      

               .pe16__std__lane28_strm1_ready         ( pe16__std__lane28_strm1_ready      ),      
               .std__pe16__lane28_strm1_cntl          ( std__pe16__lane28_strm1_cntl       ),      
               .std__pe16__lane28_strm1_data          ( std__pe16__lane28_strm1_data       ),      
               .std__pe16__lane28_strm1_data_valid    ( std__pe16__lane28_strm1_data_valid ),      
               .std__pe16__lane28_strm1_data_mask     ( std__pe16__lane28_strm1_data_mask  ),      

               // PE 16, Lane 29                 
               .pe16__std__lane29_strm0_ready         ( pe16__std__lane29_strm0_ready      ),      
               .std__pe16__lane29_strm0_cntl          ( std__pe16__lane29_strm0_cntl       ),      
               .std__pe16__lane29_strm0_data          ( std__pe16__lane29_strm0_data       ),      
               .std__pe16__lane29_strm0_data_valid    ( std__pe16__lane29_strm0_data_valid ),      
               .std__pe16__lane29_strm0_data_mask     ( std__pe16__lane29_strm0_data_mask  ),      

               .pe16__std__lane29_strm1_ready         ( pe16__std__lane29_strm1_ready      ),      
               .std__pe16__lane29_strm1_cntl          ( std__pe16__lane29_strm1_cntl       ),      
               .std__pe16__lane29_strm1_data          ( std__pe16__lane29_strm1_data       ),      
               .std__pe16__lane29_strm1_data_valid    ( std__pe16__lane29_strm1_data_valid ),      
               .std__pe16__lane29_strm1_data_mask     ( std__pe16__lane29_strm1_data_mask  ),      

               // PE 16, Lane 30                 
               .pe16__std__lane30_strm0_ready         ( pe16__std__lane30_strm0_ready      ),      
               .std__pe16__lane30_strm0_cntl          ( std__pe16__lane30_strm0_cntl       ),      
               .std__pe16__lane30_strm0_data          ( std__pe16__lane30_strm0_data       ),      
               .std__pe16__lane30_strm0_data_valid    ( std__pe16__lane30_strm0_data_valid ),      
               .std__pe16__lane30_strm0_data_mask     ( std__pe16__lane30_strm0_data_mask  ),      

               .pe16__std__lane30_strm1_ready         ( pe16__std__lane30_strm1_ready      ),      
               .std__pe16__lane30_strm1_cntl          ( std__pe16__lane30_strm1_cntl       ),      
               .std__pe16__lane30_strm1_data          ( std__pe16__lane30_strm1_data       ),      
               .std__pe16__lane30_strm1_data_valid    ( std__pe16__lane30_strm1_data_valid ),      
               .std__pe16__lane30_strm1_data_mask     ( std__pe16__lane30_strm1_data_mask  ),      

               // PE 16, Lane 31                 
               .pe16__std__lane31_strm0_ready         ( pe16__std__lane31_strm0_ready      ),      
               .std__pe16__lane31_strm0_cntl          ( std__pe16__lane31_strm0_cntl       ),      
               .std__pe16__lane31_strm0_data          ( std__pe16__lane31_strm0_data       ),      
               .std__pe16__lane31_strm0_data_valid    ( std__pe16__lane31_strm0_data_valid ),      
               .std__pe16__lane31_strm0_data_mask     ( std__pe16__lane31_strm0_data_mask  ),      

               .pe16__std__lane31_strm1_ready         ( pe16__std__lane31_strm1_ready      ),      
               .std__pe16__lane31_strm1_cntl          ( std__pe16__lane31_strm1_cntl       ),      
               .std__pe16__lane31_strm1_data          ( std__pe16__lane31_strm1_data       ),      
               .std__pe16__lane31_strm1_data_valid    ( std__pe16__lane31_strm1_data_valid ),      
               .std__pe16__lane31_strm1_data_mask     ( std__pe16__lane31_strm1_data_mask  ),      

               // PE 17, Lane 0                 
               .pe17__std__lane0_strm0_ready         ( pe17__std__lane0_strm0_ready      ),      
               .std__pe17__lane0_strm0_cntl          ( std__pe17__lane0_strm0_cntl       ),      
               .std__pe17__lane0_strm0_data          ( std__pe17__lane0_strm0_data       ),      
               .std__pe17__lane0_strm0_data_valid    ( std__pe17__lane0_strm0_data_valid ),      
               .std__pe17__lane0_strm0_data_mask     ( std__pe17__lane0_strm0_data_mask  ),      

               .pe17__std__lane0_strm1_ready         ( pe17__std__lane0_strm1_ready      ),      
               .std__pe17__lane0_strm1_cntl          ( std__pe17__lane0_strm1_cntl       ),      
               .std__pe17__lane0_strm1_data          ( std__pe17__lane0_strm1_data       ),      
               .std__pe17__lane0_strm1_data_valid    ( std__pe17__lane0_strm1_data_valid ),      
               .std__pe17__lane0_strm1_data_mask     ( std__pe17__lane0_strm1_data_mask  ),      

               // PE 17, Lane 1                 
               .pe17__std__lane1_strm0_ready         ( pe17__std__lane1_strm0_ready      ),      
               .std__pe17__lane1_strm0_cntl          ( std__pe17__lane1_strm0_cntl       ),      
               .std__pe17__lane1_strm0_data          ( std__pe17__lane1_strm0_data       ),      
               .std__pe17__lane1_strm0_data_valid    ( std__pe17__lane1_strm0_data_valid ),      
               .std__pe17__lane1_strm0_data_mask     ( std__pe17__lane1_strm0_data_mask  ),      

               .pe17__std__lane1_strm1_ready         ( pe17__std__lane1_strm1_ready      ),      
               .std__pe17__lane1_strm1_cntl          ( std__pe17__lane1_strm1_cntl       ),      
               .std__pe17__lane1_strm1_data          ( std__pe17__lane1_strm1_data       ),      
               .std__pe17__lane1_strm1_data_valid    ( std__pe17__lane1_strm1_data_valid ),      
               .std__pe17__lane1_strm1_data_mask     ( std__pe17__lane1_strm1_data_mask  ),      

               // PE 17, Lane 2                 
               .pe17__std__lane2_strm0_ready         ( pe17__std__lane2_strm0_ready      ),      
               .std__pe17__lane2_strm0_cntl          ( std__pe17__lane2_strm0_cntl       ),      
               .std__pe17__lane2_strm0_data          ( std__pe17__lane2_strm0_data       ),      
               .std__pe17__lane2_strm0_data_valid    ( std__pe17__lane2_strm0_data_valid ),      
               .std__pe17__lane2_strm0_data_mask     ( std__pe17__lane2_strm0_data_mask  ),      

               .pe17__std__lane2_strm1_ready         ( pe17__std__lane2_strm1_ready      ),      
               .std__pe17__lane2_strm1_cntl          ( std__pe17__lane2_strm1_cntl       ),      
               .std__pe17__lane2_strm1_data          ( std__pe17__lane2_strm1_data       ),      
               .std__pe17__lane2_strm1_data_valid    ( std__pe17__lane2_strm1_data_valid ),      
               .std__pe17__lane2_strm1_data_mask     ( std__pe17__lane2_strm1_data_mask  ),      

               // PE 17, Lane 3                 
               .pe17__std__lane3_strm0_ready         ( pe17__std__lane3_strm0_ready      ),      
               .std__pe17__lane3_strm0_cntl          ( std__pe17__lane3_strm0_cntl       ),      
               .std__pe17__lane3_strm0_data          ( std__pe17__lane3_strm0_data       ),      
               .std__pe17__lane3_strm0_data_valid    ( std__pe17__lane3_strm0_data_valid ),      
               .std__pe17__lane3_strm0_data_mask     ( std__pe17__lane3_strm0_data_mask  ),      

               .pe17__std__lane3_strm1_ready         ( pe17__std__lane3_strm1_ready      ),      
               .std__pe17__lane3_strm1_cntl          ( std__pe17__lane3_strm1_cntl       ),      
               .std__pe17__lane3_strm1_data          ( std__pe17__lane3_strm1_data       ),      
               .std__pe17__lane3_strm1_data_valid    ( std__pe17__lane3_strm1_data_valid ),      
               .std__pe17__lane3_strm1_data_mask     ( std__pe17__lane3_strm1_data_mask  ),      

               // PE 17, Lane 4                 
               .pe17__std__lane4_strm0_ready         ( pe17__std__lane4_strm0_ready      ),      
               .std__pe17__lane4_strm0_cntl          ( std__pe17__lane4_strm0_cntl       ),      
               .std__pe17__lane4_strm0_data          ( std__pe17__lane4_strm0_data       ),      
               .std__pe17__lane4_strm0_data_valid    ( std__pe17__lane4_strm0_data_valid ),      
               .std__pe17__lane4_strm0_data_mask     ( std__pe17__lane4_strm0_data_mask  ),      

               .pe17__std__lane4_strm1_ready         ( pe17__std__lane4_strm1_ready      ),      
               .std__pe17__lane4_strm1_cntl          ( std__pe17__lane4_strm1_cntl       ),      
               .std__pe17__lane4_strm1_data          ( std__pe17__lane4_strm1_data       ),      
               .std__pe17__lane4_strm1_data_valid    ( std__pe17__lane4_strm1_data_valid ),      
               .std__pe17__lane4_strm1_data_mask     ( std__pe17__lane4_strm1_data_mask  ),      

               // PE 17, Lane 5                 
               .pe17__std__lane5_strm0_ready         ( pe17__std__lane5_strm0_ready      ),      
               .std__pe17__lane5_strm0_cntl          ( std__pe17__lane5_strm0_cntl       ),      
               .std__pe17__lane5_strm0_data          ( std__pe17__lane5_strm0_data       ),      
               .std__pe17__lane5_strm0_data_valid    ( std__pe17__lane5_strm0_data_valid ),      
               .std__pe17__lane5_strm0_data_mask     ( std__pe17__lane5_strm0_data_mask  ),      

               .pe17__std__lane5_strm1_ready         ( pe17__std__lane5_strm1_ready      ),      
               .std__pe17__lane5_strm1_cntl          ( std__pe17__lane5_strm1_cntl       ),      
               .std__pe17__lane5_strm1_data          ( std__pe17__lane5_strm1_data       ),      
               .std__pe17__lane5_strm1_data_valid    ( std__pe17__lane5_strm1_data_valid ),      
               .std__pe17__lane5_strm1_data_mask     ( std__pe17__lane5_strm1_data_mask  ),      

               // PE 17, Lane 6                 
               .pe17__std__lane6_strm0_ready         ( pe17__std__lane6_strm0_ready      ),      
               .std__pe17__lane6_strm0_cntl          ( std__pe17__lane6_strm0_cntl       ),      
               .std__pe17__lane6_strm0_data          ( std__pe17__lane6_strm0_data       ),      
               .std__pe17__lane6_strm0_data_valid    ( std__pe17__lane6_strm0_data_valid ),      
               .std__pe17__lane6_strm0_data_mask     ( std__pe17__lane6_strm0_data_mask  ),      

               .pe17__std__lane6_strm1_ready         ( pe17__std__lane6_strm1_ready      ),      
               .std__pe17__lane6_strm1_cntl          ( std__pe17__lane6_strm1_cntl       ),      
               .std__pe17__lane6_strm1_data          ( std__pe17__lane6_strm1_data       ),      
               .std__pe17__lane6_strm1_data_valid    ( std__pe17__lane6_strm1_data_valid ),      
               .std__pe17__lane6_strm1_data_mask     ( std__pe17__lane6_strm1_data_mask  ),      

               // PE 17, Lane 7                 
               .pe17__std__lane7_strm0_ready         ( pe17__std__lane7_strm0_ready      ),      
               .std__pe17__lane7_strm0_cntl          ( std__pe17__lane7_strm0_cntl       ),      
               .std__pe17__lane7_strm0_data          ( std__pe17__lane7_strm0_data       ),      
               .std__pe17__lane7_strm0_data_valid    ( std__pe17__lane7_strm0_data_valid ),      
               .std__pe17__lane7_strm0_data_mask     ( std__pe17__lane7_strm0_data_mask  ),      

               .pe17__std__lane7_strm1_ready         ( pe17__std__lane7_strm1_ready      ),      
               .std__pe17__lane7_strm1_cntl          ( std__pe17__lane7_strm1_cntl       ),      
               .std__pe17__lane7_strm1_data          ( std__pe17__lane7_strm1_data       ),      
               .std__pe17__lane7_strm1_data_valid    ( std__pe17__lane7_strm1_data_valid ),      
               .std__pe17__lane7_strm1_data_mask     ( std__pe17__lane7_strm1_data_mask  ),      

               // PE 17, Lane 8                 
               .pe17__std__lane8_strm0_ready         ( pe17__std__lane8_strm0_ready      ),      
               .std__pe17__lane8_strm0_cntl          ( std__pe17__lane8_strm0_cntl       ),      
               .std__pe17__lane8_strm0_data          ( std__pe17__lane8_strm0_data       ),      
               .std__pe17__lane8_strm0_data_valid    ( std__pe17__lane8_strm0_data_valid ),      
               .std__pe17__lane8_strm0_data_mask     ( std__pe17__lane8_strm0_data_mask  ),      

               .pe17__std__lane8_strm1_ready         ( pe17__std__lane8_strm1_ready      ),      
               .std__pe17__lane8_strm1_cntl          ( std__pe17__lane8_strm1_cntl       ),      
               .std__pe17__lane8_strm1_data          ( std__pe17__lane8_strm1_data       ),      
               .std__pe17__lane8_strm1_data_valid    ( std__pe17__lane8_strm1_data_valid ),      
               .std__pe17__lane8_strm1_data_mask     ( std__pe17__lane8_strm1_data_mask  ),      

               // PE 17, Lane 9                 
               .pe17__std__lane9_strm0_ready         ( pe17__std__lane9_strm0_ready      ),      
               .std__pe17__lane9_strm0_cntl          ( std__pe17__lane9_strm0_cntl       ),      
               .std__pe17__lane9_strm0_data          ( std__pe17__lane9_strm0_data       ),      
               .std__pe17__lane9_strm0_data_valid    ( std__pe17__lane9_strm0_data_valid ),      
               .std__pe17__lane9_strm0_data_mask     ( std__pe17__lane9_strm0_data_mask  ),      

               .pe17__std__lane9_strm1_ready         ( pe17__std__lane9_strm1_ready      ),      
               .std__pe17__lane9_strm1_cntl          ( std__pe17__lane9_strm1_cntl       ),      
               .std__pe17__lane9_strm1_data          ( std__pe17__lane9_strm1_data       ),      
               .std__pe17__lane9_strm1_data_valid    ( std__pe17__lane9_strm1_data_valid ),      
               .std__pe17__lane9_strm1_data_mask     ( std__pe17__lane9_strm1_data_mask  ),      

               // PE 17, Lane 10                 
               .pe17__std__lane10_strm0_ready         ( pe17__std__lane10_strm0_ready      ),      
               .std__pe17__lane10_strm0_cntl          ( std__pe17__lane10_strm0_cntl       ),      
               .std__pe17__lane10_strm0_data          ( std__pe17__lane10_strm0_data       ),      
               .std__pe17__lane10_strm0_data_valid    ( std__pe17__lane10_strm0_data_valid ),      
               .std__pe17__lane10_strm0_data_mask     ( std__pe17__lane10_strm0_data_mask  ),      

               .pe17__std__lane10_strm1_ready         ( pe17__std__lane10_strm1_ready      ),      
               .std__pe17__lane10_strm1_cntl          ( std__pe17__lane10_strm1_cntl       ),      
               .std__pe17__lane10_strm1_data          ( std__pe17__lane10_strm1_data       ),      
               .std__pe17__lane10_strm1_data_valid    ( std__pe17__lane10_strm1_data_valid ),      
               .std__pe17__lane10_strm1_data_mask     ( std__pe17__lane10_strm1_data_mask  ),      

               // PE 17, Lane 11                 
               .pe17__std__lane11_strm0_ready         ( pe17__std__lane11_strm0_ready      ),      
               .std__pe17__lane11_strm0_cntl          ( std__pe17__lane11_strm0_cntl       ),      
               .std__pe17__lane11_strm0_data          ( std__pe17__lane11_strm0_data       ),      
               .std__pe17__lane11_strm0_data_valid    ( std__pe17__lane11_strm0_data_valid ),      
               .std__pe17__lane11_strm0_data_mask     ( std__pe17__lane11_strm0_data_mask  ),      

               .pe17__std__lane11_strm1_ready         ( pe17__std__lane11_strm1_ready      ),      
               .std__pe17__lane11_strm1_cntl          ( std__pe17__lane11_strm1_cntl       ),      
               .std__pe17__lane11_strm1_data          ( std__pe17__lane11_strm1_data       ),      
               .std__pe17__lane11_strm1_data_valid    ( std__pe17__lane11_strm1_data_valid ),      
               .std__pe17__lane11_strm1_data_mask     ( std__pe17__lane11_strm1_data_mask  ),      

               // PE 17, Lane 12                 
               .pe17__std__lane12_strm0_ready         ( pe17__std__lane12_strm0_ready      ),      
               .std__pe17__lane12_strm0_cntl          ( std__pe17__lane12_strm0_cntl       ),      
               .std__pe17__lane12_strm0_data          ( std__pe17__lane12_strm0_data       ),      
               .std__pe17__lane12_strm0_data_valid    ( std__pe17__lane12_strm0_data_valid ),      
               .std__pe17__lane12_strm0_data_mask     ( std__pe17__lane12_strm0_data_mask  ),      

               .pe17__std__lane12_strm1_ready         ( pe17__std__lane12_strm1_ready      ),      
               .std__pe17__lane12_strm1_cntl          ( std__pe17__lane12_strm1_cntl       ),      
               .std__pe17__lane12_strm1_data          ( std__pe17__lane12_strm1_data       ),      
               .std__pe17__lane12_strm1_data_valid    ( std__pe17__lane12_strm1_data_valid ),      
               .std__pe17__lane12_strm1_data_mask     ( std__pe17__lane12_strm1_data_mask  ),      

               // PE 17, Lane 13                 
               .pe17__std__lane13_strm0_ready         ( pe17__std__lane13_strm0_ready      ),      
               .std__pe17__lane13_strm0_cntl          ( std__pe17__lane13_strm0_cntl       ),      
               .std__pe17__lane13_strm0_data          ( std__pe17__lane13_strm0_data       ),      
               .std__pe17__lane13_strm0_data_valid    ( std__pe17__lane13_strm0_data_valid ),      
               .std__pe17__lane13_strm0_data_mask     ( std__pe17__lane13_strm0_data_mask  ),      

               .pe17__std__lane13_strm1_ready         ( pe17__std__lane13_strm1_ready      ),      
               .std__pe17__lane13_strm1_cntl          ( std__pe17__lane13_strm1_cntl       ),      
               .std__pe17__lane13_strm1_data          ( std__pe17__lane13_strm1_data       ),      
               .std__pe17__lane13_strm1_data_valid    ( std__pe17__lane13_strm1_data_valid ),      
               .std__pe17__lane13_strm1_data_mask     ( std__pe17__lane13_strm1_data_mask  ),      

               // PE 17, Lane 14                 
               .pe17__std__lane14_strm0_ready         ( pe17__std__lane14_strm0_ready      ),      
               .std__pe17__lane14_strm0_cntl          ( std__pe17__lane14_strm0_cntl       ),      
               .std__pe17__lane14_strm0_data          ( std__pe17__lane14_strm0_data       ),      
               .std__pe17__lane14_strm0_data_valid    ( std__pe17__lane14_strm0_data_valid ),      
               .std__pe17__lane14_strm0_data_mask     ( std__pe17__lane14_strm0_data_mask  ),      

               .pe17__std__lane14_strm1_ready         ( pe17__std__lane14_strm1_ready      ),      
               .std__pe17__lane14_strm1_cntl          ( std__pe17__lane14_strm1_cntl       ),      
               .std__pe17__lane14_strm1_data          ( std__pe17__lane14_strm1_data       ),      
               .std__pe17__lane14_strm1_data_valid    ( std__pe17__lane14_strm1_data_valid ),      
               .std__pe17__lane14_strm1_data_mask     ( std__pe17__lane14_strm1_data_mask  ),      

               // PE 17, Lane 15                 
               .pe17__std__lane15_strm0_ready         ( pe17__std__lane15_strm0_ready      ),      
               .std__pe17__lane15_strm0_cntl          ( std__pe17__lane15_strm0_cntl       ),      
               .std__pe17__lane15_strm0_data          ( std__pe17__lane15_strm0_data       ),      
               .std__pe17__lane15_strm0_data_valid    ( std__pe17__lane15_strm0_data_valid ),      
               .std__pe17__lane15_strm0_data_mask     ( std__pe17__lane15_strm0_data_mask  ),      

               .pe17__std__lane15_strm1_ready         ( pe17__std__lane15_strm1_ready      ),      
               .std__pe17__lane15_strm1_cntl          ( std__pe17__lane15_strm1_cntl       ),      
               .std__pe17__lane15_strm1_data          ( std__pe17__lane15_strm1_data       ),      
               .std__pe17__lane15_strm1_data_valid    ( std__pe17__lane15_strm1_data_valid ),      
               .std__pe17__lane15_strm1_data_mask     ( std__pe17__lane15_strm1_data_mask  ),      

               // PE 17, Lane 16                 
               .pe17__std__lane16_strm0_ready         ( pe17__std__lane16_strm0_ready      ),      
               .std__pe17__lane16_strm0_cntl          ( std__pe17__lane16_strm0_cntl       ),      
               .std__pe17__lane16_strm0_data          ( std__pe17__lane16_strm0_data       ),      
               .std__pe17__lane16_strm0_data_valid    ( std__pe17__lane16_strm0_data_valid ),      
               .std__pe17__lane16_strm0_data_mask     ( std__pe17__lane16_strm0_data_mask  ),      

               .pe17__std__lane16_strm1_ready         ( pe17__std__lane16_strm1_ready      ),      
               .std__pe17__lane16_strm1_cntl          ( std__pe17__lane16_strm1_cntl       ),      
               .std__pe17__lane16_strm1_data          ( std__pe17__lane16_strm1_data       ),      
               .std__pe17__lane16_strm1_data_valid    ( std__pe17__lane16_strm1_data_valid ),      
               .std__pe17__lane16_strm1_data_mask     ( std__pe17__lane16_strm1_data_mask  ),      

               // PE 17, Lane 17                 
               .pe17__std__lane17_strm0_ready         ( pe17__std__lane17_strm0_ready      ),      
               .std__pe17__lane17_strm0_cntl          ( std__pe17__lane17_strm0_cntl       ),      
               .std__pe17__lane17_strm0_data          ( std__pe17__lane17_strm0_data       ),      
               .std__pe17__lane17_strm0_data_valid    ( std__pe17__lane17_strm0_data_valid ),      
               .std__pe17__lane17_strm0_data_mask     ( std__pe17__lane17_strm0_data_mask  ),      

               .pe17__std__lane17_strm1_ready         ( pe17__std__lane17_strm1_ready      ),      
               .std__pe17__lane17_strm1_cntl          ( std__pe17__lane17_strm1_cntl       ),      
               .std__pe17__lane17_strm1_data          ( std__pe17__lane17_strm1_data       ),      
               .std__pe17__lane17_strm1_data_valid    ( std__pe17__lane17_strm1_data_valid ),      
               .std__pe17__lane17_strm1_data_mask     ( std__pe17__lane17_strm1_data_mask  ),      

               // PE 17, Lane 18                 
               .pe17__std__lane18_strm0_ready         ( pe17__std__lane18_strm0_ready      ),      
               .std__pe17__lane18_strm0_cntl          ( std__pe17__lane18_strm0_cntl       ),      
               .std__pe17__lane18_strm0_data          ( std__pe17__lane18_strm0_data       ),      
               .std__pe17__lane18_strm0_data_valid    ( std__pe17__lane18_strm0_data_valid ),      
               .std__pe17__lane18_strm0_data_mask     ( std__pe17__lane18_strm0_data_mask  ),      

               .pe17__std__lane18_strm1_ready         ( pe17__std__lane18_strm1_ready      ),      
               .std__pe17__lane18_strm1_cntl          ( std__pe17__lane18_strm1_cntl       ),      
               .std__pe17__lane18_strm1_data          ( std__pe17__lane18_strm1_data       ),      
               .std__pe17__lane18_strm1_data_valid    ( std__pe17__lane18_strm1_data_valid ),      
               .std__pe17__lane18_strm1_data_mask     ( std__pe17__lane18_strm1_data_mask  ),      

               // PE 17, Lane 19                 
               .pe17__std__lane19_strm0_ready         ( pe17__std__lane19_strm0_ready      ),      
               .std__pe17__lane19_strm0_cntl          ( std__pe17__lane19_strm0_cntl       ),      
               .std__pe17__lane19_strm0_data          ( std__pe17__lane19_strm0_data       ),      
               .std__pe17__lane19_strm0_data_valid    ( std__pe17__lane19_strm0_data_valid ),      
               .std__pe17__lane19_strm0_data_mask     ( std__pe17__lane19_strm0_data_mask  ),      

               .pe17__std__lane19_strm1_ready         ( pe17__std__lane19_strm1_ready      ),      
               .std__pe17__lane19_strm1_cntl          ( std__pe17__lane19_strm1_cntl       ),      
               .std__pe17__lane19_strm1_data          ( std__pe17__lane19_strm1_data       ),      
               .std__pe17__lane19_strm1_data_valid    ( std__pe17__lane19_strm1_data_valid ),      
               .std__pe17__lane19_strm1_data_mask     ( std__pe17__lane19_strm1_data_mask  ),      

               // PE 17, Lane 20                 
               .pe17__std__lane20_strm0_ready         ( pe17__std__lane20_strm0_ready      ),      
               .std__pe17__lane20_strm0_cntl          ( std__pe17__lane20_strm0_cntl       ),      
               .std__pe17__lane20_strm0_data          ( std__pe17__lane20_strm0_data       ),      
               .std__pe17__lane20_strm0_data_valid    ( std__pe17__lane20_strm0_data_valid ),      
               .std__pe17__lane20_strm0_data_mask     ( std__pe17__lane20_strm0_data_mask  ),      

               .pe17__std__lane20_strm1_ready         ( pe17__std__lane20_strm1_ready      ),      
               .std__pe17__lane20_strm1_cntl          ( std__pe17__lane20_strm1_cntl       ),      
               .std__pe17__lane20_strm1_data          ( std__pe17__lane20_strm1_data       ),      
               .std__pe17__lane20_strm1_data_valid    ( std__pe17__lane20_strm1_data_valid ),      
               .std__pe17__lane20_strm1_data_mask     ( std__pe17__lane20_strm1_data_mask  ),      

               // PE 17, Lane 21                 
               .pe17__std__lane21_strm0_ready         ( pe17__std__lane21_strm0_ready      ),      
               .std__pe17__lane21_strm0_cntl          ( std__pe17__lane21_strm0_cntl       ),      
               .std__pe17__lane21_strm0_data          ( std__pe17__lane21_strm0_data       ),      
               .std__pe17__lane21_strm0_data_valid    ( std__pe17__lane21_strm0_data_valid ),      
               .std__pe17__lane21_strm0_data_mask     ( std__pe17__lane21_strm0_data_mask  ),      

               .pe17__std__lane21_strm1_ready         ( pe17__std__lane21_strm1_ready      ),      
               .std__pe17__lane21_strm1_cntl          ( std__pe17__lane21_strm1_cntl       ),      
               .std__pe17__lane21_strm1_data          ( std__pe17__lane21_strm1_data       ),      
               .std__pe17__lane21_strm1_data_valid    ( std__pe17__lane21_strm1_data_valid ),      
               .std__pe17__lane21_strm1_data_mask     ( std__pe17__lane21_strm1_data_mask  ),      

               // PE 17, Lane 22                 
               .pe17__std__lane22_strm0_ready         ( pe17__std__lane22_strm0_ready      ),      
               .std__pe17__lane22_strm0_cntl          ( std__pe17__lane22_strm0_cntl       ),      
               .std__pe17__lane22_strm0_data          ( std__pe17__lane22_strm0_data       ),      
               .std__pe17__lane22_strm0_data_valid    ( std__pe17__lane22_strm0_data_valid ),      
               .std__pe17__lane22_strm0_data_mask     ( std__pe17__lane22_strm0_data_mask  ),      

               .pe17__std__lane22_strm1_ready         ( pe17__std__lane22_strm1_ready      ),      
               .std__pe17__lane22_strm1_cntl          ( std__pe17__lane22_strm1_cntl       ),      
               .std__pe17__lane22_strm1_data          ( std__pe17__lane22_strm1_data       ),      
               .std__pe17__lane22_strm1_data_valid    ( std__pe17__lane22_strm1_data_valid ),      
               .std__pe17__lane22_strm1_data_mask     ( std__pe17__lane22_strm1_data_mask  ),      

               // PE 17, Lane 23                 
               .pe17__std__lane23_strm0_ready         ( pe17__std__lane23_strm0_ready      ),      
               .std__pe17__lane23_strm0_cntl          ( std__pe17__lane23_strm0_cntl       ),      
               .std__pe17__lane23_strm0_data          ( std__pe17__lane23_strm0_data       ),      
               .std__pe17__lane23_strm0_data_valid    ( std__pe17__lane23_strm0_data_valid ),      
               .std__pe17__lane23_strm0_data_mask     ( std__pe17__lane23_strm0_data_mask  ),      

               .pe17__std__lane23_strm1_ready         ( pe17__std__lane23_strm1_ready      ),      
               .std__pe17__lane23_strm1_cntl          ( std__pe17__lane23_strm1_cntl       ),      
               .std__pe17__lane23_strm1_data          ( std__pe17__lane23_strm1_data       ),      
               .std__pe17__lane23_strm1_data_valid    ( std__pe17__lane23_strm1_data_valid ),      
               .std__pe17__lane23_strm1_data_mask     ( std__pe17__lane23_strm1_data_mask  ),      

               // PE 17, Lane 24                 
               .pe17__std__lane24_strm0_ready         ( pe17__std__lane24_strm0_ready      ),      
               .std__pe17__lane24_strm0_cntl          ( std__pe17__lane24_strm0_cntl       ),      
               .std__pe17__lane24_strm0_data          ( std__pe17__lane24_strm0_data       ),      
               .std__pe17__lane24_strm0_data_valid    ( std__pe17__lane24_strm0_data_valid ),      
               .std__pe17__lane24_strm0_data_mask     ( std__pe17__lane24_strm0_data_mask  ),      

               .pe17__std__lane24_strm1_ready         ( pe17__std__lane24_strm1_ready      ),      
               .std__pe17__lane24_strm1_cntl          ( std__pe17__lane24_strm1_cntl       ),      
               .std__pe17__lane24_strm1_data          ( std__pe17__lane24_strm1_data       ),      
               .std__pe17__lane24_strm1_data_valid    ( std__pe17__lane24_strm1_data_valid ),      
               .std__pe17__lane24_strm1_data_mask     ( std__pe17__lane24_strm1_data_mask  ),      

               // PE 17, Lane 25                 
               .pe17__std__lane25_strm0_ready         ( pe17__std__lane25_strm0_ready      ),      
               .std__pe17__lane25_strm0_cntl          ( std__pe17__lane25_strm0_cntl       ),      
               .std__pe17__lane25_strm0_data          ( std__pe17__lane25_strm0_data       ),      
               .std__pe17__lane25_strm0_data_valid    ( std__pe17__lane25_strm0_data_valid ),      
               .std__pe17__lane25_strm0_data_mask     ( std__pe17__lane25_strm0_data_mask  ),      

               .pe17__std__lane25_strm1_ready         ( pe17__std__lane25_strm1_ready      ),      
               .std__pe17__lane25_strm1_cntl          ( std__pe17__lane25_strm1_cntl       ),      
               .std__pe17__lane25_strm1_data          ( std__pe17__lane25_strm1_data       ),      
               .std__pe17__lane25_strm1_data_valid    ( std__pe17__lane25_strm1_data_valid ),      
               .std__pe17__lane25_strm1_data_mask     ( std__pe17__lane25_strm1_data_mask  ),      

               // PE 17, Lane 26                 
               .pe17__std__lane26_strm0_ready         ( pe17__std__lane26_strm0_ready      ),      
               .std__pe17__lane26_strm0_cntl          ( std__pe17__lane26_strm0_cntl       ),      
               .std__pe17__lane26_strm0_data          ( std__pe17__lane26_strm0_data       ),      
               .std__pe17__lane26_strm0_data_valid    ( std__pe17__lane26_strm0_data_valid ),      
               .std__pe17__lane26_strm0_data_mask     ( std__pe17__lane26_strm0_data_mask  ),      

               .pe17__std__lane26_strm1_ready         ( pe17__std__lane26_strm1_ready      ),      
               .std__pe17__lane26_strm1_cntl          ( std__pe17__lane26_strm1_cntl       ),      
               .std__pe17__lane26_strm1_data          ( std__pe17__lane26_strm1_data       ),      
               .std__pe17__lane26_strm1_data_valid    ( std__pe17__lane26_strm1_data_valid ),      
               .std__pe17__lane26_strm1_data_mask     ( std__pe17__lane26_strm1_data_mask  ),      

               // PE 17, Lane 27                 
               .pe17__std__lane27_strm0_ready         ( pe17__std__lane27_strm0_ready      ),      
               .std__pe17__lane27_strm0_cntl          ( std__pe17__lane27_strm0_cntl       ),      
               .std__pe17__lane27_strm0_data          ( std__pe17__lane27_strm0_data       ),      
               .std__pe17__lane27_strm0_data_valid    ( std__pe17__lane27_strm0_data_valid ),      
               .std__pe17__lane27_strm0_data_mask     ( std__pe17__lane27_strm0_data_mask  ),      

               .pe17__std__lane27_strm1_ready         ( pe17__std__lane27_strm1_ready      ),      
               .std__pe17__lane27_strm1_cntl          ( std__pe17__lane27_strm1_cntl       ),      
               .std__pe17__lane27_strm1_data          ( std__pe17__lane27_strm1_data       ),      
               .std__pe17__lane27_strm1_data_valid    ( std__pe17__lane27_strm1_data_valid ),      
               .std__pe17__lane27_strm1_data_mask     ( std__pe17__lane27_strm1_data_mask  ),      

               // PE 17, Lane 28                 
               .pe17__std__lane28_strm0_ready         ( pe17__std__lane28_strm0_ready      ),      
               .std__pe17__lane28_strm0_cntl          ( std__pe17__lane28_strm0_cntl       ),      
               .std__pe17__lane28_strm0_data          ( std__pe17__lane28_strm0_data       ),      
               .std__pe17__lane28_strm0_data_valid    ( std__pe17__lane28_strm0_data_valid ),      
               .std__pe17__lane28_strm0_data_mask     ( std__pe17__lane28_strm0_data_mask  ),      

               .pe17__std__lane28_strm1_ready         ( pe17__std__lane28_strm1_ready      ),      
               .std__pe17__lane28_strm1_cntl          ( std__pe17__lane28_strm1_cntl       ),      
               .std__pe17__lane28_strm1_data          ( std__pe17__lane28_strm1_data       ),      
               .std__pe17__lane28_strm1_data_valid    ( std__pe17__lane28_strm1_data_valid ),      
               .std__pe17__lane28_strm1_data_mask     ( std__pe17__lane28_strm1_data_mask  ),      

               // PE 17, Lane 29                 
               .pe17__std__lane29_strm0_ready         ( pe17__std__lane29_strm0_ready      ),      
               .std__pe17__lane29_strm0_cntl          ( std__pe17__lane29_strm0_cntl       ),      
               .std__pe17__lane29_strm0_data          ( std__pe17__lane29_strm0_data       ),      
               .std__pe17__lane29_strm0_data_valid    ( std__pe17__lane29_strm0_data_valid ),      
               .std__pe17__lane29_strm0_data_mask     ( std__pe17__lane29_strm0_data_mask  ),      

               .pe17__std__lane29_strm1_ready         ( pe17__std__lane29_strm1_ready      ),      
               .std__pe17__lane29_strm1_cntl          ( std__pe17__lane29_strm1_cntl       ),      
               .std__pe17__lane29_strm1_data          ( std__pe17__lane29_strm1_data       ),      
               .std__pe17__lane29_strm1_data_valid    ( std__pe17__lane29_strm1_data_valid ),      
               .std__pe17__lane29_strm1_data_mask     ( std__pe17__lane29_strm1_data_mask  ),      

               // PE 17, Lane 30                 
               .pe17__std__lane30_strm0_ready         ( pe17__std__lane30_strm0_ready      ),      
               .std__pe17__lane30_strm0_cntl          ( std__pe17__lane30_strm0_cntl       ),      
               .std__pe17__lane30_strm0_data          ( std__pe17__lane30_strm0_data       ),      
               .std__pe17__lane30_strm0_data_valid    ( std__pe17__lane30_strm0_data_valid ),      
               .std__pe17__lane30_strm0_data_mask     ( std__pe17__lane30_strm0_data_mask  ),      

               .pe17__std__lane30_strm1_ready         ( pe17__std__lane30_strm1_ready      ),      
               .std__pe17__lane30_strm1_cntl          ( std__pe17__lane30_strm1_cntl       ),      
               .std__pe17__lane30_strm1_data          ( std__pe17__lane30_strm1_data       ),      
               .std__pe17__lane30_strm1_data_valid    ( std__pe17__lane30_strm1_data_valid ),      
               .std__pe17__lane30_strm1_data_mask     ( std__pe17__lane30_strm1_data_mask  ),      

               // PE 17, Lane 31                 
               .pe17__std__lane31_strm0_ready         ( pe17__std__lane31_strm0_ready      ),      
               .std__pe17__lane31_strm0_cntl          ( std__pe17__lane31_strm0_cntl       ),      
               .std__pe17__lane31_strm0_data          ( std__pe17__lane31_strm0_data       ),      
               .std__pe17__lane31_strm0_data_valid    ( std__pe17__lane31_strm0_data_valid ),      
               .std__pe17__lane31_strm0_data_mask     ( std__pe17__lane31_strm0_data_mask  ),      

               .pe17__std__lane31_strm1_ready         ( pe17__std__lane31_strm1_ready      ),      
               .std__pe17__lane31_strm1_cntl          ( std__pe17__lane31_strm1_cntl       ),      
               .std__pe17__lane31_strm1_data          ( std__pe17__lane31_strm1_data       ),      
               .std__pe17__lane31_strm1_data_valid    ( std__pe17__lane31_strm1_data_valid ),      
               .std__pe17__lane31_strm1_data_mask     ( std__pe17__lane31_strm1_data_mask  ),      

               // PE 18, Lane 0                 
               .pe18__std__lane0_strm0_ready         ( pe18__std__lane0_strm0_ready      ),      
               .std__pe18__lane0_strm0_cntl          ( std__pe18__lane0_strm0_cntl       ),      
               .std__pe18__lane0_strm0_data          ( std__pe18__lane0_strm0_data       ),      
               .std__pe18__lane0_strm0_data_valid    ( std__pe18__lane0_strm0_data_valid ),      
               .std__pe18__lane0_strm0_data_mask     ( std__pe18__lane0_strm0_data_mask  ),      

               .pe18__std__lane0_strm1_ready         ( pe18__std__lane0_strm1_ready      ),      
               .std__pe18__lane0_strm1_cntl          ( std__pe18__lane0_strm1_cntl       ),      
               .std__pe18__lane0_strm1_data          ( std__pe18__lane0_strm1_data       ),      
               .std__pe18__lane0_strm1_data_valid    ( std__pe18__lane0_strm1_data_valid ),      
               .std__pe18__lane0_strm1_data_mask     ( std__pe18__lane0_strm1_data_mask  ),      

               // PE 18, Lane 1                 
               .pe18__std__lane1_strm0_ready         ( pe18__std__lane1_strm0_ready      ),      
               .std__pe18__lane1_strm0_cntl          ( std__pe18__lane1_strm0_cntl       ),      
               .std__pe18__lane1_strm0_data          ( std__pe18__lane1_strm0_data       ),      
               .std__pe18__lane1_strm0_data_valid    ( std__pe18__lane1_strm0_data_valid ),      
               .std__pe18__lane1_strm0_data_mask     ( std__pe18__lane1_strm0_data_mask  ),      

               .pe18__std__lane1_strm1_ready         ( pe18__std__lane1_strm1_ready      ),      
               .std__pe18__lane1_strm1_cntl          ( std__pe18__lane1_strm1_cntl       ),      
               .std__pe18__lane1_strm1_data          ( std__pe18__lane1_strm1_data       ),      
               .std__pe18__lane1_strm1_data_valid    ( std__pe18__lane1_strm1_data_valid ),      
               .std__pe18__lane1_strm1_data_mask     ( std__pe18__lane1_strm1_data_mask  ),      

               // PE 18, Lane 2                 
               .pe18__std__lane2_strm0_ready         ( pe18__std__lane2_strm0_ready      ),      
               .std__pe18__lane2_strm0_cntl          ( std__pe18__lane2_strm0_cntl       ),      
               .std__pe18__lane2_strm0_data          ( std__pe18__lane2_strm0_data       ),      
               .std__pe18__lane2_strm0_data_valid    ( std__pe18__lane2_strm0_data_valid ),      
               .std__pe18__lane2_strm0_data_mask     ( std__pe18__lane2_strm0_data_mask  ),      

               .pe18__std__lane2_strm1_ready         ( pe18__std__lane2_strm1_ready      ),      
               .std__pe18__lane2_strm1_cntl          ( std__pe18__lane2_strm1_cntl       ),      
               .std__pe18__lane2_strm1_data          ( std__pe18__lane2_strm1_data       ),      
               .std__pe18__lane2_strm1_data_valid    ( std__pe18__lane2_strm1_data_valid ),      
               .std__pe18__lane2_strm1_data_mask     ( std__pe18__lane2_strm1_data_mask  ),      

               // PE 18, Lane 3                 
               .pe18__std__lane3_strm0_ready         ( pe18__std__lane3_strm0_ready      ),      
               .std__pe18__lane3_strm0_cntl          ( std__pe18__lane3_strm0_cntl       ),      
               .std__pe18__lane3_strm0_data          ( std__pe18__lane3_strm0_data       ),      
               .std__pe18__lane3_strm0_data_valid    ( std__pe18__lane3_strm0_data_valid ),      
               .std__pe18__lane3_strm0_data_mask     ( std__pe18__lane3_strm0_data_mask  ),      

               .pe18__std__lane3_strm1_ready         ( pe18__std__lane3_strm1_ready      ),      
               .std__pe18__lane3_strm1_cntl          ( std__pe18__lane3_strm1_cntl       ),      
               .std__pe18__lane3_strm1_data          ( std__pe18__lane3_strm1_data       ),      
               .std__pe18__lane3_strm1_data_valid    ( std__pe18__lane3_strm1_data_valid ),      
               .std__pe18__lane3_strm1_data_mask     ( std__pe18__lane3_strm1_data_mask  ),      

               // PE 18, Lane 4                 
               .pe18__std__lane4_strm0_ready         ( pe18__std__lane4_strm0_ready      ),      
               .std__pe18__lane4_strm0_cntl          ( std__pe18__lane4_strm0_cntl       ),      
               .std__pe18__lane4_strm0_data          ( std__pe18__lane4_strm0_data       ),      
               .std__pe18__lane4_strm0_data_valid    ( std__pe18__lane4_strm0_data_valid ),      
               .std__pe18__lane4_strm0_data_mask     ( std__pe18__lane4_strm0_data_mask  ),      

               .pe18__std__lane4_strm1_ready         ( pe18__std__lane4_strm1_ready      ),      
               .std__pe18__lane4_strm1_cntl          ( std__pe18__lane4_strm1_cntl       ),      
               .std__pe18__lane4_strm1_data          ( std__pe18__lane4_strm1_data       ),      
               .std__pe18__lane4_strm1_data_valid    ( std__pe18__lane4_strm1_data_valid ),      
               .std__pe18__lane4_strm1_data_mask     ( std__pe18__lane4_strm1_data_mask  ),      

               // PE 18, Lane 5                 
               .pe18__std__lane5_strm0_ready         ( pe18__std__lane5_strm0_ready      ),      
               .std__pe18__lane5_strm0_cntl          ( std__pe18__lane5_strm0_cntl       ),      
               .std__pe18__lane5_strm0_data          ( std__pe18__lane5_strm0_data       ),      
               .std__pe18__lane5_strm0_data_valid    ( std__pe18__lane5_strm0_data_valid ),      
               .std__pe18__lane5_strm0_data_mask     ( std__pe18__lane5_strm0_data_mask  ),      

               .pe18__std__lane5_strm1_ready         ( pe18__std__lane5_strm1_ready      ),      
               .std__pe18__lane5_strm1_cntl          ( std__pe18__lane5_strm1_cntl       ),      
               .std__pe18__lane5_strm1_data          ( std__pe18__lane5_strm1_data       ),      
               .std__pe18__lane5_strm1_data_valid    ( std__pe18__lane5_strm1_data_valid ),      
               .std__pe18__lane5_strm1_data_mask     ( std__pe18__lane5_strm1_data_mask  ),      

               // PE 18, Lane 6                 
               .pe18__std__lane6_strm0_ready         ( pe18__std__lane6_strm0_ready      ),      
               .std__pe18__lane6_strm0_cntl          ( std__pe18__lane6_strm0_cntl       ),      
               .std__pe18__lane6_strm0_data          ( std__pe18__lane6_strm0_data       ),      
               .std__pe18__lane6_strm0_data_valid    ( std__pe18__lane6_strm0_data_valid ),      
               .std__pe18__lane6_strm0_data_mask     ( std__pe18__lane6_strm0_data_mask  ),      

               .pe18__std__lane6_strm1_ready         ( pe18__std__lane6_strm1_ready      ),      
               .std__pe18__lane6_strm1_cntl          ( std__pe18__lane6_strm1_cntl       ),      
               .std__pe18__lane6_strm1_data          ( std__pe18__lane6_strm1_data       ),      
               .std__pe18__lane6_strm1_data_valid    ( std__pe18__lane6_strm1_data_valid ),      
               .std__pe18__lane6_strm1_data_mask     ( std__pe18__lane6_strm1_data_mask  ),      

               // PE 18, Lane 7                 
               .pe18__std__lane7_strm0_ready         ( pe18__std__lane7_strm0_ready      ),      
               .std__pe18__lane7_strm0_cntl          ( std__pe18__lane7_strm0_cntl       ),      
               .std__pe18__lane7_strm0_data          ( std__pe18__lane7_strm0_data       ),      
               .std__pe18__lane7_strm0_data_valid    ( std__pe18__lane7_strm0_data_valid ),      
               .std__pe18__lane7_strm0_data_mask     ( std__pe18__lane7_strm0_data_mask  ),      

               .pe18__std__lane7_strm1_ready         ( pe18__std__lane7_strm1_ready      ),      
               .std__pe18__lane7_strm1_cntl          ( std__pe18__lane7_strm1_cntl       ),      
               .std__pe18__lane7_strm1_data          ( std__pe18__lane7_strm1_data       ),      
               .std__pe18__lane7_strm1_data_valid    ( std__pe18__lane7_strm1_data_valid ),      
               .std__pe18__lane7_strm1_data_mask     ( std__pe18__lane7_strm1_data_mask  ),      

               // PE 18, Lane 8                 
               .pe18__std__lane8_strm0_ready         ( pe18__std__lane8_strm0_ready      ),      
               .std__pe18__lane8_strm0_cntl          ( std__pe18__lane8_strm0_cntl       ),      
               .std__pe18__lane8_strm0_data          ( std__pe18__lane8_strm0_data       ),      
               .std__pe18__lane8_strm0_data_valid    ( std__pe18__lane8_strm0_data_valid ),      
               .std__pe18__lane8_strm0_data_mask     ( std__pe18__lane8_strm0_data_mask  ),      

               .pe18__std__lane8_strm1_ready         ( pe18__std__lane8_strm1_ready      ),      
               .std__pe18__lane8_strm1_cntl          ( std__pe18__lane8_strm1_cntl       ),      
               .std__pe18__lane8_strm1_data          ( std__pe18__lane8_strm1_data       ),      
               .std__pe18__lane8_strm1_data_valid    ( std__pe18__lane8_strm1_data_valid ),      
               .std__pe18__lane8_strm1_data_mask     ( std__pe18__lane8_strm1_data_mask  ),      

               // PE 18, Lane 9                 
               .pe18__std__lane9_strm0_ready         ( pe18__std__lane9_strm0_ready      ),      
               .std__pe18__lane9_strm0_cntl          ( std__pe18__lane9_strm0_cntl       ),      
               .std__pe18__lane9_strm0_data          ( std__pe18__lane9_strm0_data       ),      
               .std__pe18__lane9_strm0_data_valid    ( std__pe18__lane9_strm0_data_valid ),      
               .std__pe18__lane9_strm0_data_mask     ( std__pe18__lane9_strm0_data_mask  ),      

               .pe18__std__lane9_strm1_ready         ( pe18__std__lane9_strm1_ready      ),      
               .std__pe18__lane9_strm1_cntl          ( std__pe18__lane9_strm1_cntl       ),      
               .std__pe18__lane9_strm1_data          ( std__pe18__lane9_strm1_data       ),      
               .std__pe18__lane9_strm1_data_valid    ( std__pe18__lane9_strm1_data_valid ),      
               .std__pe18__lane9_strm1_data_mask     ( std__pe18__lane9_strm1_data_mask  ),      

               // PE 18, Lane 10                 
               .pe18__std__lane10_strm0_ready         ( pe18__std__lane10_strm0_ready      ),      
               .std__pe18__lane10_strm0_cntl          ( std__pe18__lane10_strm0_cntl       ),      
               .std__pe18__lane10_strm0_data          ( std__pe18__lane10_strm0_data       ),      
               .std__pe18__lane10_strm0_data_valid    ( std__pe18__lane10_strm0_data_valid ),      
               .std__pe18__lane10_strm0_data_mask     ( std__pe18__lane10_strm0_data_mask  ),      

               .pe18__std__lane10_strm1_ready         ( pe18__std__lane10_strm1_ready      ),      
               .std__pe18__lane10_strm1_cntl          ( std__pe18__lane10_strm1_cntl       ),      
               .std__pe18__lane10_strm1_data          ( std__pe18__lane10_strm1_data       ),      
               .std__pe18__lane10_strm1_data_valid    ( std__pe18__lane10_strm1_data_valid ),      
               .std__pe18__lane10_strm1_data_mask     ( std__pe18__lane10_strm1_data_mask  ),      

               // PE 18, Lane 11                 
               .pe18__std__lane11_strm0_ready         ( pe18__std__lane11_strm0_ready      ),      
               .std__pe18__lane11_strm0_cntl          ( std__pe18__lane11_strm0_cntl       ),      
               .std__pe18__lane11_strm0_data          ( std__pe18__lane11_strm0_data       ),      
               .std__pe18__lane11_strm0_data_valid    ( std__pe18__lane11_strm0_data_valid ),      
               .std__pe18__lane11_strm0_data_mask     ( std__pe18__lane11_strm0_data_mask  ),      

               .pe18__std__lane11_strm1_ready         ( pe18__std__lane11_strm1_ready      ),      
               .std__pe18__lane11_strm1_cntl          ( std__pe18__lane11_strm1_cntl       ),      
               .std__pe18__lane11_strm1_data          ( std__pe18__lane11_strm1_data       ),      
               .std__pe18__lane11_strm1_data_valid    ( std__pe18__lane11_strm1_data_valid ),      
               .std__pe18__lane11_strm1_data_mask     ( std__pe18__lane11_strm1_data_mask  ),      

               // PE 18, Lane 12                 
               .pe18__std__lane12_strm0_ready         ( pe18__std__lane12_strm0_ready      ),      
               .std__pe18__lane12_strm0_cntl          ( std__pe18__lane12_strm0_cntl       ),      
               .std__pe18__lane12_strm0_data          ( std__pe18__lane12_strm0_data       ),      
               .std__pe18__lane12_strm0_data_valid    ( std__pe18__lane12_strm0_data_valid ),      
               .std__pe18__lane12_strm0_data_mask     ( std__pe18__lane12_strm0_data_mask  ),      

               .pe18__std__lane12_strm1_ready         ( pe18__std__lane12_strm1_ready      ),      
               .std__pe18__lane12_strm1_cntl          ( std__pe18__lane12_strm1_cntl       ),      
               .std__pe18__lane12_strm1_data          ( std__pe18__lane12_strm1_data       ),      
               .std__pe18__lane12_strm1_data_valid    ( std__pe18__lane12_strm1_data_valid ),      
               .std__pe18__lane12_strm1_data_mask     ( std__pe18__lane12_strm1_data_mask  ),      

               // PE 18, Lane 13                 
               .pe18__std__lane13_strm0_ready         ( pe18__std__lane13_strm0_ready      ),      
               .std__pe18__lane13_strm0_cntl          ( std__pe18__lane13_strm0_cntl       ),      
               .std__pe18__lane13_strm0_data          ( std__pe18__lane13_strm0_data       ),      
               .std__pe18__lane13_strm0_data_valid    ( std__pe18__lane13_strm0_data_valid ),      
               .std__pe18__lane13_strm0_data_mask     ( std__pe18__lane13_strm0_data_mask  ),      

               .pe18__std__lane13_strm1_ready         ( pe18__std__lane13_strm1_ready      ),      
               .std__pe18__lane13_strm1_cntl          ( std__pe18__lane13_strm1_cntl       ),      
               .std__pe18__lane13_strm1_data          ( std__pe18__lane13_strm1_data       ),      
               .std__pe18__lane13_strm1_data_valid    ( std__pe18__lane13_strm1_data_valid ),      
               .std__pe18__lane13_strm1_data_mask     ( std__pe18__lane13_strm1_data_mask  ),      

               // PE 18, Lane 14                 
               .pe18__std__lane14_strm0_ready         ( pe18__std__lane14_strm0_ready      ),      
               .std__pe18__lane14_strm0_cntl          ( std__pe18__lane14_strm0_cntl       ),      
               .std__pe18__lane14_strm0_data          ( std__pe18__lane14_strm0_data       ),      
               .std__pe18__lane14_strm0_data_valid    ( std__pe18__lane14_strm0_data_valid ),      
               .std__pe18__lane14_strm0_data_mask     ( std__pe18__lane14_strm0_data_mask  ),      

               .pe18__std__lane14_strm1_ready         ( pe18__std__lane14_strm1_ready      ),      
               .std__pe18__lane14_strm1_cntl          ( std__pe18__lane14_strm1_cntl       ),      
               .std__pe18__lane14_strm1_data          ( std__pe18__lane14_strm1_data       ),      
               .std__pe18__lane14_strm1_data_valid    ( std__pe18__lane14_strm1_data_valid ),      
               .std__pe18__lane14_strm1_data_mask     ( std__pe18__lane14_strm1_data_mask  ),      

               // PE 18, Lane 15                 
               .pe18__std__lane15_strm0_ready         ( pe18__std__lane15_strm0_ready      ),      
               .std__pe18__lane15_strm0_cntl          ( std__pe18__lane15_strm0_cntl       ),      
               .std__pe18__lane15_strm0_data          ( std__pe18__lane15_strm0_data       ),      
               .std__pe18__lane15_strm0_data_valid    ( std__pe18__lane15_strm0_data_valid ),      
               .std__pe18__lane15_strm0_data_mask     ( std__pe18__lane15_strm0_data_mask  ),      

               .pe18__std__lane15_strm1_ready         ( pe18__std__lane15_strm1_ready      ),      
               .std__pe18__lane15_strm1_cntl          ( std__pe18__lane15_strm1_cntl       ),      
               .std__pe18__lane15_strm1_data          ( std__pe18__lane15_strm1_data       ),      
               .std__pe18__lane15_strm1_data_valid    ( std__pe18__lane15_strm1_data_valid ),      
               .std__pe18__lane15_strm1_data_mask     ( std__pe18__lane15_strm1_data_mask  ),      

               // PE 18, Lane 16                 
               .pe18__std__lane16_strm0_ready         ( pe18__std__lane16_strm0_ready      ),      
               .std__pe18__lane16_strm0_cntl          ( std__pe18__lane16_strm0_cntl       ),      
               .std__pe18__lane16_strm0_data          ( std__pe18__lane16_strm0_data       ),      
               .std__pe18__lane16_strm0_data_valid    ( std__pe18__lane16_strm0_data_valid ),      
               .std__pe18__lane16_strm0_data_mask     ( std__pe18__lane16_strm0_data_mask  ),      

               .pe18__std__lane16_strm1_ready         ( pe18__std__lane16_strm1_ready      ),      
               .std__pe18__lane16_strm1_cntl          ( std__pe18__lane16_strm1_cntl       ),      
               .std__pe18__lane16_strm1_data          ( std__pe18__lane16_strm1_data       ),      
               .std__pe18__lane16_strm1_data_valid    ( std__pe18__lane16_strm1_data_valid ),      
               .std__pe18__lane16_strm1_data_mask     ( std__pe18__lane16_strm1_data_mask  ),      

               // PE 18, Lane 17                 
               .pe18__std__lane17_strm0_ready         ( pe18__std__lane17_strm0_ready      ),      
               .std__pe18__lane17_strm0_cntl          ( std__pe18__lane17_strm0_cntl       ),      
               .std__pe18__lane17_strm0_data          ( std__pe18__lane17_strm0_data       ),      
               .std__pe18__lane17_strm0_data_valid    ( std__pe18__lane17_strm0_data_valid ),      
               .std__pe18__lane17_strm0_data_mask     ( std__pe18__lane17_strm0_data_mask  ),      

               .pe18__std__lane17_strm1_ready         ( pe18__std__lane17_strm1_ready      ),      
               .std__pe18__lane17_strm1_cntl          ( std__pe18__lane17_strm1_cntl       ),      
               .std__pe18__lane17_strm1_data          ( std__pe18__lane17_strm1_data       ),      
               .std__pe18__lane17_strm1_data_valid    ( std__pe18__lane17_strm1_data_valid ),      
               .std__pe18__lane17_strm1_data_mask     ( std__pe18__lane17_strm1_data_mask  ),      

               // PE 18, Lane 18                 
               .pe18__std__lane18_strm0_ready         ( pe18__std__lane18_strm0_ready      ),      
               .std__pe18__lane18_strm0_cntl          ( std__pe18__lane18_strm0_cntl       ),      
               .std__pe18__lane18_strm0_data          ( std__pe18__lane18_strm0_data       ),      
               .std__pe18__lane18_strm0_data_valid    ( std__pe18__lane18_strm0_data_valid ),      
               .std__pe18__lane18_strm0_data_mask     ( std__pe18__lane18_strm0_data_mask  ),      

               .pe18__std__lane18_strm1_ready         ( pe18__std__lane18_strm1_ready      ),      
               .std__pe18__lane18_strm1_cntl          ( std__pe18__lane18_strm1_cntl       ),      
               .std__pe18__lane18_strm1_data          ( std__pe18__lane18_strm1_data       ),      
               .std__pe18__lane18_strm1_data_valid    ( std__pe18__lane18_strm1_data_valid ),      
               .std__pe18__lane18_strm1_data_mask     ( std__pe18__lane18_strm1_data_mask  ),      

               // PE 18, Lane 19                 
               .pe18__std__lane19_strm0_ready         ( pe18__std__lane19_strm0_ready      ),      
               .std__pe18__lane19_strm0_cntl          ( std__pe18__lane19_strm0_cntl       ),      
               .std__pe18__lane19_strm0_data          ( std__pe18__lane19_strm0_data       ),      
               .std__pe18__lane19_strm0_data_valid    ( std__pe18__lane19_strm0_data_valid ),      
               .std__pe18__lane19_strm0_data_mask     ( std__pe18__lane19_strm0_data_mask  ),      

               .pe18__std__lane19_strm1_ready         ( pe18__std__lane19_strm1_ready      ),      
               .std__pe18__lane19_strm1_cntl          ( std__pe18__lane19_strm1_cntl       ),      
               .std__pe18__lane19_strm1_data          ( std__pe18__lane19_strm1_data       ),      
               .std__pe18__lane19_strm1_data_valid    ( std__pe18__lane19_strm1_data_valid ),      
               .std__pe18__lane19_strm1_data_mask     ( std__pe18__lane19_strm1_data_mask  ),      

               // PE 18, Lane 20                 
               .pe18__std__lane20_strm0_ready         ( pe18__std__lane20_strm0_ready      ),      
               .std__pe18__lane20_strm0_cntl          ( std__pe18__lane20_strm0_cntl       ),      
               .std__pe18__lane20_strm0_data          ( std__pe18__lane20_strm0_data       ),      
               .std__pe18__lane20_strm0_data_valid    ( std__pe18__lane20_strm0_data_valid ),      
               .std__pe18__lane20_strm0_data_mask     ( std__pe18__lane20_strm0_data_mask  ),      

               .pe18__std__lane20_strm1_ready         ( pe18__std__lane20_strm1_ready      ),      
               .std__pe18__lane20_strm1_cntl          ( std__pe18__lane20_strm1_cntl       ),      
               .std__pe18__lane20_strm1_data          ( std__pe18__lane20_strm1_data       ),      
               .std__pe18__lane20_strm1_data_valid    ( std__pe18__lane20_strm1_data_valid ),      
               .std__pe18__lane20_strm1_data_mask     ( std__pe18__lane20_strm1_data_mask  ),      

               // PE 18, Lane 21                 
               .pe18__std__lane21_strm0_ready         ( pe18__std__lane21_strm0_ready      ),      
               .std__pe18__lane21_strm0_cntl          ( std__pe18__lane21_strm0_cntl       ),      
               .std__pe18__lane21_strm0_data          ( std__pe18__lane21_strm0_data       ),      
               .std__pe18__lane21_strm0_data_valid    ( std__pe18__lane21_strm0_data_valid ),      
               .std__pe18__lane21_strm0_data_mask     ( std__pe18__lane21_strm0_data_mask  ),      

               .pe18__std__lane21_strm1_ready         ( pe18__std__lane21_strm1_ready      ),      
               .std__pe18__lane21_strm1_cntl          ( std__pe18__lane21_strm1_cntl       ),      
               .std__pe18__lane21_strm1_data          ( std__pe18__lane21_strm1_data       ),      
               .std__pe18__lane21_strm1_data_valid    ( std__pe18__lane21_strm1_data_valid ),      
               .std__pe18__lane21_strm1_data_mask     ( std__pe18__lane21_strm1_data_mask  ),      

               // PE 18, Lane 22                 
               .pe18__std__lane22_strm0_ready         ( pe18__std__lane22_strm0_ready      ),      
               .std__pe18__lane22_strm0_cntl          ( std__pe18__lane22_strm0_cntl       ),      
               .std__pe18__lane22_strm0_data          ( std__pe18__lane22_strm0_data       ),      
               .std__pe18__lane22_strm0_data_valid    ( std__pe18__lane22_strm0_data_valid ),      
               .std__pe18__lane22_strm0_data_mask     ( std__pe18__lane22_strm0_data_mask  ),      

               .pe18__std__lane22_strm1_ready         ( pe18__std__lane22_strm1_ready      ),      
               .std__pe18__lane22_strm1_cntl          ( std__pe18__lane22_strm1_cntl       ),      
               .std__pe18__lane22_strm1_data          ( std__pe18__lane22_strm1_data       ),      
               .std__pe18__lane22_strm1_data_valid    ( std__pe18__lane22_strm1_data_valid ),      
               .std__pe18__lane22_strm1_data_mask     ( std__pe18__lane22_strm1_data_mask  ),      

               // PE 18, Lane 23                 
               .pe18__std__lane23_strm0_ready         ( pe18__std__lane23_strm0_ready      ),      
               .std__pe18__lane23_strm0_cntl          ( std__pe18__lane23_strm0_cntl       ),      
               .std__pe18__lane23_strm0_data          ( std__pe18__lane23_strm0_data       ),      
               .std__pe18__lane23_strm0_data_valid    ( std__pe18__lane23_strm0_data_valid ),      
               .std__pe18__lane23_strm0_data_mask     ( std__pe18__lane23_strm0_data_mask  ),      

               .pe18__std__lane23_strm1_ready         ( pe18__std__lane23_strm1_ready      ),      
               .std__pe18__lane23_strm1_cntl          ( std__pe18__lane23_strm1_cntl       ),      
               .std__pe18__lane23_strm1_data          ( std__pe18__lane23_strm1_data       ),      
               .std__pe18__lane23_strm1_data_valid    ( std__pe18__lane23_strm1_data_valid ),      
               .std__pe18__lane23_strm1_data_mask     ( std__pe18__lane23_strm1_data_mask  ),      

               // PE 18, Lane 24                 
               .pe18__std__lane24_strm0_ready         ( pe18__std__lane24_strm0_ready      ),      
               .std__pe18__lane24_strm0_cntl          ( std__pe18__lane24_strm0_cntl       ),      
               .std__pe18__lane24_strm0_data          ( std__pe18__lane24_strm0_data       ),      
               .std__pe18__lane24_strm0_data_valid    ( std__pe18__lane24_strm0_data_valid ),      
               .std__pe18__lane24_strm0_data_mask     ( std__pe18__lane24_strm0_data_mask  ),      

               .pe18__std__lane24_strm1_ready         ( pe18__std__lane24_strm1_ready      ),      
               .std__pe18__lane24_strm1_cntl          ( std__pe18__lane24_strm1_cntl       ),      
               .std__pe18__lane24_strm1_data          ( std__pe18__lane24_strm1_data       ),      
               .std__pe18__lane24_strm1_data_valid    ( std__pe18__lane24_strm1_data_valid ),      
               .std__pe18__lane24_strm1_data_mask     ( std__pe18__lane24_strm1_data_mask  ),      

               // PE 18, Lane 25                 
               .pe18__std__lane25_strm0_ready         ( pe18__std__lane25_strm0_ready      ),      
               .std__pe18__lane25_strm0_cntl          ( std__pe18__lane25_strm0_cntl       ),      
               .std__pe18__lane25_strm0_data          ( std__pe18__lane25_strm0_data       ),      
               .std__pe18__lane25_strm0_data_valid    ( std__pe18__lane25_strm0_data_valid ),      
               .std__pe18__lane25_strm0_data_mask     ( std__pe18__lane25_strm0_data_mask  ),      

               .pe18__std__lane25_strm1_ready         ( pe18__std__lane25_strm1_ready      ),      
               .std__pe18__lane25_strm1_cntl          ( std__pe18__lane25_strm1_cntl       ),      
               .std__pe18__lane25_strm1_data          ( std__pe18__lane25_strm1_data       ),      
               .std__pe18__lane25_strm1_data_valid    ( std__pe18__lane25_strm1_data_valid ),      
               .std__pe18__lane25_strm1_data_mask     ( std__pe18__lane25_strm1_data_mask  ),      

               // PE 18, Lane 26                 
               .pe18__std__lane26_strm0_ready         ( pe18__std__lane26_strm0_ready      ),      
               .std__pe18__lane26_strm0_cntl          ( std__pe18__lane26_strm0_cntl       ),      
               .std__pe18__lane26_strm0_data          ( std__pe18__lane26_strm0_data       ),      
               .std__pe18__lane26_strm0_data_valid    ( std__pe18__lane26_strm0_data_valid ),      
               .std__pe18__lane26_strm0_data_mask     ( std__pe18__lane26_strm0_data_mask  ),      

               .pe18__std__lane26_strm1_ready         ( pe18__std__lane26_strm1_ready      ),      
               .std__pe18__lane26_strm1_cntl          ( std__pe18__lane26_strm1_cntl       ),      
               .std__pe18__lane26_strm1_data          ( std__pe18__lane26_strm1_data       ),      
               .std__pe18__lane26_strm1_data_valid    ( std__pe18__lane26_strm1_data_valid ),      
               .std__pe18__lane26_strm1_data_mask     ( std__pe18__lane26_strm1_data_mask  ),      

               // PE 18, Lane 27                 
               .pe18__std__lane27_strm0_ready         ( pe18__std__lane27_strm0_ready      ),      
               .std__pe18__lane27_strm0_cntl          ( std__pe18__lane27_strm0_cntl       ),      
               .std__pe18__lane27_strm0_data          ( std__pe18__lane27_strm0_data       ),      
               .std__pe18__lane27_strm0_data_valid    ( std__pe18__lane27_strm0_data_valid ),      
               .std__pe18__lane27_strm0_data_mask     ( std__pe18__lane27_strm0_data_mask  ),      

               .pe18__std__lane27_strm1_ready         ( pe18__std__lane27_strm1_ready      ),      
               .std__pe18__lane27_strm1_cntl          ( std__pe18__lane27_strm1_cntl       ),      
               .std__pe18__lane27_strm1_data          ( std__pe18__lane27_strm1_data       ),      
               .std__pe18__lane27_strm1_data_valid    ( std__pe18__lane27_strm1_data_valid ),      
               .std__pe18__lane27_strm1_data_mask     ( std__pe18__lane27_strm1_data_mask  ),      

               // PE 18, Lane 28                 
               .pe18__std__lane28_strm0_ready         ( pe18__std__lane28_strm0_ready      ),      
               .std__pe18__lane28_strm0_cntl          ( std__pe18__lane28_strm0_cntl       ),      
               .std__pe18__lane28_strm0_data          ( std__pe18__lane28_strm0_data       ),      
               .std__pe18__lane28_strm0_data_valid    ( std__pe18__lane28_strm0_data_valid ),      
               .std__pe18__lane28_strm0_data_mask     ( std__pe18__lane28_strm0_data_mask  ),      

               .pe18__std__lane28_strm1_ready         ( pe18__std__lane28_strm1_ready      ),      
               .std__pe18__lane28_strm1_cntl          ( std__pe18__lane28_strm1_cntl       ),      
               .std__pe18__lane28_strm1_data          ( std__pe18__lane28_strm1_data       ),      
               .std__pe18__lane28_strm1_data_valid    ( std__pe18__lane28_strm1_data_valid ),      
               .std__pe18__lane28_strm1_data_mask     ( std__pe18__lane28_strm1_data_mask  ),      

               // PE 18, Lane 29                 
               .pe18__std__lane29_strm0_ready         ( pe18__std__lane29_strm0_ready      ),      
               .std__pe18__lane29_strm0_cntl          ( std__pe18__lane29_strm0_cntl       ),      
               .std__pe18__lane29_strm0_data          ( std__pe18__lane29_strm0_data       ),      
               .std__pe18__lane29_strm0_data_valid    ( std__pe18__lane29_strm0_data_valid ),      
               .std__pe18__lane29_strm0_data_mask     ( std__pe18__lane29_strm0_data_mask  ),      

               .pe18__std__lane29_strm1_ready         ( pe18__std__lane29_strm1_ready      ),      
               .std__pe18__lane29_strm1_cntl          ( std__pe18__lane29_strm1_cntl       ),      
               .std__pe18__lane29_strm1_data          ( std__pe18__lane29_strm1_data       ),      
               .std__pe18__lane29_strm1_data_valid    ( std__pe18__lane29_strm1_data_valid ),      
               .std__pe18__lane29_strm1_data_mask     ( std__pe18__lane29_strm1_data_mask  ),      

               // PE 18, Lane 30                 
               .pe18__std__lane30_strm0_ready         ( pe18__std__lane30_strm0_ready      ),      
               .std__pe18__lane30_strm0_cntl          ( std__pe18__lane30_strm0_cntl       ),      
               .std__pe18__lane30_strm0_data          ( std__pe18__lane30_strm0_data       ),      
               .std__pe18__lane30_strm0_data_valid    ( std__pe18__lane30_strm0_data_valid ),      
               .std__pe18__lane30_strm0_data_mask     ( std__pe18__lane30_strm0_data_mask  ),      

               .pe18__std__lane30_strm1_ready         ( pe18__std__lane30_strm1_ready      ),      
               .std__pe18__lane30_strm1_cntl          ( std__pe18__lane30_strm1_cntl       ),      
               .std__pe18__lane30_strm1_data          ( std__pe18__lane30_strm1_data       ),      
               .std__pe18__lane30_strm1_data_valid    ( std__pe18__lane30_strm1_data_valid ),      
               .std__pe18__lane30_strm1_data_mask     ( std__pe18__lane30_strm1_data_mask  ),      

               // PE 18, Lane 31                 
               .pe18__std__lane31_strm0_ready         ( pe18__std__lane31_strm0_ready      ),      
               .std__pe18__lane31_strm0_cntl          ( std__pe18__lane31_strm0_cntl       ),      
               .std__pe18__lane31_strm0_data          ( std__pe18__lane31_strm0_data       ),      
               .std__pe18__lane31_strm0_data_valid    ( std__pe18__lane31_strm0_data_valid ),      
               .std__pe18__lane31_strm0_data_mask     ( std__pe18__lane31_strm0_data_mask  ),      

               .pe18__std__lane31_strm1_ready         ( pe18__std__lane31_strm1_ready      ),      
               .std__pe18__lane31_strm1_cntl          ( std__pe18__lane31_strm1_cntl       ),      
               .std__pe18__lane31_strm1_data          ( std__pe18__lane31_strm1_data       ),      
               .std__pe18__lane31_strm1_data_valid    ( std__pe18__lane31_strm1_data_valid ),      
               .std__pe18__lane31_strm1_data_mask     ( std__pe18__lane31_strm1_data_mask  ),      

               // PE 19, Lane 0                 
               .pe19__std__lane0_strm0_ready         ( pe19__std__lane0_strm0_ready      ),      
               .std__pe19__lane0_strm0_cntl          ( std__pe19__lane0_strm0_cntl       ),      
               .std__pe19__lane0_strm0_data          ( std__pe19__lane0_strm0_data       ),      
               .std__pe19__lane0_strm0_data_valid    ( std__pe19__lane0_strm0_data_valid ),      
               .std__pe19__lane0_strm0_data_mask     ( std__pe19__lane0_strm0_data_mask  ),      

               .pe19__std__lane0_strm1_ready         ( pe19__std__lane0_strm1_ready      ),      
               .std__pe19__lane0_strm1_cntl          ( std__pe19__lane0_strm1_cntl       ),      
               .std__pe19__lane0_strm1_data          ( std__pe19__lane0_strm1_data       ),      
               .std__pe19__lane0_strm1_data_valid    ( std__pe19__lane0_strm1_data_valid ),      
               .std__pe19__lane0_strm1_data_mask     ( std__pe19__lane0_strm1_data_mask  ),      

               // PE 19, Lane 1                 
               .pe19__std__lane1_strm0_ready         ( pe19__std__lane1_strm0_ready      ),      
               .std__pe19__lane1_strm0_cntl          ( std__pe19__lane1_strm0_cntl       ),      
               .std__pe19__lane1_strm0_data          ( std__pe19__lane1_strm0_data       ),      
               .std__pe19__lane1_strm0_data_valid    ( std__pe19__lane1_strm0_data_valid ),      
               .std__pe19__lane1_strm0_data_mask     ( std__pe19__lane1_strm0_data_mask  ),      

               .pe19__std__lane1_strm1_ready         ( pe19__std__lane1_strm1_ready      ),      
               .std__pe19__lane1_strm1_cntl          ( std__pe19__lane1_strm1_cntl       ),      
               .std__pe19__lane1_strm1_data          ( std__pe19__lane1_strm1_data       ),      
               .std__pe19__lane1_strm1_data_valid    ( std__pe19__lane1_strm1_data_valid ),      
               .std__pe19__lane1_strm1_data_mask     ( std__pe19__lane1_strm1_data_mask  ),      

               // PE 19, Lane 2                 
               .pe19__std__lane2_strm0_ready         ( pe19__std__lane2_strm0_ready      ),      
               .std__pe19__lane2_strm0_cntl          ( std__pe19__lane2_strm0_cntl       ),      
               .std__pe19__lane2_strm0_data          ( std__pe19__lane2_strm0_data       ),      
               .std__pe19__lane2_strm0_data_valid    ( std__pe19__lane2_strm0_data_valid ),      
               .std__pe19__lane2_strm0_data_mask     ( std__pe19__lane2_strm0_data_mask  ),      

               .pe19__std__lane2_strm1_ready         ( pe19__std__lane2_strm1_ready      ),      
               .std__pe19__lane2_strm1_cntl          ( std__pe19__lane2_strm1_cntl       ),      
               .std__pe19__lane2_strm1_data          ( std__pe19__lane2_strm1_data       ),      
               .std__pe19__lane2_strm1_data_valid    ( std__pe19__lane2_strm1_data_valid ),      
               .std__pe19__lane2_strm1_data_mask     ( std__pe19__lane2_strm1_data_mask  ),      

               // PE 19, Lane 3                 
               .pe19__std__lane3_strm0_ready         ( pe19__std__lane3_strm0_ready      ),      
               .std__pe19__lane3_strm0_cntl          ( std__pe19__lane3_strm0_cntl       ),      
               .std__pe19__lane3_strm0_data          ( std__pe19__lane3_strm0_data       ),      
               .std__pe19__lane3_strm0_data_valid    ( std__pe19__lane3_strm0_data_valid ),      
               .std__pe19__lane3_strm0_data_mask     ( std__pe19__lane3_strm0_data_mask  ),      

               .pe19__std__lane3_strm1_ready         ( pe19__std__lane3_strm1_ready      ),      
               .std__pe19__lane3_strm1_cntl          ( std__pe19__lane3_strm1_cntl       ),      
               .std__pe19__lane3_strm1_data          ( std__pe19__lane3_strm1_data       ),      
               .std__pe19__lane3_strm1_data_valid    ( std__pe19__lane3_strm1_data_valid ),      
               .std__pe19__lane3_strm1_data_mask     ( std__pe19__lane3_strm1_data_mask  ),      

               // PE 19, Lane 4                 
               .pe19__std__lane4_strm0_ready         ( pe19__std__lane4_strm0_ready      ),      
               .std__pe19__lane4_strm0_cntl          ( std__pe19__lane4_strm0_cntl       ),      
               .std__pe19__lane4_strm0_data          ( std__pe19__lane4_strm0_data       ),      
               .std__pe19__lane4_strm0_data_valid    ( std__pe19__lane4_strm0_data_valid ),      
               .std__pe19__lane4_strm0_data_mask     ( std__pe19__lane4_strm0_data_mask  ),      

               .pe19__std__lane4_strm1_ready         ( pe19__std__lane4_strm1_ready      ),      
               .std__pe19__lane4_strm1_cntl          ( std__pe19__lane4_strm1_cntl       ),      
               .std__pe19__lane4_strm1_data          ( std__pe19__lane4_strm1_data       ),      
               .std__pe19__lane4_strm1_data_valid    ( std__pe19__lane4_strm1_data_valid ),      
               .std__pe19__lane4_strm1_data_mask     ( std__pe19__lane4_strm1_data_mask  ),      

               // PE 19, Lane 5                 
               .pe19__std__lane5_strm0_ready         ( pe19__std__lane5_strm0_ready      ),      
               .std__pe19__lane5_strm0_cntl          ( std__pe19__lane5_strm0_cntl       ),      
               .std__pe19__lane5_strm0_data          ( std__pe19__lane5_strm0_data       ),      
               .std__pe19__lane5_strm0_data_valid    ( std__pe19__lane5_strm0_data_valid ),      
               .std__pe19__lane5_strm0_data_mask     ( std__pe19__lane5_strm0_data_mask  ),      

               .pe19__std__lane5_strm1_ready         ( pe19__std__lane5_strm1_ready      ),      
               .std__pe19__lane5_strm1_cntl          ( std__pe19__lane5_strm1_cntl       ),      
               .std__pe19__lane5_strm1_data          ( std__pe19__lane5_strm1_data       ),      
               .std__pe19__lane5_strm1_data_valid    ( std__pe19__lane5_strm1_data_valid ),      
               .std__pe19__lane5_strm1_data_mask     ( std__pe19__lane5_strm1_data_mask  ),      

               // PE 19, Lane 6                 
               .pe19__std__lane6_strm0_ready         ( pe19__std__lane6_strm0_ready      ),      
               .std__pe19__lane6_strm0_cntl          ( std__pe19__lane6_strm0_cntl       ),      
               .std__pe19__lane6_strm0_data          ( std__pe19__lane6_strm0_data       ),      
               .std__pe19__lane6_strm0_data_valid    ( std__pe19__lane6_strm0_data_valid ),      
               .std__pe19__lane6_strm0_data_mask     ( std__pe19__lane6_strm0_data_mask  ),      

               .pe19__std__lane6_strm1_ready         ( pe19__std__lane6_strm1_ready      ),      
               .std__pe19__lane6_strm1_cntl          ( std__pe19__lane6_strm1_cntl       ),      
               .std__pe19__lane6_strm1_data          ( std__pe19__lane6_strm1_data       ),      
               .std__pe19__lane6_strm1_data_valid    ( std__pe19__lane6_strm1_data_valid ),      
               .std__pe19__lane6_strm1_data_mask     ( std__pe19__lane6_strm1_data_mask  ),      

               // PE 19, Lane 7                 
               .pe19__std__lane7_strm0_ready         ( pe19__std__lane7_strm0_ready      ),      
               .std__pe19__lane7_strm0_cntl          ( std__pe19__lane7_strm0_cntl       ),      
               .std__pe19__lane7_strm0_data          ( std__pe19__lane7_strm0_data       ),      
               .std__pe19__lane7_strm0_data_valid    ( std__pe19__lane7_strm0_data_valid ),      
               .std__pe19__lane7_strm0_data_mask     ( std__pe19__lane7_strm0_data_mask  ),      

               .pe19__std__lane7_strm1_ready         ( pe19__std__lane7_strm1_ready      ),      
               .std__pe19__lane7_strm1_cntl          ( std__pe19__lane7_strm1_cntl       ),      
               .std__pe19__lane7_strm1_data          ( std__pe19__lane7_strm1_data       ),      
               .std__pe19__lane7_strm1_data_valid    ( std__pe19__lane7_strm1_data_valid ),      
               .std__pe19__lane7_strm1_data_mask     ( std__pe19__lane7_strm1_data_mask  ),      

               // PE 19, Lane 8                 
               .pe19__std__lane8_strm0_ready         ( pe19__std__lane8_strm0_ready      ),      
               .std__pe19__lane8_strm0_cntl          ( std__pe19__lane8_strm0_cntl       ),      
               .std__pe19__lane8_strm0_data          ( std__pe19__lane8_strm0_data       ),      
               .std__pe19__lane8_strm0_data_valid    ( std__pe19__lane8_strm0_data_valid ),      
               .std__pe19__lane8_strm0_data_mask     ( std__pe19__lane8_strm0_data_mask  ),      

               .pe19__std__lane8_strm1_ready         ( pe19__std__lane8_strm1_ready      ),      
               .std__pe19__lane8_strm1_cntl          ( std__pe19__lane8_strm1_cntl       ),      
               .std__pe19__lane8_strm1_data          ( std__pe19__lane8_strm1_data       ),      
               .std__pe19__lane8_strm1_data_valid    ( std__pe19__lane8_strm1_data_valid ),      
               .std__pe19__lane8_strm1_data_mask     ( std__pe19__lane8_strm1_data_mask  ),      

               // PE 19, Lane 9                 
               .pe19__std__lane9_strm0_ready         ( pe19__std__lane9_strm0_ready      ),      
               .std__pe19__lane9_strm0_cntl          ( std__pe19__lane9_strm0_cntl       ),      
               .std__pe19__lane9_strm0_data          ( std__pe19__lane9_strm0_data       ),      
               .std__pe19__lane9_strm0_data_valid    ( std__pe19__lane9_strm0_data_valid ),      
               .std__pe19__lane9_strm0_data_mask     ( std__pe19__lane9_strm0_data_mask  ),      

               .pe19__std__lane9_strm1_ready         ( pe19__std__lane9_strm1_ready      ),      
               .std__pe19__lane9_strm1_cntl          ( std__pe19__lane9_strm1_cntl       ),      
               .std__pe19__lane9_strm1_data          ( std__pe19__lane9_strm1_data       ),      
               .std__pe19__lane9_strm1_data_valid    ( std__pe19__lane9_strm1_data_valid ),      
               .std__pe19__lane9_strm1_data_mask     ( std__pe19__lane9_strm1_data_mask  ),      

               // PE 19, Lane 10                 
               .pe19__std__lane10_strm0_ready         ( pe19__std__lane10_strm0_ready      ),      
               .std__pe19__lane10_strm0_cntl          ( std__pe19__lane10_strm0_cntl       ),      
               .std__pe19__lane10_strm0_data          ( std__pe19__lane10_strm0_data       ),      
               .std__pe19__lane10_strm0_data_valid    ( std__pe19__lane10_strm0_data_valid ),      
               .std__pe19__lane10_strm0_data_mask     ( std__pe19__lane10_strm0_data_mask  ),      

               .pe19__std__lane10_strm1_ready         ( pe19__std__lane10_strm1_ready      ),      
               .std__pe19__lane10_strm1_cntl          ( std__pe19__lane10_strm1_cntl       ),      
               .std__pe19__lane10_strm1_data          ( std__pe19__lane10_strm1_data       ),      
               .std__pe19__lane10_strm1_data_valid    ( std__pe19__lane10_strm1_data_valid ),      
               .std__pe19__lane10_strm1_data_mask     ( std__pe19__lane10_strm1_data_mask  ),      

               // PE 19, Lane 11                 
               .pe19__std__lane11_strm0_ready         ( pe19__std__lane11_strm0_ready      ),      
               .std__pe19__lane11_strm0_cntl          ( std__pe19__lane11_strm0_cntl       ),      
               .std__pe19__lane11_strm0_data          ( std__pe19__lane11_strm0_data       ),      
               .std__pe19__lane11_strm0_data_valid    ( std__pe19__lane11_strm0_data_valid ),      
               .std__pe19__lane11_strm0_data_mask     ( std__pe19__lane11_strm0_data_mask  ),      

               .pe19__std__lane11_strm1_ready         ( pe19__std__lane11_strm1_ready      ),      
               .std__pe19__lane11_strm1_cntl          ( std__pe19__lane11_strm1_cntl       ),      
               .std__pe19__lane11_strm1_data          ( std__pe19__lane11_strm1_data       ),      
               .std__pe19__lane11_strm1_data_valid    ( std__pe19__lane11_strm1_data_valid ),      
               .std__pe19__lane11_strm1_data_mask     ( std__pe19__lane11_strm1_data_mask  ),      

               // PE 19, Lane 12                 
               .pe19__std__lane12_strm0_ready         ( pe19__std__lane12_strm0_ready      ),      
               .std__pe19__lane12_strm0_cntl          ( std__pe19__lane12_strm0_cntl       ),      
               .std__pe19__lane12_strm0_data          ( std__pe19__lane12_strm0_data       ),      
               .std__pe19__lane12_strm0_data_valid    ( std__pe19__lane12_strm0_data_valid ),      
               .std__pe19__lane12_strm0_data_mask     ( std__pe19__lane12_strm0_data_mask  ),      

               .pe19__std__lane12_strm1_ready         ( pe19__std__lane12_strm1_ready      ),      
               .std__pe19__lane12_strm1_cntl          ( std__pe19__lane12_strm1_cntl       ),      
               .std__pe19__lane12_strm1_data          ( std__pe19__lane12_strm1_data       ),      
               .std__pe19__lane12_strm1_data_valid    ( std__pe19__lane12_strm1_data_valid ),      
               .std__pe19__lane12_strm1_data_mask     ( std__pe19__lane12_strm1_data_mask  ),      

               // PE 19, Lane 13                 
               .pe19__std__lane13_strm0_ready         ( pe19__std__lane13_strm0_ready      ),      
               .std__pe19__lane13_strm0_cntl          ( std__pe19__lane13_strm0_cntl       ),      
               .std__pe19__lane13_strm0_data          ( std__pe19__lane13_strm0_data       ),      
               .std__pe19__lane13_strm0_data_valid    ( std__pe19__lane13_strm0_data_valid ),      
               .std__pe19__lane13_strm0_data_mask     ( std__pe19__lane13_strm0_data_mask  ),      

               .pe19__std__lane13_strm1_ready         ( pe19__std__lane13_strm1_ready      ),      
               .std__pe19__lane13_strm1_cntl          ( std__pe19__lane13_strm1_cntl       ),      
               .std__pe19__lane13_strm1_data          ( std__pe19__lane13_strm1_data       ),      
               .std__pe19__lane13_strm1_data_valid    ( std__pe19__lane13_strm1_data_valid ),      
               .std__pe19__lane13_strm1_data_mask     ( std__pe19__lane13_strm1_data_mask  ),      

               // PE 19, Lane 14                 
               .pe19__std__lane14_strm0_ready         ( pe19__std__lane14_strm0_ready      ),      
               .std__pe19__lane14_strm0_cntl          ( std__pe19__lane14_strm0_cntl       ),      
               .std__pe19__lane14_strm0_data          ( std__pe19__lane14_strm0_data       ),      
               .std__pe19__lane14_strm0_data_valid    ( std__pe19__lane14_strm0_data_valid ),      
               .std__pe19__lane14_strm0_data_mask     ( std__pe19__lane14_strm0_data_mask  ),      

               .pe19__std__lane14_strm1_ready         ( pe19__std__lane14_strm1_ready      ),      
               .std__pe19__lane14_strm1_cntl          ( std__pe19__lane14_strm1_cntl       ),      
               .std__pe19__lane14_strm1_data          ( std__pe19__lane14_strm1_data       ),      
               .std__pe19__lane14_strm1_data_valid    ( std__pe19__lane14_strm1_data_valid ),      
               .std__pe19__lane14_strm1_data_mask     ( std__pe19__lane14_strm1_data_mask  ),      

               // PE 19, Lane 15                 
               .pe19__std__lane15_strm0_ready         ( pe19__std__lane15_strm0_ready      ),      
               .std__pe19__lane15_strm0_cntl          ( std__pe19__lane15_strm0_cntl       ),      
               .std__pe19__lane15_strm0_data          ( std__pe19__lane15_strm0_data       ),      
               .std__pe19__lane15_strm0_data_valid    ( std__pe19__lane15_strm0_data_valid ),      
               .std__pe19__lane15_strm0_data_mask     ( std__pe19__lane15_strm0_data_mask  ),      

               .pe19__std__lane15_strm1_ready         ( pe19__std__lane15_strm1_ready      ),      
               .std__pe19__lane15_strm1_cntl          ( std__pe19__lane15_strm1_cntl       ),      
               .std__pe19__lane15_strm1_data          ( std__pe19__lane15_strm1_data       ),      
               .std__pe19__lane15_strm1_data_valid    ( std__pe19__lane15_strm1_data_valid ),      
               .std__pe19__lane15_strm1_data_mask     ( std__pe19__lane15_strm1_data_mask  ),      

               // PE 19, Lane 16                 
               .pe19__std__lane16_strm0_ready         ( pe19__std__lane16_strm0_ready      ),      
               .std__pe19__lane16_strm0_cntl          ( std__pe19__lane16_strm0_cntl       ),      
               .std__pe19__lane16_strm0_data          ( std__pe19__lane16_strm0_data       ),      
               .std__pe19__lane16_strm0_data_valid    ( std__pe19__lane16_strm0_data_valid ),      
               .std__pe19__lane16_strm0_data_mask     ( std__pe19__lane16_strm0_data_mask  ),      

               .pe19__std__lane16_strm1_ready         ( pe19__std__lane16_strm1_ready      ),      
               .std__pe19__lane16_strm1_cntl          ( std__pe19__lane16_strm1_cntl       ),      
               .std__pe19__lane16_strm1_data          ( std__pe19__lane16_strm1_data       ),      
               .std__pe19__lane16_strm1_data_valid    ( std__pe19__lane16_strm1_data_valid ),      
               .std__pe19__lane16_strm1_data_mask     ( std__pe19__lane16_strm1_data_mask  ),      

               // PE 19, Lane 17                 
               .pe19__std__lane17_strm0_ready         ( pe19__std__lane17_strm0_ready      ),      
               .std__pe19__lane17_strm0_cntl          ( std__pe19__lane17_strm0_cntl       ),      
               .std__pe19__lane17_strm0_data          ( std__pe19__lane17_strm0_data       ),      
               .std__pe19__lane17_strm0_data_valid    ( std__pe19__lane17_strm0_data_valid ),      
               .std__pe19__lane17_strm0_data_mask     ( std__pe19__lane17_strm0_data_mask  ),      

               .pe19__std__lane17_strm1_ready         ( pe19__std__lane17_strm1_ready      ),      
               .std__pe19__lane17_strm1_cntl          ( std__pe19__lane17_strm1_cntl       ),      
               .std__pe19__lane17_strm1_data          ( std__pe19__lane17_strm1_data       ),      
               .std__pe19__lane17_strm1_data_valid    ( std__pe19__lane17_strm1_data_valid ),      
               .std__pe19__lane17_strm1_data_mask     ( std__pe19__lane17_strm1_data_mask  ),      

               // PE 19, Lane 18                 
               .pe19__std__lane18_strm0_ready         ( pe19__std__lane18_strm0_ready      ),      
               .std__pe19__lane18_strm0_cntl          ( std__pe19__lane18_strm0_cntl       ),      
               .std__pe19__lane18_strm0_data          ( std__pe19__lane18_strm0_data       ),      
               .std__pe19__lane18_strm0_data_valid    ( std__pe19__lane18_strm0_data_valid ),      
               .std__pe19__lane18_strm0_data_mask     ( std__pe19__lane18_strm0_data_mask  ),      

               .pe19__std__lane18_strm1_ready         ( pe19__std__lane18_strm1_ready      ),      
               .std__pe19__lane18_strm1_cntl          ( std__pe19__lane18_strm1_cntl       ),      
               .std__pe19__lane18_strm1_data          ( std__pe19__lane18_strm1_data       ),      
               .std__pe19__lane18_strm1_data_valid    ( std__pe19__lane18_strm1_data_valid ),      
               .std__pe19__lane18_strm1_data_mask     ( std__pe19__lane18_strm1_data_mask  ),      

               // PE 19, Lane 19                 
               .pe19__std__lane19_strm0_ready         ( pe19__std__lane19_strm0_ready      ),      
               .std__pe19__lane19_strm0_cntl          ( std__pe19__lane19_strm0_cntl       ),      
               .std__pe19__lane19_strm0_data          ( std__pe19__lane19_strm0_data       ),      
               .std__pe19__lane19_strm0_data_valid    ( std__pe19__lane19_strm0_data_valid ),      
               .std__pe19__lane19_strm0_data_mask     ( std__pe19__lane19_strm0_data_mask  ),      

               .pe19__std__lane19_strm1_ready         ( pe19__std__lane19_strm1_ready      ),      
               .std__pe19__lane19_strm1_cntl          ( std__pe19__lane19_strm1_cntl       ),      
               .std__pe19__lane19_strm1_data          ( std__pe19__lane19_strm1_data       ),      
               .std__pe19__lane19_strm1_data_valid    ( std__pe19__lane19_strm1_data_valid ),      
               .std__pe19__lane19_strm1_data_mask     ( std__pe19__lane19_strm1_data_mask  ),      

               // PE 19, Lane 20                 
               .pe19__std__lane20_strm0_ready         ( pe19__std__lane20_strm0_ready      ),      
               .std__pe19__lane20_strm0_cntl          ( std__pe19__lane20_strm0_cntl       ),      
               .std__pe19__lane20_strm0_data          ( std__pe19__lane20_strm0_data       ),      
               .std__pe19__lane20_strm0_data_valid    ( std__pe19__lane20_strm0_data_valid ),      
               .std__pe19__lane20_strm0_data_mask     ( std__pe19__lane20_strm0_data_mask  ),      

               .pe19__std__lane20_strm1_ready         ( pe19__std__lane20_strm1_ready      ),      
               .std__pe19__lane20_strm1_cntl          ( std__pe19__lane20_strm1_cntl       ),      
               .std__pe19__lane20_strm1_data          ( std__pe19__lane20_strm1_data       ),      
               .std__pe19__lane20_strm1_data_valid    ( std__pe19__lane20_strm1_data_valid ),      
               .std__pe19__lane20_strm1_data_mask     ( std__pe19__lane20_strm1_data_mask  ),      

               // PE 19, Lane 21                 
               .pe19__std__lane21_strm0_ready         ( pe19__std__lane21_strm0_ready      ),      
               .std__pe19__lane21_strm0_cntl          ( std__pe19__lane21_strm0_cntl       ),      
               .std__pe19__lane21_strm0_data          ( std__pe19__lane21_strm0_data       ),      
               .std__pe19__lane21_strm0_data_valid    ( std__pe19__lane21_strm0_data_valid ),      
               .std__pe19__lane21_strm0_data_mask     ( std__pe19__lane21_strm0_data_mask  ),      

               .pe19__std__lane21_strm1_ready         ( pe19__std__lane21_strm1_ready      ),      
               .std__pe19__lane21_strm1_cntl          ( std__pe19__lane21_strm1_cntl       ),      
               .std__pe19__lane21_strm1_data          ( std__pe19__lane21_strm1_data       ),      
               .std__pe19__lane21_strm1_data_valid    ( std__pe19__lane21_strm1_data_valid ),      
               .std__pe19__lane21_strm1_data_mask     ( std__pe19__lane21_strm1_data_mask  ),      

               // PE 19, Lane 22                 
               .pe19__std__lane22_strm0_ready         ( pe19__std__lane22_strm0_ready      ),      
               .std__pe19__lane22_strm0_cntl          ( std__pe19__lane22_strm0_cntl       ),      
               .std__pe19__lane22_strm0_data          ( std__pe19__lane22_strm0_data       ),      
               .std__pe19__lane22_strm0_data_valid    ( std__pe19__lane22_strm0_data_valid ),      
               .std__pe19__lane22_strm0_data_mask     ( std__pe19__lane22_strm0_data_mask  ),      

               .pe19__std__lane22_strm1_ready         ( pe19__std__lane22_strm1_ready      ),      
               .std__pe19__lane22_strm1_cntl          ( std__pe19__lane22_strm1_cntl       ),      
               .std__pe19__lane22_strm1_data          ( std__pe19__lane22_strm1_data       ),      
               .std__pe19__lane22_strm1_data_valid    ( std__pe19__lane22_strm1_data_valid ),      
               .std__pe19__lane22_strm1_data_mask     ( std__pe19__lane22_strm1_data_mask  ),      

               // PE 19, Lane 23                 
               .pe19__std__lane23_strm0_ready         ( pe19__std__lane23_strm0_ready      ),      
               .std__pe19__lane23_strm0_cntl          ( std__pe19__lane23_strm0_cntl       ),      
               .std__pe19__lane23_strm0_data          ( std__pe19__lane23_strm0_data       ),      
               .std__pe19__lane23_strm0_data_valid    ( std__pe19__lane23_strm0_data_valid ),      
               .std__pe19__lane23_strm0_data_mask     ( std__pe19__lane23_strm0_data_mask  ),      

               .pe19__std__lane23_strm1_ready         ( pe19__std__lane23_strm1_ready      ),      
               .std__pe19__lane23_strm1_cntl          ( std__pe19__lane23_strm1_cntl       ),      
               .std__pe19__lane23_strm1_data          ( std__pe19__lane23_strm1_data       ),      
               .std__pe19__lane23_strm1_data_valid    ( std__pe19__lane23_strm1_data_valid ),      
               .std__pe19__lane23_strm1_data_mask     ( std__pe19__lane23_strm1_data_mask  ),      

               // PE 19, Lane 24                 
               .pe19__std__lane24_strm0_ready         ( pe19__std__lane24_strm0_ready      ),      
               .std__pe19__lane24_strm0_cntl          ( std__pe19__lane24_strm0_cntl       ),      
               .std__pe19__lane24_strm0_data          ( std__pe19__lane24_strm0_data       ),      
               .std__pe19__lane24_strm0_data_valid    ( std__pe19__lane24_strm0_data_valid ),      
               .std__pe19__lane24_strm0_data_mask     ( std__pe19__lane24_strm0_data_mask  ),      

               .pe19__std__lane24_strm1_ready         ( pe19__std__lane24_strm1_ready      ),      
               .std__pe19__lane24_strm1_cntl          ( std__pe19__lane24_strm1_cntl       ),      
               .std__pe19__lane24_strm1_data          ( std__pe19__lane24_strm1_data       ),      
               .std__pe19__lane24_strm1_data_valid    ( std__pe19__lane24_strm1_data_valid ),      
               .std__pe19__lane24_strm1_data_mask     ( std__pe19__lane24_strm1_data_mask  ),      

               // PE 19, Lane 25                 
               .pe19__std__lane25_strm0_ready         ( pe19__std__lane25_strm0_ready      ),      
               .std__pe19__lane25_strm0_cntl          ( std__pe19__lane25_strm0_cntl       ),      
               .std__pe19__lane25_strm0_data          ( std__pe19__lane25_strm0_data       ),      
               .std__pe19__lane25_strm0_data_valid    ( std__pe19__lane25_strm0_data_valid ),      
               .std__pe19__lane25_strm0_data_mask     ( std__pe19__lane25_strm0_data_mask  ),      

               .pe19__std__lane25_strm1_ready         ( pe19__std__lane25_strm1_ready      ),      
               .std__pe19__lane25_strm1_cntl          ( std__pe19__lane25_strm1_cntl       ),      
               .std__pe19__lane25_strm1_data          ( std__pe19__lane25_strm1_data       ),      
               .std__pe19__lane25_strm1_data_valid    ( std__pe19__lane25_strm1_data_valid ),      
               .std__pe19__lane25_strm1_data_mask     ( std__pe19__lane25_strm1_data_mask  ),      

               // PE 19, Lane 26                 
               .pe19__std__lane26_strm0_ready         ( pe19__std__lane26_strm0_ready      ),      
               .std__pe19__lane26_strm0_cntl          ( std__pe19__lane26_strm0_cntl       ),      
               .std__pe19__lane26_strm0_data          ( std__pe19__lane26_strm0_data       ),      
               .std__pe19__lane26_strm0_data_valid    ( std__pe19__lane26_strm0_data_valid ),      
               .std__pe19__lane26_strm0_data_mask     ( std__pe19__lane26_strm0_data_mask  ),      

               .pe19__std__lane26_strm1_ready         ( pe19__std__lane26_strm1_ready      ),      
               .std__pe19__lane26_strm1_cntl          ( std__pe19__lane26_strm1_cntl       ),      
               .std__pe19__lane26_strm1_data          ( std__pe19__lane26_strm1_data       ),      
               .std__pe19__lane26_strm1_data_valid    ( std__pe19__lane26_strm1_data_valid ),      
               .std__pe19__lane26_strm1_data_mask     ( std__pe19__lane26_strm1_data_mask  ),      

               // PE 19, Lane 27                 
               .pe19__std__lane27_strm0_ready         ( pe19__std__lane27_strm0_ready      ),      
               .std__pe19__lane27_strm0_cntl          ( std__pe19__lane27_strm0_cntl       ),      
               .std__pe19__lane27_strm0_data          ( std__pe19__lane27_strm0_data       ),      
               .std__pe19__lane27_strm0_data_valid    ( std__pe19__lane27_strm0_data_valid ),      
               .std__pe19__lane27_strm0_data_mask     ( std__pe19__lane27_strm0_data_mask  ),      

               .pe19__std__lane27_strm1_ready         ( pe19__std__lane27_strm1_ready      ),      
               .std__pe19__lane27_strm1_cntl          ( std__pe19__lane27_strm1_cntl       ),      
               .std__pe19__lane27_strm1_data          ( std__pe19__lane27_strm1_data       ),      
               .std__pe19__lane27_strm1_data_valid    ( std__pe19__lane27_strm1_data_valid ),      
               .std__pe19__lane27_strm1_data_mask     ( std__pe19__lane27_strm1_data_mask  ),      

               // PE 19, Lane 28                 
               .pe19__std__lane28_strm0_ready         ( pe19__std__lane28_strm0_ready      ),      
               .std__pe19__lane28_strm0_cntl          ( std__pe19__lane28_strm0_cntl       ),      
               .std__pe19__lane28_strm0_data          ( std__pe19__lane28_strm0_data       ),      
               .std__pe19__lane28_strm0_data_valid    ( std__pe19__lane28_strm0_data_valid ),      
               .std__pe19__lane28_strm0_data_mask     ( std__pe19__lane28_strm0_data_mask  ),      

               .pe19__std__lane28_strm1_ready         ( pe19__std__lane28_strm1_ready      ),      
               .std__pe19__lane28_strm1_cntl          ( std__pe19__lane28_strm1_cntl       ),      
               .std__pe19__lane28_strm1_data          ( std__pe19__lane28_strm1_data       ),      
               .std__pe19__lane28_strm1_data_valid    ( std__pe19__lane28_strm1_data_valid ),      
               .std__pe19__lane28_strm1_data_mask     ( std__pe19__lane28_strm1_data_mask  ),      

               // PE 19, Lane 29                 
               .pe19__std__lane29_strm0_ready         ( pe19__std__lane29_strm0_ready      ),      
               .std__pe19__lane29_strm0_cntl          ( std__pe19__lane29_strm0_cntl       ),      
               .std__pe19__lane29_strm0_data          ( std__pe19__lane29_strm0_data       ),      
               .std__pe19__lane29_strm0_data_valid    ( std__pe19__lane29_strm0_data_valid ),      
               .std__pe19__lane29_strm0_data_mask     ( std__pe19__lane29_strm0_data_mask  ),      

               .pe19__std__lane29_strm1_ready         ( pe19__std__lane29_strm1_ready      ),      
               .std__pe19__lane29_strm1_cntl          ( std__pe19__lane29_strm1_cntl       ),      
               .std__pe19__lane29_strm1_data          ( std__pe19__lane29_strm1_data       ),      
               .std__pe19__lane29_strm1_data_valid    ( std__pe19__lane29_strm1_data_valid ),      
               .std__pe19__lane29_strm1_data_mask     ( std__pe19__lane29_strm1_data_mask  ),      

               // PE 19, Lane 30                 
               .pe19__std__lane30_strm0_ready         ( pe19__std__lane30_strm0_ready      ),      
               .std__pe19__lane30_strm0_cntl          ( std__pe19__lane30_strm0_cntl       ),      
               .std__pe19__lane30_strm0_data          ( std__pe19__lane30_strm0_data       ),      
               .std__pe19__lane30_strm0_data_valid    ( std__pe19__lane30_strm0_data_valid ),      
               .std__pe19__lane30_strm0_data_mask     ( std__pe19__lane30_strm0_data_mask  ),      

               .pe19__std__lane30_strm1_ready         ( pe19__std__lane30_strm1_ready      ),      
               .std__pe19__lane30_strm1_cntl          ( std__pe19__lane30_strm1_cntl       ),      
               .std__pe19__lane30_strm1_data          ( std__pe19__lane30_strm1_data       ),      
               .std__pe19__lane30_strm1_data_valid    ( std__pe19__lane30_strm1_data_valid ),      
               .std__pe19__lane30_strm1_data_mask     ( std__pe19__lane30_strm1_data_mask  ),      

               // PE 19, Lane 31                 
               .pe19__std__lane31_strm0_ready         ( pe19__std__lane31_strm0_ready      ),      
               .std__pe19__lane31_strm0_cntl          ( std__pe19__lane31_strm0_cntl       ),      
               .std__pe19__lane31_strm0_data          ( std__pe19__lane31_strm0_data       ),      
               .std__pe19__lane31_strm0_data_valid    ( std__pe19__lane31_strm0_data_valid ),      
               .std__pe19__lane31_strm0_data_mask     ( std__pe19__lane31_strm0_data_mask  ),      

               .pe19__std__lane31_strm1_ready         ( pe19__std__lane31_strm1_ready      ),      
               .std__pe19__lane31_strm1_cntl          ( std__pe19__lane31_strm1_cntl       ),      
               .std__pe19__lane31_strm1_data          ( std__pe19__lane31_strm1_data       ),      
               .std__pe19__lane31_strm1_data_valid    ( std__pe19__lane31_strm1_data_valid ),      
               .std__pe19__lane31_strm1_data_mask     ( std__pe19__lane31_strm1_data_mask  ),      

               // PE 20, Lane 0                 
               .pe20__std__lane0_strm0_ready         ( pe20__std__lane0_strm0_ready      ),      
               .std__pe20__lane0_strm0_cntl          ( std__pe20__lane0_strm0_cntl       ),      
               .std__pe20__lane0_strm0_data          ( std__pe20__lane0_strm0_data       ),      
               .std__pe20__lane0_strm0_data_valid    ( std__pe20__lane0_strm0_data_valid ),      
               .std__pe20__lane0_strm0_data_mask     ( std__pe20__lane0_strm0_data_mask  ),      

               .pe20__std__lane0_strm1_ready         ( pe20__std__lane0_strm1_ready      ),      
               .std__pe20__lane0_strm1_cntl          ( std__pe20__lane0_strm1_cntl       ),      
               .std__pe20__lane0_strm1_data          ( std__pe20__lane0_strm1_data       ),      
               .std__pe20__lane0_strm1_data_valid    ( std__pe20__lane0_strm1_data_valid ),      
               .std__pe20__lane0_strm1_data_mask     ( std__pe20__lane0_strm1_data_mask  ),      

               // PE 20, Lane 1                 
               .pe20__std__lane1_strm0_ready         ( pe20__std__lane1_strm0_ready      ),      
               .std__pe20__lane1_strm0_cntl          ( std__pe20__lane1_strm0_cntl       ),      
               .std__pe20__lane1_strm0_data          ( std__pe20__lane1_strm0_data       ),      
               .std__pe20__lane1_strm0_data_valid    ( std__pe20__lane1_strm0_data_valid ),      
               .std__pe20__lane1_strm0_data_mask     ( std__pe20__lane1_strm0_data_mask  ),      

               .pe20__std__lane1_strm1_ready         ( pe20__std__lane1_strm1_ready      ),      
               .std__pe20__lane1_strm1_cntl          ( std__pe20__lane1_strm1_cntl       ),      
               .std__pe20__lane1_strm1_data          ( std__pe20__lane1_strm1_data       ),      
               .std__pe20__lane1_strm1_data_valid    ( std__pe20__lane1_strm1_data_valid ),      
               .std__pe20__lane1_strm1_data_mask     ( std__pe20__lane1_strm1_data_mask  ),      

               // PE 20, Lane 2                 
               .pe20__std__lane2_strm0_ready         ( pe20__std__lane2_strm0_ready      ),      
               .std__pe20__lane2_strm0_cntl          ( std__pe20__lane2_strm0_cntl       ),      
               .std__pe20__lane2_strm0_data          ( std__pe20__lane2_strm0_data       ),      
               .std__pe20__lane2_strm0_data_valid    ( std__pe20__lane2_strm0_data_valid ),      
               .std__pe20__lane2_strm0_data_mask     ( std__pe20__lane2_strm0_data_mask  ),      

               .pe20__std__lane2_strm1_ready         ( pe20__std__lane2_strm1_ready      ),      
               .std__pe20__lane2_strm1_cntl          ( std__pe20__lane2_strm1_cntl       ),      
               .std__pe20__lane2_strm1_data          ( std__pe20__lane2_strm1_data       ),      
               .std__pe20__lane2_strm1_data_valid    ( std__pe20__lane2_strm1_data_valid ),      
               .std__pe20__lane2_strm1_data_mask     ( std__pe20__lane2_strm1_data_mask  ),      

               // PE 20, Lane 3                 
               .pe20__std__lane3_strm0_ready         ( pe20__std__lane3_strm0_ready      ),      
               .std__pe20__lane3_strm0_cntl          ( std__pe20__lane3_strm0_cntl       ),      
               .std__pe20__lane3_strm0_data          ( std__pe20__lane3_strm0_data       ),      
               .std__pe20__lane3_strm0_data_valid    ( std__pe20__lane3_strm0_data_valid ),      
               .std__pe20__lane3_strm0_data_mask     ( std__pe20__lane3_strm0_data_mask  ),      

               .pe20__std__lane3_strm1_ready         ( pe20__std__lane3_strm1_ready      ),      
               .std__pe20__lane3_strm1_cntl          ( std__pe20__lane3_strm1_cntl       ),      
               .std__pe20__lane3_strm1_data          ( std__pe20__lane3_strm1_data       ),      
               .std__pe20__lane3_strm1_data_valid    ( std__pe20__lane3_strm1_data_valid ),      
               .std__pe20__lane3_strm1_data_mask     ( std__pe20__lane3_strm1_data_mask  ),      

               // PE 20, Lane 4                 
               .pe20__std__lane4_strm0_ready         ( pe20__std__lane4_strm0_ready      ),      
               .std__pe20__lane4_strm0_cntl          ( std__pe20__lane4_strm0_cntl       ),      
               .std__pe20__lane4_strm0_data          ( std__pe20__lane4_strm0_data       ),      
               .std__pe20__lane4_strm0_data_valid    ( std__pe20__lane4_strm0_data_valid ),      
               .std__pe20__lane4_strm0_data_mask     ( std__pe20__lane4_strm0_data_mask  ),      

               .pe20__std__lane4_strm1_ready         ( pe20__std__lane4_strm1_ready      ),      
               .std__pe20__lane4_strm1_cntl          ( std__pe20__lane4_strm1_cntl       ),      
               .std__pe20__lane4_strm1_data          ( std__pe20__lane4_strm1_data       ),      
               .std__pe20__lane4_strm1_data_valid    ( std__pe20__lane4_strm1_data_valid ),      
               .std__pe20__lane4_strm1_data_mask     ( std__pe20__lane4_strm1_data_mask  ),      

               // PE 20, Lane 5                 
               .pe20__std__lane5_strm0_ready         ( pe20__std__lane5_strm0_ready      ),      
               .std__pe20__lane5_strm0_cntl          ( std__pe20__lane5_strm0_cntl       ),      
               .std__pe20__lane5_strm0_data          ( std__pe20__lane5_strm0_data       ),      
               .std__pe20__lane5_strm0_data_valid    ( std__pe20__lane5_strm0_data_valid ),      
               .std__pe20__lane5_strm0_data_mask     ( std__pe20__lane5_strm0_data_mask  ),      

               .pe20__std__lane5_strm1_ready         ( pe20__std__lane5_strm1_ready      ),      
               .std__pe20__lane5_strm1_cntl          ( std__pe20__lane5_strm1_cntl       ),      
               .std__pe20__lane5_strm1_data          ( std__pe20__lane5_strm1_data       ),      
               .std__pe20__lane5_strm1_data_valid    ( std__pe20__lane5_strm1_data_valid ),      
               .std__pe20__lane5_strm1_data_mask     ( std__pe20__lane5_strm1_data_mask  ),      

               // PE 20, Lane 6                 
               .pe20__std__lane6_strm0_ready         ( pe20__std__lane6_strm0_ready      ),      
               .std__pe20__lane6_strm0_cntl          ( std__pe20__lane6_strm0_cntl       ),      
               .std__pe20__lane6_strm0_data          ( std__pe20__lane6_strm0_data       ),      
               .std__pe20__lane6_strm0_data_valid    ( std__pe20__lane6_strm0_data_valid ),      
               .std__pe20__lane6_strm0_data_mask     ( std__pe20__lane6_strm0_data_mask  ),      

               .pe20__std__lane6_strm1_ready         ( pe20__std__lane6_strm1_ready      ),      
               .std__pe20__lane6_strm1_cntl          ( std__pe20__lane6_strm1_cntl       ),      
               .std__pe20__lane6_strm1_data          ( std__pe20__lane6_strm1_data       ),      
               .std__pe20__lane6_strm1_data_valid    ( std__pe20__lane6_strm1_data_valid ),      
               .std__pe20__lane6_strm1_data_mask     ( std__pe20__lane6_strm1_data_mask  ),      

               // PE 20, Lane 7                 
               .pe20__std__lane7_strm0_ready         ( pe20__std__lane7_strm0_ready      ),      
               .std__pe20__lane7_strm0_cntl          ( std__pe20__lane7_strm0_cntl       ),      
               .std__pe20__lane7_strm0_data          ( std__pe20__lane7_strm0_data       ),      
               .std__pe20__lane7_strm0_data_valid    ( std__pe20__lane7_strm0_data_valid ),      
               .std__pe20__lane7_strm0_data_mask     ( std__pe20__lane7_strm0_data_mask  ),      

               .pe20__std__lane7_strm1_ready         ( pe20__std__lane7_strm1_ready      ),      
               .std__pe20__lane7_strm1_cntl          ( std__pe20__lane7_strm1_cntl       ),      
               .std__pe20__lane7_strm1_data          ( std__pe20__lane7_strm1_data       ),      
               .std__pe20__lane7_strm1_data_valid    ( std__pe20__lane7_strm1_data_valid ),      
               .std__pe20__lane7_strm1_data_mask     ( std__pe20__lane7_strm1_data_mask  ),      

               // PE 20, Lane 8                 
               .pe20__std__lane8_strm0_ready         ( pe20__std__lane8_strm0_ready      ),      
               .std__pe20__lane8_strm0_cntl          ( std__pe20__lane8_strm0_cntl       ),      
               .std__pe20__lane8_strm0_data          ( std__pe20__lane8_strm0_data       ),      
               .std__pe20__lane8_strm0_data_valid    ( std__pe20__lane8_strm0_data_valid ),      
               .std__pe20__lane8_strm0_data_mask     ( std__pe20__lane8_strm0_data_mask  ),      

               .pe20__std__lane8_strm1_ready         ( pe20__std__lane8_strm1_ready      ),      
               .std__pe20__lane8_strm1_cntl          ( std__pe20__lane8_strm1_cntl       ),      
               .std__pe20__lane8_strm1_data          ( std__pe20__lane8_strm1_data       ),      
               .std__pe20__lane8_strm1_data_valid    ( std__pe20__lane8_strm1_data_valid ),      
               .std__pe20__lane8_strm1_data_mask     ( std__pe20__lane8_strm1_data_mask  ),      

               // PE 20, Lane 9                 
               .pe20__std__lane9_strm0_ready         ( pe20__std__lane9_strm0_ready      ),      
               .std__pe20__lane9_strm0_cntl          ( std__pe20__lane9_strm0_cntl       ),      
               .std__pe20__lane9_strm0_data          ( std__pe20__lane9_strm0_data       ),      
               .std__pe20__lane9_strm0_data_valid    ( std__pe20__lane9_strm0_data_valid ),      
               .std__pe20__lane9_strm0_data_mask     ( std__pe20__lane9_strm0_data_mask  ),      

               .pe20__std__lane9_strm1_ready         ( pe20__std__lane9_strm1_ready      ),      
               .std__pe20__lane9_strm1_cntl          ( std__pe20__lane9_strm1_cntl       ),      
               .std__pe20__lane9_strm1_data          ( std__pe20__lane9_strm1_data       ),      
               .std__pe20__lane9_strm1_data_valid    ( std__pe20__lane9_strm1_data_valid ),      
               .std__pe20__lane9_strm1_data_mask     ( std__pe20__lane9_strm1_data_mask  ),      

               // PE 20, Lane 10                 
               .pe20__std__lane10_strm0_ready         ( pe20__std__lane10_strm0_ready      ),      
               .std__pe20__lane10_strm0_cntl          ( std__pe20__lane10_strm0_cntl       ),      
               .std__pe20__lane10_strm0_data          ( std__pe20__lane10_strm0_data       ),      
               .std__pe20__lane10_strm0_data_valid    ( std__pe20__lane10_strm0_data_valid ),      
               .std__pe20__lane10_strm0_data_mask     ( std__pe20__lane10_strm0_data_mask  ),      

               .pe20__std__lane10_strm1_ready         ( pe20__std__lane10_strm1_ready      ),      
               .std__pe20__lane10_strm1_cntl          ( std__pe20__lane10_strm1_cntl       ),      
               .std__pe20__lane10_strm1_data          ( std__pe20__lane10_strm1_data       ),      
               .std__pe20__lane10_strm1_data_valid    ( std__pe20__lane10_strm1_data_valid ),      
               .std__pe20__lane10_strm1_data_mask     ( std__pe20__lane10_strm1_data_mask  ),      

               // PE 20, Lane 11                 
               .pe20__std__lane11_strm0_ready         ( pe20__std__lane11_strm0_ready      ),      
               .std__pe20__lane11_strm0_cntl          ( std__pe20__lane11_strm0_cntl       ),      
               .std__pe20__lane11_strm0_data          ( std__pe20__lane11_strm0_data       ),      
               .std__pe20__lane11_strm0_data_valid    ( std__pe20__lane11_strm0_data_valid ),      
               .std__pe20__lane11_strm0_data_mask     ( std__pe20__lane11_strm0_data_mask  ),      

               .pe20__std__lane11_strm1_ready         ( pe20__std__lane11_strm1_ready      ),      
               .std__pe20__lane11_strm1_cntl          ( std__pe20__lane11_strm1_cntl       ),      
               .std__pe20__lane11_strm1_data          ( std__pe20__lane11_strm1_data       ),      
               .std__pe20__lane11_strm1_data_valid    ( std__pe20__lane11_strm1_data_valid ),      
               .std__pe20__lane11_strm1_data_mask     ( std__pe20__lane11_strm1_data_mask  ),      

               // PE 20, Lane 12                 
               .pe20__std__lane12_strm0_ready         ( pe20__std__lane12_strm0_ready      ),      
               .std__pe20__lane12_strm0_cntl          ( std__pe20__lane12_strm0_cntl       ),      
               .std__pe20__lane12_strm0_data          ( std__pe20__lane12_strm0_data       ),      
               .std__pe20__lane12_strm0_data_valid    ( std__pe20__lane12_strm0_data_valid ),      
               .std__pe20__lane12_strm0_data_mask     ( std__pe20__lane12_strm0_data_mask  ),      

               .pe20__std__lane12_strm1_ready         ( pe20__std__lane12_strm1_ready      ),      
               .std__pe20__lane12_strm1_cntl          ( std__pe20__lane12_strm1_cntl       ),      
               .std__pe20__lane12_strm1_data          ( std__pe20__lane12_strm1_data       ),      
               .std__pe20__lane12_strm1_data_valid    ( std__pe20__lane12_strm1_data_valid ),      
               .std__pe20__lane12_strm1_data_mask     ( std__pe20__lane12_strm1_data_mask  ),      

               // PE 20, Lane 13                 
               .pe20__std__lane13_strm0_ready         ( pe20__std__lane13_strm0_ready      ),      
               .std__pe20__lane13_strm0_cntl          ( std__pe20__lane13_strm0_cntl       ),      
               .std__pe20__lane13_strm0_data          ( std__pe20__lane13_strm0_data       ),      
               .std__pe20__lane13_strm0_data_valid    ( std__pe20__lane13_strm0_data_valid ),      
               .std__pe20__lane13_strm0_data_mask     ( std__pe20__lane13_strm0_data_mask  ),      

               .pe20__std__lane13_strm1_ready         ( pe20__std__lane13_strm1_ready      ),      
               .std__pe20__lane13_strm1_cntl          ( std__pe20__lane13_strm1_cntl       ),      
               .std__pe20__lane13_strm1_data          ( std__pe20__lane13_strm1_data       ),      
               .std__pe20__lane13_strm1_data_valid    ( std__pe20__lane13_strm1_data_valid ),      
               .std__pe20__lane13_strm1_data_mask     ( std__pe20__lane13_strm1_data_mask  ),      

               // PE 20, Lane 14                 
               .pe20__std__lane14_strm0_ready         ( pe20__std__lane14_strm0_ready      ),      
               .std__pe20__lane14_strm0_cntl          ( std__pe20__lane14_strm0_cntl       ),      
               .std__pe20__lane14_strm0_data          ( std__pe20__lane14_strm0_data       ),      
               .std__pe20__lane14_strm0_data_valid    ( std__pe20__lane14_strm0_data_valid ),      
               .std__pe20__lane14_strm0_data_mask     ( std__pe20__lane14_strm0_data_mask  ),      

               .pe20__std__lane14_strm1_ready         ( pe20__std__lane14_strm1_ready      ),      
               .std__pe20__lane14_strm1_cntl          ( std__pe20__lane14_strm1_cntl       ),      
               .std__pe20__lane14_strm1_data          ( std__pe20__lane14_strm1_data       ),      
               .std__pe20__lane14_strm1_data_valid    ( std__pe20__lane14_strm1_data_valid ),      
               .std__pe20__lane14_strm1_data_mask     ( std__pe20__lane14_strm1_data_mask  ),      

               // PE 20, Lane 15                 
               .pe20__std__lane15_strm0_ready         ( pe20__std__lane15_strm0_ready      ),      
               .std__pe20__lane15_strm0_cntl          ( std__pe20__lane15_strm0_cntl       ),      
               .std__pe20__lane15_strm0_data          ( std__pe20__lane15_strm0_data       ),      
               .std__pe20__lane15_strm0_data_valid    ( std__pe20__lane15_strm0_data_valid ),      
               .std__pe20__lane15_strm0_data_mask     ( std__pe20__lane15_strm0_data_mask  ),      

               .pe20__std__lane15_strm1_ready         ( pe20__std__lane15_strm1_ready      ),      
               .std__pe20__lane15_strm1_cntl          ( std__pe20__lane15_strm1_cntl       ),      
               .std__pe20__lane15_strm1_data          ( std__pe20__lane15_strm1_data       ),      
               .std__pe20__lane15_strm1_data_valid    ( std__pe20__lane15_strm1_data_valid ),      
               .std__pe20__lane15_strm1_data_mask     ( std__pe20__lane15_strm1_data_mask  ),      

               // PE 20, Lane 16                 
               .pe20__std__lane16_strm0_ready         ( pe20__std__lane16_strm0_ready      ),      
               .std__pe20__lane16_strm0_cntl          ( std__pe20__lane16_strm0_cntl       ),      
               .std__pe20__lane16_strm0_data          ( std__pe20__lane16_strm0_data       ),      
               .std__pe20__lane16_strm0_data_valid    ( std__pe20__lane16_strm0_data_valid ),      
               .std__pe20__lane16_strm0_data_mask     ( std__pe20__lane16_strm0_data_mask  ),      

               .pe20__std__lane16_strm1_ready         ( pe20__std__lane16_strm1_ready      ),      
               .std__pe20__lane16_strm1_cntl          ( std__pe20__lane16_strm1_cntl       ),      
               .std__pe20__lane16_strm1_data          ( std__pe20__lane16_strm1_data       ),      
               .std__pe20__lane16_strm1_data_valid    ( std__pe20__lane16_strm1_data_valid ),      
               .std__pe20__lane16_strm1_data_mask     ( std__pe20__lane16_strm1_data_mask  ),      

               // PE 20, Lane 17                 
               .pe20__std__lane17_strm0_ready         ( pe20__std__lane17_strm0_ready      ),      
               .std__pe20__lane17_strm0_cntl          ( std__pe20__lane17_strm0_cntl       ),      
               .std__pe20__lane17_strm0_data          ( std__pe20__lane17_strm0_data       ),      
               .std__pe20__lane17_strm0_data_valid    ( std__pe20__lane17_strm0_data_valid ),      
               .std__pe20__lane17_strm0_data_mask     ( std__pe20__lane17_strm0_data_mask  ),      

               .pe20__std__lane17_strm1_ready         ( pe20__std__lane17_strm1_ready      ),      
               .std__pe20__lane17_strm1_cntl          ( std__pe20__lane17_strm1_cntl       ),      
               .std__pe20__lane17_strm1_data          ( std__pe20__lane17_strm1_data       ),      
               .std__pe20__lane17_strm1_data_valid    ( std__pe20__lane17_strm1_data_valid ),      
               .std__pe20__lane17_strm1_data_mask     ( std__pe20__lane17_strm1_data_mask  ),      

               // PE 20, Lane 18                 
               .pe20__std__lane18_strm0_ready         ( pe20__std__lane18_strm0_ready      ),      
               .std__pe20__lane18_strm0_cntl          ( std__pe20__lane18_strm0_cntl       ),      
               .std__pe20__lane18_strm0_data          ( std__pe20__lane18_strm0_data       ),      
               .std__pe20__lane18_strm0_data_valid    ( std__pe20__lane18_strm0_data_valid ),      
               .std__pe20__lane18_strm0_data_mask     ( std__pe20__lane18_strm0_data_mask  ),      

               .pe20__std__lane18_strm1_ready         ( pe20__std__lane18_strm1_ready      ),      
               .std__pe20__lane18_strm1_cntl          ( std__pe20__lane18_strm1_cntl       ),      
               .std__pe20__lane18_strm1_data          ( std__pe20__lane18_strm1_data       ),      
               .std__pe20__lane18_strm1_data_valid    ( std__pe20__lane18_strm1_data_valid ),      
               .std__pe20__lane18_strm1_data_mask     ( std__pe20__lane18_strm1_data_mask  ),      

               // PE 20, Lane 19                 
               .pe20__std__lane19_strm0_ready         ( pe20__std__lane19_strm0_ready      ),      
               .std__pe20__lane19_strm0_cntl          ( std__pe20__lane19_strm0_cntl       ),      
               .std__pe20__lane19_strm0_data          ( std__pe20__lane19_strm0_data       ),      
               .std__pe20__lane19_strm0_data_valid    ( std__pe20__lane19_strm0_data_valid ),      
               .std__pe20__lane19_strm0_data_mask     ( std__pe20__lane19_strm0_data_mask  ),      

               .pe20__std__lane19_strm1_ready         ( pe20__std__lane19_strm1_ready      ),      
               .std__pe20__lane19_strm1_cntl          ( std__pe20__lane19_strm1_cntl       ),      
               .std__pe20__lane19_strm1_data          ( std__pe20__lane19_strm1_data       ),      
               .std__pe20__lane19_strm1_data_valid    ( std__pe20__lane19_strm1_data_valid ),      
               .std__pe20__lane19_strm1_data_mask     ( std__pe20__lane19_strm1_data_mask  ),      

               // PE 20, Lane 20                 
               .pe20__std__lane20_strm0_ready         ( pe20__std__lane20_strm0_ready      ),      
               .std__pe20__lane20_strm0_cntl          ( std__pe20__lane20_strm0_cntl       ),      
               .std__pe20__lane20_strm0_data          ( std__pe20__lane20_strm0_data       ),      
               .std__pe20__lane20_strm0_data_valid    ( std__pe20__lane20_strm0_data_valid ),      
               .std__pe20__lane20_strm0_data_mask     ( std__pe20__lane20_strm0_data_mask  ),      

               .pe20__std__lane20_strm1_ready         ( pe20__std__lane20_strm1_ready      ),      
               .std__pe20__lane20_strm1_cntl          ( std__pe20__lane20_strm1_cntl       ),      
               .std__pe20__lane20_strm1_data          ( std__pe20__lane20_strm1_data       ),      
               .std__pe20__lane20_strm1_data_valid    ( std__pe20__lane20_strm1_data_valid ),      
               .std__pe20__lane20_strm1_data_mask     ( std__pe20__lane20_strm1_data_mask  ),      

               // PE 20, Lane 21                 
               .pe20__std__lane21_strm0_ready         ( pe20__std__lane21_strm0_ready      ),      
               .std__pe20__lane21_strm0_cntl          ( std__pe20__lane21_strm0_cntl       ),      
               .std__pe20__lane21_strm0_data          ( std__pe20__lane21_strm0_data       ),      
               .std__pe20__lane21_strm0_data_valid    ( std__pe20__lane21_strm0_data_valid ),      
               .std__pe20__lane21_strm0_data_mask     ( std__pe20__lane21_strm0_data_mask  ),      

               .pe20__std__lane21_strm1_ready         ( pe20__std__lane21_strm1_ready      ),      
               .std__pe20__lane21_strm1_cntl          ( std__pe20__lane21_strm1_cntl       ),      
               .std__pe20__lane21_strm1_data          ( std__pe20__lane21_strm1_data       ),      
               .std__pe20__lane21_strm1_data_valid    ( std__pe20__lane21_strm1_data_valid ),      
               .std__pe20__lane21_strm1_data_mask     ( std__pe20__lane21_strm1_data_mask  ),      

               // PE 20, Lane 22                 
               .pe20__std__lane22_strm0_ready         ( pe20__std__lane22_strm0_ready      ),      
               .std__pe20__lane22_strm0_cntl          ( std__pe20__lane22_strm0_cntl       ),      
               .std__pe20__lane22_strm0_data          ( std__pe20__lane22_strm0_data       ),      
               .std__pe20__lane22_strm0_data_valid    ( std__pe20__lane22_strm0_data_valid ),      
               .std__pe20__lane22_strm0_data_mask     ( std__pe20__lane22_strm0_data_mask  ),      

               .pe20__std__lane22_strm1_ready         ( pe20__std__lane22_strm1_ready      ),      
               .std__pe20__lane22_strm1_cntl          ( std__pe20__lane22_strm1_cntl       ),      
               .std__pe20__lane22_strm1_data          ( std__pe20__lane22_strm1_data       ),      
               .std__pe20__lane22_strm1_data_valid    ( std__pe20__lane22_strm1_data_valid ),      
               .std__pe20__lane22_strm1_data_mask     ( std__pe20__lane22_strm1_data_mask  ),      

               // PE 20, Lane 23                 
               .pe20__std__lane23_strm0_ready         ( pe20__std__lane23_strm0_ready      ),      
               .std__pe20__lane23_strm0_cntl          ( std__pe20__lane23_strm0_cntl       ),      
               .std__pe20__lane23_strm0_data          ( std__pe20__lane23_strm0_data       ),      
               .std__pe20__lane23_strm0_data_valid    ( std__pe20__lane23_strm0_data_valid ),      
               .std__pe20__lane23_strm0_data_mask     ( std__pe20__lane23_strm0_data_mask  ),      

               .pe20__std__lane23_strm1_ready         ( pe20__std__lane23_strm1_ready      ),      
               .std__pe20__lane23_strm1_cntl          ( std__pe20__lane23_strm1_cntl       ),      
               .std__pe20__lane23_strm1_data          ( std__pe20__lane23_strm1_data       ),      
               .std__pe20__lane23_strm1_data_valid    ( std__pe20__lane23_strm1_data_valid ),      
               .std__pe20__lane23_strm1_data_mask     ( std__pe20__lane23_strm1_data_mask  ),      

               // PE 20, Lane 24                 
               .pe20__std__lane24_strm0_ready         ( pe20__std__lane24_strm0_ready      ),      
               .std__pe20__lane24_strm0_cntl          ( std__pe20__lane24_strm0_cntl       ),      
               .std__pe20__lane24_strm0_data          ( std__pe20__lane24_strm0_data       ),      
               .std__pe20__lane24_strm0_data_valid    ( std__pe20__lane24_strm0_data_valid ),      
               .std__pe20__lane24_strm0_data_mask     ( std__pe20__lane24_strm0_data_mask  ),      

               .pe20__std__lane24_strm1_ready         ( pe20__std__lane24_strm1_ready      ),      
               .std__pe20__lane24_strm1_cntl          ( std__pe20__lane24_strm1_cntl       ),      
               .std__pe20__lane24_strm1_data          ( std__pe20__lane24_strm1_data       ),      
               .std__pe20__lane24_strm1_data_valid    ( std__pe20__lane24_strm1_data_valid ),      
               .std__pe20__lane24_strm1_data_mask     ( std__pe20__lane24_strm1_data_mask  ),      

               // PE 20, Lane 25                 
               .pe20__std__lane25_strm0_ready         ( pe20__std__lane25_strm0_ready      ),      
               .std__pe20__lane25_strm0_cntl          ( std__pe20__lane25_strm0_cntl       ),      
               .std__pe20__lane25_strm0_data          ( std__pe20__lane25_strm0_data       ),      
               .std__pe20__lane25_strm0_data_valid    ( std__pe20__lane25_strm0_data_valid ),      
               .std__pe20__lane25_strm0_data_mask     ( std__pe20__lane25_strm0_data_mask  ),      

               .pe20__std__lane25_strm1_ready         ( pe20__std__lane25_strm1_ready      ),      
               .std__pe20__lane25_strm1_cntl          ( std__pe20__lane25_strm1_cntl       ),      
               .std__pe20__lane25_strm1_data          ( std__pe20__lane25_strm1_data       ),      
               .std__pe20__lane25_strm1_data_valid    ( std__pe20__lane25_strm1_data_valid ),      
               .std__pe20__lane25_strm1_data_mask     ( std__pe20__lane25_strm1_data_mask  ),      

               // PE 20, Lane 26                 
               .pe20__std__lane26_strm0_ready         ( pe20__std__lane26_strm0_ready      ),      
               .std__pe20__lane26_strm0_cntl          ( std__pe20__lane26_strm0_cntl       ),      
               .std__pe20__lane26_strm0_data          ( std__pe20__lane26_strm0_data       ),      
               .std__pe20__lane26_strm0_data_valid    ( std__pe20__lane26_strm0_data_valid ),      
               .std__pe20__lane26_strm0_data_mask     ( std__pe20__lane26_strm0_data_mask  ),      

               .pe20__std__lane26_strm1_ready         ( pe20__std__lane26_strm1_ready      ),      
               .std__pe20__lane26_strm1_cntl          ( std__pe20__lane26_strm1_cntl       ),      
               .std__pe20__lane26_strm1_data          ( std__pe20__lane26_strm1_data       ),      
               .std__pe20__lane26_strm1_data_valid    ( std__pe20__lane26_strm1_data_valid ),      
               .std__pe20__lane26_strm1_data_mask     ( std__pe20__lane26_strm1_data_mask  ),      

               // PE 20, Lane 27                 
               .pe20__std__lane27_strm0_ready         ( pe20__std__lane27_strm0_ready      ),      
               .std__pe20__lane27_strm0_cntl          ( std__pe20__lane27_strm0_cntl       ),      
               .std__pe20__lane27_strm0_data          ( std__pe20__lane27_strm0_data       ),      
               .std__pe20__lane27_strm0_data_valid    ( std__pe20__lane27_strm0_data_valid ),      
               .std__pe20__lane27_strm0_data_mask     ( std__pe20__lane27_strm0_data_mask  ),      

               .pe20__std__lane27_strm1_ready         ( pe20__std__lane27_strm1_ready      ),      
               .std__pe20__lane27_strm1_cntl          ( std__pe20__lane27_strm1_cntl       ),      
               .std__pe20__lane27_strm1_data          ( std__pe20__lane27_strm1_data       ),      
               .std__pe20__lane27_strm1_data_valid    ( std__pe20__lane27_strm1_data_valid ),      
               .std__pe20__lane27_strm1_data_mask     ( std__pe20__lane27_strm1_data_mask  ),      

               // PE 20, Lane 28                 
               .pe20__std__lane28_strm0_ready         ( pe20__std__lane28_strm0_ready      ),      
               .std__pe20__lane28_strm0_cntl          ( std__pe20__lane28_strm0_cntl       ),      
               .std__pe20__lane28_strm0_data          ( std__pe20__lane28_strm0_data       ),      
               .std__pe20__lane28_strm0_data_valid    ( std__pe20__lane28_strm0_data_valid ),      
               .std__pe20__lane28_strm0_data_mask     ( std__pe20__lane28_strm0_data_mask  ),      

               .pe20__std__lane28_strm1_ready         ( pe20__std__lane28_strm1_ready      ),      
               .std__pe20__lane28_strm1_cntl          ( std__pe20__lane28_strm1_cntl       ),      
               .std__pe20__lane28_strm1_data          ( std__pe20__lane28_strm1_data       ),      
               .std__pe20__lane28_strm1_data_valid    ( std__pe20__lane28_strm1_data_valid ),      
               .std__pe20__lane28_strm1_data_mask     ( std__pe20__lane28_strm1_data_mask  ),      

               // PE 20, Lane 29                 
               .pe20__std__lane29_strm0_ready         ( pe20__std__lane29_strm0_ready      ),      
               .std__pe20__lane29_strm0_cntl          ( std__pe20__lane29_strm0_cntl       ),      
               .std__pe20__lane29_strm0_data          ( std__pe20__lane29_strm0_data       ),      
               .std__pe20__lane29_strm0_data_valid    ( std__pe20__lane29_strm0_data_valid ),      
               .std__pe20__lane29_strm0_data_mask     ( std__pe20__lane29_strm0_data_mask  ),      

               .pe20__std__lane29_strm1_ready         ( pe20__std__lane29_strm1_ready      ),      
               .std__pe20__lane29_strm1_cntl          ( std__pe20__lane29_strm1_cntl       ),      
               .std__pe20__lane29_strm1_data          ( std__pe20__lane29_strm1_data       ),      
               .std__pe20__lane29_strm1_data_valid    ( std__pe20__lane29_strm1_data_valid ),      
               .std__pe20__lane29_strm1_data_mask     ( std__pe20__lane29_strm1_data_mask  ),      

               // PE 20, Lane 30                 
               .pe20__std__lane30_strm0_ready         ( pe20__std__lane30_strm0_ready      ),      
               .std__pe20__lane30_strm0_cntl          ( std__pe20__lane30_strm0_cntl       ),      
               .std__pe20__lane30_strm0_data          ( std__pe20__lane30_strm0_data       ),      
               .std__pe20__lane30_strm0_data_valid    ( std__pe20__lane30_strm0_data_valid ),      
               .std__pe20__lane30_strm0_data_mask     ( std__pe20__lane30_strm0_data_mask  ),      

               .pe20__std__lane30_strm1_ready         ( pe20__std__lane30_strm1_ready      ),      
               .std__pe20__lane30_strm1_cntl          ( std__pe20__lane30_strm1_cntl       ),      
               .std__pe20__lane30_strm1_data          ( std__pe20__lane30_strm1_data       ),      
               .std__pe20__lane30_strm1_data_valid    ( std__pe20__lane30_strm1_data_valid ),      
               .std__pe20__lane30_strm1_data_mask     ( std__pe20__lane30_strm1_data_mask  ),      

               // PE 20, Lane 31                 
               .pe20__std__lane31_strm0_ready         ( pe20__std__lane31_strm0_ready      ),      
               .std__pe20__lane31_strm0_cntl          ( std__pe20__lane31_strm0_cntl       ),      
               .std__pe20__lane31_strm0_data          ( std__pe20__lane31_strm0_data       ),      
               .std__pe20__lane31_strm0_data_valid    ( std__pe20__lane31_strm0_data_valid ),      
               .std__pe20__lane31_strm0_data_mask     ( std__pe20__lane31_strm0_data_mask  ),      

               .pe20__std__lane31_strm1_ready         ( pe20__std__lane31_strm1_ready      ),      
               .std__pe20__lane31_strm1_cntl          ( std__pe20__lane31_strm1_cntl       ),      
               .std__pe20__lane31_strm1_data          ( std__pe20__lane31_strm1_data       ),      
               .std__pe20__lane31_strm1_data_valid    ( std__pe20__lane31_strm1_data_valid ),      
               .std__pe20__lane31_strm1_data_mask     ( std__pe20__lane31_strm1_data_mask  ),      

               // PE 21, Lane 0                 
               .pe21__std__lane0_strm0_ready         ( pe21__std__lane0_strm0_ready      ),      
               .std__pe21__lane0_strm0_cntl          ( std__pe21__lane0_strm0_cntl       ),      
               .std__pe21__lane0_strm0_data          ( std__pe21__lane0_strm0_data       ),      
               .std__pe21__lane0_strm0_data_valid    ( std__pe21__lane0_strm0_data_valid ),      
               .std__pe21__lane0_strm0_data_mask     ( std__pe21__lane0_strm0_data_mask  ),      

               .pe21__std__lane0_strm1_ready         ( pe21__std__lane0_strm1_ready      ),      
               .std__pe21__lane0_strm1_cntl          ( std__pe21__lane0_strm1_cntl       ),      
               .std__pe21__lane0_strm1_data          ( std__pe21__lane0_strm1_data       ),      
               .std__pe21__lane0_strm1_data_valid    ( std__pe21__lane0_strm1_data_valid ),      
               .std__pe21__lane0_strm1_data_mask     ( std__pe21__lane0_strm1_data_mask  ),      

               // PE 21, Lane 1                 
               .pe21__std__lane1_strm0_ready         ( pe21__std__lane1_strm0_ready      ),      
               .std__pe21__lane1_strm0_cntl          ( std__pe21__lane1_strm0_cntl       ),      
               .std__pe21__lane1_strm0_data          ( std__pe21__lane1_strm0_data       ),      
               .std__pe21__lane1_strm0_data_valid    ( std__pe21__lane1_strm0_data_valid ),      
               .std__pe21__lane1_strm0_data_mask     ( std__pe21__lane1_strm0_data_mask  ),      

               .pe21__std__lane1_strm1_ready         ( pe21__std__lane1_strm1_ready      ),      
               .std__pe21__lane1_strm1_cntl          ( std__pe21__lane1_strm1_cntl       ),      
               .std__pe21__lane1_strm1_data          ( std__pe21__lane1_strm1_data       ),      
               .std__pe21__lane1_strm1_data_valid    ( std__pe21__lane1_strm1_data_valid ),      
               .std__pe21__lane1_strm1_data_mask     ( std__pe21__lane1_strm1_data_mask  ),      

               // PE 21, Lane 2                 
               .pe21__std__lane2_strm0_ready         ( pe21__std__lane2_strm0_ready      ),      
               .std__pe21__lane2_strm0_cntl          ( std__pe21__lane2_strm0_cntl       ),      
               .std__pe21__lane2_strm0_data          ( std__pe21__lane2_strm0_data       ),      
               .std__pe21__lane2_strm0_data_valid    ( std__pe21__lane2_strm0_data_valid ),      
               .std__pe21__lane2_strm0_data_mask     ( std__pe21__lane2_strm0_data_mask  ),      

               .pe21__std__lane2_strm1_ready         ( pe21__std__lane2_strm1_ready      ),      
               .std__pe21__lane2_strm1_cntl          ( std__pe21__lane2_strm1_cntl       ),      
               .std__pe21__lane2_strm1_data          ( std__pe21__lane2_strm1_data       ),      
               .std__pe21__lane2_strm1_data_valid    ( std__pe21__lane2_strm1_data_valid ),      
               .std__pe21__lane2_strm1_data_mask     ( std__pe21__lane2_strm1_data_mask  ),      

               // PE 21, Lane 3                 
               .pe21__std__lane3_strm0_ready         ( pe21__std__lane3_strm0_ready      ),      
               .std__pe21__lane3_strm0_cntl          ( std__pe21__lane3_strm0_cntl       ),      
               .std__pe21__lane3_strm0_data          ( std__pe21__lane3_strm0_data       ),      
               .std__pe21__lane3_strm0_data_valid    ( std__pe21__lane3_strm0_data_valid ),      
               .std__pe21__lane3_strm0_data_mask     ( std__pe21__lane3_strm0_data_mask  ),      

               .pe21__std__lane3_strm1_ready         ( pe21__std__lane3_strm1_ready      ),      
               .std__pe21__lane3_strm1_cntl          ( std__pe21__lane3_strm1_cntl       ),      
               .std__pe21__lane3_strm1_data          ( std__pe21__lane3_strm1_data       ),      
               .std__pe21__lane3_strm1_data_valid    ( std__pe21__lane3_strm1_data_valid ),      
               .std__pe21__lane3_strm1_data_mask     ( std__pe21__lane3_strm1_data_mask  ),      

               // PE 21, Lane 4                 
               .pe21__std__lane4_strm0_ready         ( pe21__std__lane4_strm0_ready      ),      
               .std__pe21__lane4_strm0_cntl          ( std__pe21__lane4_strm0_cntl       ),      
               .std__pe21__lane4_strm0_data          ( std__pe21__lane4_strm0_data       ),      
               .std__pe21__lane4_strm0_data_valid    ( std__pe21__lane4_strm0_data_valid ),      
               .std__pe21__lane4_strm0_data_mask     ( std__pe21__lane4_strm0_data_mask  ),      

               .pe21__std__lane4_strm1_ready         ( pe21__std__lane4_strm1_ready      ),      
               .std__pe21__lane4_strm1_cntl          ( std__pe21__lane4_strm1_cntl       ),      
               .std__pe21__lane4_strm1_data          ( std__pe21__lane4_strm1_data       ),      
               .std__pe21__lane4_strm1_data_valid    ( std__pe21__lane4_strm1_data_valid ),      
               .std__pe21__lane4_strm1_data_mask     ( std__pe21__lane4_strm1_data_mask  ),      

               // PE 21, Lane 5                 
               .pe21__std__lane5_strm0_ready         ( pe21__std__lane5_strm0_ready      ),      
               .std__pe21__lane5_strm0_cntl          ( std__pe21__lane5_strm0_cntl       ),      
               .std__pe21__lane5_strm0_data          ( std__pe21__lane5_strm0_data       ),      
               .std__pe21__lane5_strm0_data_valid    ( std__pe21__lane5_strm0_data_valid ),      
               .std__pe21__lane5_strm0_data_mask     ( std__pe21__lane5_strm0_data_mask  ),      

               .pe21__std__lane5_strm1_ready         ( pe21__std__lane5_strm1_ready      ),      
               .std__pe21__lane5_strm1_cntl          ( std__pe21__lane5_strm1_cntl       ),      
               .std__pe21__lane5_strm1_data          ( std__pe21__lane5_strm1_data       ),      
               .std__pe21__lane5_strm1_data_valid    ( std__pe21__lane5_strm1_data_valid ),      
               .std__pe21__lane5_strm1_data_mask     ( std__pe21__lane5_strm1_data_mask  ),      

               // PE 21, Lane 6                 
               .pe21__std__lane6_strm0_ready         ( pe21__std__lane6_strm0_ready      ),      
               .std__pe21__lane6_strm0_cntl          ( std__pe21__lane6_strm0_cntl       ),      
               .std__pe21__lane6_strm0_data          ( std__pe21__lane6_strm0_data       ),      
               .std__pe21__lane6_strm0_data_valid    ( std__pe21__lane6_strm0_data_valid ),      
               .std__pe21__lane6_strm0_data_mask     ( std__pe21__lane6_strm0_data_mask  ),      

               .pe21__std__lane6_strm1_ready         ( pe21__std__lane6_strm1_ready      ),      
               .std__pe21__lane6_strm1_cntl          ( std__pe21__lane6_strm1_cntl       ),      
               .std__pe21__lane6_strm1_data          ( std__pe21__lane6_strm1_data       ),      
               .std__pe21__lane6_strm1_data_valid    ( std__pe21__lane6_strm1_data_valid ),      
               .std__pe21__lane6_strm1_data_mask     ( std__pe21__lane6_strm1_data_mask  ),      

               // PE 21, Lane 7                 
               .pe21__std__lane7_strm0_ready         ( pe21__std__lane7_strm0_ready      ),      
               .std__pe21__lane7_strm0_cntl          ( std__pe21__lane7_strm0_cntl       ),      
               .std__pe21__lane7_strm0_data          ( std__pe21__lane7_strm0_data       ),      
               .std__pe21__lane7_strm0_data_valid    ( std__pe21__lane7_strm0_data_valid ),      
               .std__pe21__lane7_strm0_data_mask     ( std__pe21__lane7_strm0_data_mask  ),      

               .pe21__std__lane7_strm1_ready         ( pe21__std__lane7_strm1_ready      ),      
               .std__pe21__lane7_strm1_cntl          ( std__pe21__lane7_strm1_cntl       ),      
               .std__pe21__lane7_strm1_data          ( std__pe21__lane7_strm1_data       ),      
               .std__pe21__lane7_strm1_data_valid    ( std__pe21__lane7_strm1_data_valid ),      
               .std__pe21__lane7_strm1_data_mask     ( std__pe21__lane7_strm1_data_mask  ),      

               // PE 21, Lane 8                 
               .pe21__std__lane8_strm0_ready         ( pe21__std__lane8_strm0_ready      ),      
               .std__pe21__lane8_strm0_cntl          ( std__pe21__lane8_strm0_cntl       ),      
               .std__pe21__lane8_strm0_data          ( std__pe21__lane8_strm0_data       ),      
               .std__pe21__lane8_strm0_data_valid    ( std__pe21__lane8_strm0_data_valid ),      
               .std__pe21__lane8_strm0_data_mask     ( std__pe21__lane8_strm0_data_mask  ),      

               .pe21__std__lane8_strm1_ready         ( pe21__std__lane8_strm1_ready      ),      
               .std__pe21__lane8_strm1_cntl          ( std__pe21__lane8_strm1_cntl       ),      
               .std__pe21__lane8_strm1_data          ( std__pe21__lane8_strm1_data       ),      
               .std__pe21__lane8_strm1_data_valid    ( std__pe21__lane8_strm1_data_valid ),      
               .std__pe21__lane8_strm1_data_mask     ( std__pe21__lane8_strm1_data_mask  ),      

               // PE 21, Lane 9                 
               .pe21__std__lane9_strm0_ready         ( pe21__std__lane9_strm0_ready      ),      
               .std__pe21__lane9_strm0_cntl          ( std__pe21__lane9_strm0_cntl       ),      
               .std__pe21__lane9_strm0_data          ( std__pe21__lane9_strm0_data       ),      
               .std__pe21__lane9_strm0_data_valid    ( std__pe21__lane9_strm0_data_valid ),      
               .std__pe21__lane9_strm0_data_mask     ( std__pe21__lane9_strm0_data_mask  ),      

               .pe21__std__lane9_strm1_ready         ( pe21__std__lane9_strm1_ready      ),      
               .std__pe21__lane9_strm1_cntl          ( std__pe21__lane9_strm1_cntl       ),      
               .std__pe21__lane9_strm1_data          ( std__pe21__lane9_strm1_data       ),      
               .std__pe21__lane9_strm1_data_valid    ( std__pe21__lane9_strm1_data_valid ),      
               .std__pe21__lane9_strm1_data_mask     ( std__pe21__lane9_strm1_data_mask  ),      

               // PE 21, Lane 10                 
               .pe21__std__lane10_strm0_ready         ( pe21__std__lane10_strm0_ready      ),      
               .std__pe21__lane10_strm0_cntl          ( std__pe21__lane10_strm0_cntl       ),      
               .std__pe21__lane10_strm0_data          ( std__pe21__lane10_strm0_data       ),      
               .std__pe21__lane10_strm0_data_valid    ( std__pe21__lane10_strm0_data_valid ),      
               .std__pe21__lane10_strm0_data_mask     ( std__pe21__lane10_strm0_data_mask  ),      

               .pe21__std__lane10_strm1_ready         ( pe21__std__lane10_strm1_ready      ),      
               .std__pe21__lane10_strm1_cntl          ( std__pe21__lane10_strm1_cntl       ),      
               .std__pe21__lane10_strm1_data          ( std__pe21__lane10_strm1_data       ),      
               .std__pe21__lane10_strm1_data_valid    ( std__pe21__lane10_strm1_data_valid ),      
               .std__pe21__lane10_strm1_data_mask     ( std__pe21__lane10_strm1_data_mask  ),      

               // PE 21, Lane 11                 
               .pe21__std__lane11_strm0_ready         ( pe21__std__lane11_strm0_ready      ),      
               .std__pe21__lane11_strm0_cntl          ( std__pe21__lane11_strm0_cntl       ),      
               .std__pe21__lane11_strm0_data          ( std__pe21__lane11_strm0_data       ),      
               .std__pe21__lane11_strm0_data_valid    ( std__pe21__lane11_strm0_data_valid ),      
               .std__pe21__lane11_strm0_data_mask     ( std__pe21__lane11_strm0_data_mask  ),      

               .pe21__std__lane11_strm1_ready         ( pe21__std__lane11_strm1_ready      ),      
               .std__pe21__lane11_strm1_cntl          ( std__pe21__lane11_strm1_cntl       ),      
               .std__pe21__lane11_strm1_data          ( std__pe21__lane11_strm1_data       ),      
               .std__pe21__lane11_strm1_data_valid    ( std__pe21__lane11_strm1_data_valid ),      
               .std__pe21__lane11_strm1_data_mask     ( std__pe21__lane11_strm1_data_mask  ),      

               // PE 21, Lane 12                 
               .pe21__std__lane12_strm0_ready         ( pe21__std__lane12_strm0_ready      ),      
               .std__pe21__lane12_strm0_cntl          ( std__pe21__lane12_strm0_cntl       ),      
               .std__pe21__lane12_strm0_data          ( std__pe21__lane12_strm0_data       ),      
               .std__pe21__lane12_strm0_data_valid    ( std__pe21__lane12_strm0_data_valid ),      
               .std__pe21__lane12_strm0_data_mask     ( std__pe21__lane12_strm0_data_mask  ),      

               .pe21__std__lane12_strm1_ready         ( pe21__std__lane12_strm1_ready      ),      
               .std__pe21__lane12_strm1_cntl          ( std__pe21__lane12_strm1_cntl       ),      
               .std__pe21__lane12_strm1_data          ( std__pe21__lane12_strm1_data       ),      
               .std__pe21__lane12_strm1_data_valid    ( std__pe21__lane12_strm1_data_valid ),      
               .std__pe21__lane12_strm1_data_mask     ( std__pe21__lane12_strm1_data_mask  ),      

               // PE 21, Lane 13                 
               .pe21__std__lane13_strm0_ready         ( pe21__std__lane13_strm0_ready      ),      
               .std__pe21__lane13_strm0_cntl          ( std__pe21__lane13_strm0_cntl       ),      
               .std__pe21__lane13_strm0_data          ( std__pe21__lane13_strm0_data       ),      
               .std__pe21__lane13_strm0_data_valid    ( std__pe21__lane13_strm0_data_valid ),      
               .std__pe21__lane13_strm0_data_mask     ( std__pe21__lane13_strm0_data_mask  ),      

               .pe21__std__lane13_strm1_ready         ( pe21__std__lane13_strm1_ready      ),      
               .std__pe21__lane13_strm1_cntl          ( std__pe21__lane13_strm1_cntl       ),      
               .std__pe21__lane13_strm1_data          ( std__pe21__lane13_strm1_data       ),      
               .std__pe21__lane13_strm1_data_valid    ( std__pe21__lane13_strm1_data_valid ),      
               .std__pe21__lane13_strm1_data_mask     ( std__pe21__lane13_strm1_data_mask  ),      

               // PE 21, Lane 14                 
               .pe21__std__lane14_strm0_ready         ( pe21__std__lane14_strm0_ready      ),      
               .std__pe21__lane14_strm0_cntl          ( std__pe21__lane14_strm0_cntl       ),      
               .std__pe21__lane14_strm0_data          ( std__pe21__lane14_strm0_data       ),      
               .std__pe21__lane14_strm0_data_valid    ( std__pe21__lane14_strm0_data_valid ),      
               .std__pe21__lane14_strm0_data_mask     ( std__pe21__lane14_strm0_data_mask  ),      

               .pe21__std__lane14_strm1_ready         ( pe21__std__lane14_strm1_ready      ),      
               .std__pe21__lane14_strm1_cntl          ( std__pe21__lane14_strm1_cntl       ),      
               .std__pe21__lane14_strm1_data          ( std__pe21__lane14_strm1_data       ),      
               .std__pe21__lane14_strm1_data_valid    ( std__pe21__lane14_strm1_data_valid ),      
               .std__pe21__lane14_strm1_data_mask     ( std__pe21__lane14_strm1_data_mask  ),      

               // PE 21, Lane 15                 
               .pe21__std__lane15_strm0_ready         ( pe21__std__lane15_strm0_ready      ),      
               .std__pe21__lane15_strm0_cntl          ( std__pe21__lane15_strm0_cntl       ),      
               .std__pe21__lane15_strm0_data          ( std__pe21__lane15_strm0_data       ),      
               .std__pe21__lane15_strm0_data_valid    ( std__pe21__lane15_strm0_data_valid ),      
               .std__pe21__lane15_strm0_data_mask     ( std__pe21__lane15_strm0_data_mask  ),      

               .pe21__std__lane15_strm1_ready         ( pe21__std__lane15_strm1_ready      ),      
               .std__pe21__lane15_strm1_cntl          ( std__pe21__lane15_strm1_cntl       ),      
               .std__pe21__lane15_strm1_data          ( std__pe21__lane15_strm1_data       ),      
               .std__pe21__lane15_strm1_data_valid    ( std__pe21__lane15_strm1_data_valid ),      
               .std__pe21__lane15_strm1_data_mask     ( std__pe21__lane15_strm1_data_mask  ),      

               // PE 21, Lane 16                 
               .pe21__std__lane16_strm0_ready         ( pe21__std__lane16_strm0_ready      ),      
               .std__pe21__lane16_strm0_cntl          ( std__pe21__lane16_strm0_cntl       ),      
               .std__pe21__lane16_strm0_data          ( std__pe21__lane16_strm0_data       ),      
               .std__pe21__lane16_strm0_data_valid    ( std__pe21__lane16_strm0_data_valid ),      
               .std__pe21__lane16_strm0_data_mask     ( std__pe21__lane16_strm0_data_mask  ),      

               .pe21__std__lane16_strm1_ready         ( pe21__std__lane16_strm1_ready      ),      
               .std__pe21__lane16_strm1_cntl          ( std__pe21__lane16_strm1_cntl       ),      
               .std__pe21__lane16_strm1_data          ( std__pe21__lane16_strm1_data       ),      
               .std__pe21__lane16_strm1_data_valid    ( std__pe21__lane16_strm1_data_valid ),      
               .std__pe21__lane16_strm1_data_mask     ( std__pe21__lane16_strm1_data_mask  ),      

               // PE 21, Lane 17                 
               .pe21__std__lane17_strm0_ready         ( pe21__std__lane17_strm0_ready      ),      
               .std__pe21__lane17_strm0_cntl          ( std__pe21__lane17_strm0_cntl       ),      
               .std__pe21__lane17_strm0_data          ( std__pe21__lane17_strm0_data       ),      
               .std__pe21__lane17_strm0_data_valid    ( std__pe21__lane17_strm0_data_valid ),      
               .std__pe21__lane17_strm0_data_mask     ( std__pe21__lane17_strm0_data_mask  ),      

               .pe21__std__lane17_strm1_ready         ( pe21__std__lane17_strm1_ready      ),      
               .std__pe21__lane17_strm1_cntl          ( std__pe21__lane17_strm1_cntl       ),      
               .std__pe21__lane17_strm1_data          ( std__pe21__lane17_strm1_data       ),      
               .std__pe21__lane17_strm1_data_valid    ( std__pe21__lane17_strm1_data_valid ),      
               .std__pe21__lane17_strm1_data_mask     ( std__pe21__lane17_strm1_data_mask  ),      

               // PE 21, Lane 18                 
               .pe21__std__lane18_strm0_ready         ( pe21__std__lane18_strm0_ready      ),      
               .std__pe21__lane18_strm0_cntl          ( std__pe21__lane18_strm0_cntl       ),      
               .std__pe21__lane18_strm0_data          ( std__pe21__lane18_strm0_data       ),      
               .std__pe21__lane18_strm0_data_valid    ( std__pe21__lane18_strm0_data_valid ),      
               .std__pe21__lane18_strm0_data_mask     ( std__pe21__lane18_strm0_data_mask  ),      

               .pe21__std__lane18_strm1_ready         ( pe21__std__lane18_strm1_ready      ),      
               .std__pe21__lane18_strm1_cntl          ( std__pe21__lane18_strm1_cntl       ),      
               .std__pe21__lane18_strm1_data          ( std__pe21__lane18_strm1_data       ),      
               .std__pe21__lane18_strm1_data_valid    ( std__pe21__lane18_strm1_data_valid ),      
               .std__pe21__lane18_strm1_data_mask     ( std__pe21__lane18_strm1_data_mask  ),      

               // PE 21, Lane 19                 
               .pe21__std__lane19_strm0_ready         ( pe21__std__lane19_strm0_ready      ),      
               .std__pe21__lane19_strm0_cntl          ( std__pe21__lane19_strm0_cntl       ),      
               .std__pe21__lane19_strm0_data          ( std__pe21__lane19_strm0_data       ),      
               .std__pe21__lane19_strm0_data_valid    ( std__pe21__lane19_strm0_data_valid ),      
               .std__pe21__lane19_strm0_data_mask     ( std__pe21__lane19_strm0_data_mask  ),      

               .pe21__std__lane19_strm1_ready         ( pe21__std__lane19_strm1_ready      ),      
               .std__pe21__lane19_strm1_cntl          ( std__pe21__lane19_strm1_cntl       ),      
               .std__pe21__lane19_strm1_data          ( std__pe21__lane19_strm1_data       ),      
               .std__pe21__lane19_strm1_data_valid    ( std__pe21__lane19_strm1_data_valid ),      
               .std__pe21__lane19_strm1_data_mask     ( std__pe21__lane19_strm1_data_mask  ),      

               // PE 21, Lane 20                 
               .pe21__std__lane20_strm0_ready         ( pe21__std__lane20_strm0_ready      ),      
               .std__pe21__lane20_strm0_cntl          ( std__pe21__lane20_strm0_cntl       ),      
               .std__pe21__lane20_strm0_data          ( std__pe21__lane20_strm0_data       ),      
               .std__pe21__lane20_strm0_data_valid    ( std__pe21__lane20_strm0_data_valid ),      
               .std__pe21__lane20_strm0_data_mask     ( std__pe21__lane20_strm0_data_mask  ),      

               .pe21__std__lane20_strm1_ready         ( pe21__std__lane20_strm1_ready      ),      
               .std__pe21__lane20_strm1_cntl          ( std__pe21__lane20_strm1_cntl       ),      
               .std__pe21__lane20_strm1_data          ( std__pe21__lane20_strm1_data       ),      
               .std__pe21__lane20_strm1_data_valid    ( std__pe21__lane20_strm1_data_valid ),      
               .std__pe21__lane20_strm1_data_mask     ( std__pe21__lane20_strm1_data_mask  ),      

               // PE 21, Lane 21                 
               .pe21__std__lane21_strm0_ready         ( pe21__std__lane21_strm0_ready      ),      
               .std__pe21__lane21_strm0_cntl          ( std__pe21__lane21_strm0_cntl       ),      
               .std__pe21__lane21_strm0_data          ( std__pe21__lane21_strm0_data       ),      
               .std__pe21__lane21_strm0_data_valid    ( std__pe21__lane21_strm0_data_valid ),      
               .std__pe21__lane21_strm0_data_mask     ( std__pe21__lane21_strm0_data_mask  ),      

               .pe21__std__lane21_strm1_ready         ( pe21__std__lane21_strm1_ready      ),      
               .std__pe21__lane21_strm1_cntl          ( std__pe21__lane21_strm1_cntl       ),      
               .std__pe21__lane21_strm1_data          ( std__pe21__lane21_strm1_data       ),      
               .std__pe21__lane21_strm1_data_valid    ( std__pe21__lane21_strm1_data_valid ),      
               .std__pe21__lane21_strm1_data_mask     ( std__pe21__lane21_strm1_data_mask  ),      

               // PE 21, Lane 22                 
               .pe21__std__lane22_strm0_ready         ( pe21__std__lane22_strm0_ready      ),      
               .std__pe21__lane22_strm0_cntl          ( std__pe21__lane22_strm0_cntl       ),      
               .std__pe21__lane22_strm0_data          ( std__pe21__lane22_strm0_data       ),      
               .std__pe21__lane22_strm0_data_valid    ( std__pe21__lane22_strm0_data_valid ),      
               .std__pe21__lane22_strm0_data_mask     ( std__pe21__lane22_strm0_data_mask  ),      

               .pe21__std__lane22_strm1_ready         ( pe21__std__lane22_strm1_ready      ),      
               .std__pe21__lane22_strm1_cntl          ( std__pe21__lane22_strm1_cntl       ),      
               .std__pe21__lane22_strm1_data          ( std__pe21__lane22_strm1_data       ),      
               .std__pe21__lane22_strm1_data_valid    ( std__pe21__lane22_strm1_data_valid ),      
               .std__pe21__lane22_strm1_data_mask     ( std__pe21__lane22_strm1_data_mask  ),      

               // PE 21, Lane 23                 
               .pe21__std__lane23_strm0_ready         ( pe21__std__lane23_strm0_ready      ),      
               .std__pe21__lane23_strm0_cntl          ( std__pe21__lane23_strm0_cntl       ),      
               .std__pe21__lane23_strm0_data          ( std__pe21__lane23_strm0_data       ),      
               .std__pe21__lane23_strm0_data_valid    ( std__pe21__lane23_strm0_data_valid ),      
               .std__pe21__lane23_strm0_data_mask     ( std__pe21__lane23_strm0_data_mask  ),      

               .pe21__std__lane23_strm1_ready         ( pe21__std__lane23_strm1_ready      ),      
               .std__pe21__lane23_strm1_cntl          ( std__pe21__lane23_strm1_cntl       ),      
               .std__pe21__lane23_strm1_data          ( std__pe21__lane23_strm1_data       ),      
               .std__pe21__lane23_strm1_data_valid    ( std__pe21__lane23_strm1_data_valid ),      
               .std__pe21__lane23_strm1_data_mask     ( std__pe21__lane23_strm1_data_mask  ),      

               // PE 21, Lane 24                 
               .pe21__std__lane24_strm0_ready         ( pe21__std__lane24_strm0_ready      ),      
               .std__pe21__lane24_strm0_cntl          ( std__pe21__lane24_strm0_cntl       ),      
               .std__pe21__lane24_strm0_data          ( std__pe21__lane24_strm0_data       ),      
               .std__pe21__lane24_strm0_data_valid    ( std__pe21__lane24_strm0_data_valid ),      
               .std__pe21__lane24_strm0_data_mask     ( std__pe21__lane24_strm0_data_mask  ),      

               .pe21__std__lane24_strm1_ready         ( pe21__std__lane24_strm1_ready      ),      
               .std__pe21__lane24_strm1_cntl          ( std__pe21__lane24_strm1_cntl       ),      
               .std__pe21__lane24_strm1_data          ( std__pe21__lane24_strm1_data       ),      
               .std__pe21__lane24_strm1_data_valid    ( std__pe21__lane24_strm1_data_valid ),      
               .std__pe21__lane24_strm1_data_mask     ( std__pe21__lane24_strm1_data_mask  ),      

               // PE 21, Lane 25                 
               .pe21__std__lane25_strm0_ready         ( pe21__std__lane25_strm0_ready      ),      
               .std__pe21__lane25_strm0_cntl          ( std__pe21__lane25_strm0_cntl       ),      
               .std__pe21__lane25_strm0_data          ( std__pe21__lane25_strm0_data       ),      
               .std__pe21__lane25_strm0_data_valid    ( std__pe21__lane25_strm0_data_valid ),      
               .std__pe21__lane25_strm0_data_mask     ( std__pe21__lane25_strm0_data_mask  ),      

               .pe21__std__lane25_strm1_ready         ( pe21__std__lane25_strm1_ready      ),      
               .std__pe21__lane25_strm1_cntl          ( std__pe21__lane25_strm1_cntl       ),      
               .std__pe21__lane25_strm1_data          ( std__pe21__lane25_strm1_data       ),      
               .std__pe21__lane25_strm1_data_valid    ( std__pe21__lane25_strm1_data_valid ),      
               .std__pe21__lane25_strm1_data_mask     ( std__pe21__lane25_strm1_data_mask  ),      

               // PE 21, Lane 26                 
               .pe21__std__lane26_strm0_ready         ( pe21__std__lane26_strm0_ready      ),      
               .std__pe21__lane26_strm0_cntl          ( std__pe21__lane26_strm0_cntl       ),      
               .std__pe21__lane26_strm0_data          ( std__pe21__lane26_strm0_data       ),      
               .std__pe21__lane26_strm0_data_valid    ( std__pe21__lane26_strm0_data_valid ),      
               .std__pe21__lane26_strm0_data_mask     ( std__pe21__lane26_strm0_data_mask  ),      

               .pe21__std__lane26_strm1_ready         ( pe21__std__lane26_strm1_ready      ),      
               .std__pe21__lane26_strm1_cntl          ( std__pe21__lane26_strm1_cntl       ),      
               .std__pe21__lane26_strm1_data          ( std__pe21__lane26_strm1_data       ),      
               .std__pe21__lane26_strm1_data_valid    ( std__pe21__lane26_strm1_data_valid ),      
               .std__pe21__lane26_strm1_data_mask     ( std__pe21__lane26_strm1_data_mask  ),      

               // PE 21, Lane 27                 
               .pe21__std__lane27_strm0_ready         ( pe21__std__lane27_strm0_ready      ),      
               .std__pe21__lane27_strm0_cntl          ( std__pe21__lane27_strm0_cntl       ),      
               .std__pe21__lane27_strm0_data          ( std__pe21__lane27_strm0_data       ),      
               .std__pe21__lane27_strm0_data_valid    ( std__pe21__lane27_strm0_data_valid ),      
               .std__pe21__lane27_strm0_data_mask     ( std__pe21__lane27_strm0_data_mask  ),      

               .pe21__std__lane27_strm1_ready         ( pe21__std__lane27_strm1_ready      ),      
               .std__pe21__lane27_strm1_cntl          ( std__pe21__lane27_strm1_cntl       ),      
               .std__pe21__lane27_strm1_data          ( std__pe21__lane27_strm1_data       ),      
               .std__pe21__lane27_strm1_data_valid    ( std__pe21__lane27_strm1_data_valid ),      
               .std__pe21__lane27_strm1_data_mask     ( std__pe21__lane27_strm1_data_mask  ),      

               // PE 21, Lane 28                 
               .pe21__std__lane28_strm0_ready         ( pe21__std__lane28_strm0_ready      ),      
               .std__pe21__lane28_strm0_cntl          ( std__pe21__lane28_strm0_cntl       ),      
               .std__pe21__lane28_strm0_data          ( std__pe21__lane28_strm0_data       ),      
               .std__pe21__lane28_strm0_data_valid    ( std__pe21__lane28_strm0_data_valid ),      
               .std__pe21__lane28_strm0_data_mask     ( std__pe21__lane28_strm0_data_mask  ),      

               .pe21__std__lane28_strm1_ready         ( pe21__std__lane28_strm1_ready      ),      
               .std__pe21__lane28_strm1_cntl          ( std__pe21__lane28_strm1_cntl       ),      
               .std__pe21__lane28_strm1_data          ( std__pe21__lane28_strm1_data       ),      
               .std__pe21__lane28_strm1_data_valid    ( std__pe21__lane28_strm1_data_valid ),      
               .std__pe21__lane28_strm1_data_mask     ( std__pe21__lane28_strm1_data_mask  ),      

               // PE 21, Lane 29                 
               .pe21__std__lane29_strm0_ready         ( pe21__std__lane29_strm0_ready      ),      
               .std__pe21__lane29_strm0_cntl          ( std__pe21__lane29_strm0_cntl       ),      
               .std__pe21__lane29_strm0_data          ( std__pe21__lane29_strm0_data       ),      
               .std__pe21__lane29_strm0_data_valid    ( std__pe21__lane29_strm0_data_valid ),      
               .std__pe21__lane29_strm0_data_mask     ( std__pe21__lane29_strm0_data_mask  ),      

               .pe21__std__lane29_strm1_ready         ( pe21__std__lane29_strm1_ready      ),      
               .std__pe21__lane29_strm1_cntl          ( std__pe21__lane29_strm1_cntl       ),      
               .std__pe21__lane29_strm1_data          ( std__pe21__lane29_strm1_data       ),      
               .std__pe21__lane29_strm1_data_valid    ( std__pe21__lane29_strm1_data_valid ),      
               .std__pe21__lane29_strm1_data_mask     ( std__pe21__lane29_strm1_data_mask  ),      

               // PE 21, Lane 30                 
               .pe21__std__lane30_strm0_ready         ( pe21__std__lane30_strm0_ready      ),      
               .std__pe21__lane30_strm0_cntl          ( std__pe21__lane30_strm0_cntl       ),      
               .std__pe21__lane30_strm0_data          ( std__pe21__lane30_strm0_data       ),      
               .std__pe21__lane30_strm0_data_valid    ( std__pe21__lane30_strm0_data_valid ),      
               .std__pe21__lane30_strm0_data_mask     ( std__pe21__lane30_strm0_data_mask  ),      

               .pe21__std__lane30_strm1_ready         ( pe21__std__lane30_strm1_ready      ),      
               .std__pe21__lane30_strm1_cntl          ( std__pe21__lane30_strm1_cntl       ),      
               .std__pe21__lane30_strm1_data          ( std__pe21__lane30_strm1_data       ),      
               .std__pe21__lane30_strm1_data_valid    ( std__pe21__lane30_strm1_data_valid ),      
               .std__pe21__lane30_strm1_data_mask     ( std__pe21__lane30_strm1_data_mask  ),      

               // PE 21, Lane 31                 
               .pe21__std__lane31_strm0_ready         ( pe21__std__lane31_strm0_ready      ),      
               .std__pe21__lane31_strm0_cntl          ( std__pe21__lane31_strm0_cntl       ),      
               .std__pe21__lane31_strm0_data          ( std__pe21__lane31_strm0_data       ),      
               .std__pe21__lane31_strm0_data_valid    ( std__pe21__lane31_strm0_data_valid ),      
               .std__pe21__lane31_strm0_data_mask     ( std__pe21__lane31_strm0_data_mask  ),      

               .pe21__std__lane31_strm1_ready         ( pe21__std__lane31_strm1_ready      ),      
               .std__pe21__lane31_strm1_cntl          ( std__pe21__lane31_strm1_cntl       ),      
               .std__pe21__lane31_strm1_data          ( std__pe21__lane31_strm1_data       ),      
               .std__pe21__lane31_strm1_data_valid    ( std__pe21__lane31_strm1_data_valid ),      
               .std__pe21__lane31_strm1_data_mask     ( std__pe21__lane31_strm1_data_mask  ),      

               // PE 22, Lane 0                 
               .pe22__std__lane0_strm0_ready         ( pe22__std__lane0_strm0_ready      ),      
               .std__pe22__lane0_strm0_cntl          ( std__pe22__lane0_strm0_cntl       ),      
               .std__pe22__lane0_strm0_data          ( std__pe22__lane0_strm0_data       ),      
               .std__pe22__lane0_strm0_data_valid    ( std__pe22__lane0_strm0_data_valid ),      
               .std__pe22__lane0_strm0_data_mask     ( std__pe22__lane0_strm0_data_mask  ),      

               .pe22__std__lane0_strm1_ready         ( pe22__std__lane0_strm1_ready      ),      
               .std__pe22__lane0_strm1_cntl          ( std__pe22__lane0_strm1_cntl       ),      
               .std__pe22__lane0_strm1_data          ( std__pe22__lane0_strm1_data       ),      
               .std__pe22__lane0_strm1_data_valid    ( std__pe22__lane0_strm1_data_valid ),      
               .std__pe22__lane0_strm1_data_mask     ( std__pe22__lane0_strm1_data_mask  ),      

               // PE 22, Lane 1                 
               .pe22__std__lane1_strm0_ready         ( pe22__std__lane1_strm0_ready      ),      
               .std__pe22__lane1_strm0_cntl          ( std__pe22__lane1_strm0_cntl       ),      
               .std__pe22__lane1_strm0_data          ( std__pe22__lane1_strm0_data       ),      
               .std__pe22__lane1_strm0_data_valid    ( std__pe22__lane1_strm0_data_valid ),      
               .std__pe22__lane1_strm0_data_mask     ( std__pe22__lane1_strm0_data_mask  ),      

               .pe22__std__lane1_strm1_ready         ( pe22__std__lane1_strm1_ready      ),      
               .std__pe22__lane1_strm1_cntl          ( std__pe22__lane1_strm1_cntl       ),      
               .std__pe22__lane1_strm1_data          ( std__pe22__lane1_strm1_data       ),      
               .std__pe22__lane1_strm1_data_valid    ( std__pe22__lane1_strm1_data_valid ),      
               .std__pe22__lane1_strm1_data_mask     ( std__pe22__lane1_strm1_data_mask  ),      

               // PE 22, Lane 2                 
               .pe22__std__lane2_strm0_ready         ( pe22__std__lane2_strm0_ready      ),      
               .std__pe22__lane2_strm0_cntl          ( std__pe22__lane2_strm0_cntl       ),      
               .std__pe22__lane2_strm0_data          ( std__pe22__lane2_strm0_data       ),      
               .std__pe22__lane2_strm0_data_valid    ( std__pe22__lane2_strm0_data_valid ),      
               .std__pe22__lane2_strm0_data_mask     ( std__pe22__lane2_strm0_data_mask  ),      

               .pe22__std__lane2_strm1_ready         ( pe22__std__lane2_strm1_ready      ),      
               .std__pe22__lane2_strm1_cntl          ( std__pe22__lane2_strm1_cntl       ),      
               .std__pe22__lane2_strm1_data          ( std__pe22__lane2_strm1_data       ),      
               .std__pe22__lane2_strm1_data_valid    ( std__pe22__lane2_strm1_data_valid ),      
               .std__pe22__lane2_strm1_data_mask     ( std__pe22__lane2_strm1_data_mask  ),      

               // PE 22, Lane 3                 
               .pe22__std__lane3_strm0_ready         ( pe22__std__lane3_strm0_ready      ),      
               .std__pe22__lane3_strm0_cntl          ( std__pe22__lane3_strm0_cntl       ),      
               .std__pe22__lane3_strm0_data          ( std__pe22__lane3_strm0_data       ),      
               .std__pe22__lane3_strm0_data_valid    ( std__pe22__lane3_strm0_data_valid ),      
               .std__pe22__lane3_strm0_data_mask     ( std__pe22__lane3_strm0_data_mask  ),      

               .pe22__std__lane3_strm1_ready         ( pe22__std__lane3_strm1_ready      ),      
               .std__pe22__lane3_strm1_cntl          ( std__pe22__lane3_strm1_cntl       ),      
               .std__pe22__lane3_strm1_data          ( std__pe22__lane3_strm1_data       ),      
               .std__pe22__lane3_strm1_data_valid    ( std__pe22__lane3_strm1_data_valid ),      
               .std__pe22__lane3_strm1_data_mask     ( std__pe22__lane3_strm1_data_mask  ),      

               // PE 22, Lane 4                 
               .pe22__std__lane4_strm0_ready         ( pe22__std__lane4_strm0_ready      ),      
               .std__pe22__lane4_strm0_cntl          ( std__pe22__lane4_strm0_cntl       ),      
               .std__pe22__lane4_strm0_data          ( std__pe22__lane4_strm0_data       ),      
               .std__pe22__lane4_strm0_data_valid    ( std__pe22__lane4_strm0_data_valid ),      
               .std__pe22__lane4_strm0_data_mask     ( std__pe22__lane4_strm0_data_mask  ),      

               .pe22__std__lane4_strm1_ready         ( pe22__std__lane4_strm1_ready      ),      
               .std__pe22__lane4_strm1_cntl          ( std__pe22__lane4_strm1_cntl       ),      
               .std__pe22__lane4_strm1_data          ( std__pe22__lane4_strm1_data       ),      
               .std__pe22__lane4_strm1_data_valid    ( std__pe22__lane4_strm1_data_valid ),      
               .std__pe22__lane4_strm1_data_mask     ( std__pe22__lane4_strm1_data_mask  ),      

               // PE 22, Lane 5                 
               .pe22__std__lane5_strm0_ready         ( pe22__std__lane5_strm0_ready      ),      
               .std__pe22__lane5_strm0_cntl          ( std__pe22__lane5_strm0_cntl       ),      
               .std__pe22__lane5_strm0_data          ( std__pe22__lane5_strm0_data       ),      
               .std__pe22__lane5_strm0_data_valid    ( std__pe22__lane5_strm0_data_valid ),      
               .std__pe22__lane5_strm0_data_mask     ( std__pe22__lane5_strm0_data_mask  ),      

               .pe22__std__lane5_strm1_ready         ( pe22__std__lane5_strm1_ready      ),      
               .std__pe22__lane5_strm1_cntl          ( std__pe22__lane5_strm1_cntl       ),      
               .std__pe22__lane5_strm1_data          ( std__pe22__lane5_strm1_data       ),      
               .std__pe22__lane5_strm1_data_valid    ( std__pe22__lane5_strm1_data_valid ),      
               .std__pe22__lane5_strm1_data_mask     ( std__pe22__lane5_strm1_data_mask  ),      

               // PE 22, Lane 6                 
               .pe22__std__lane6_strm0_ready         ( pe22__std__lane6_strm0_ready      ),      
               .std__pe22__lane6_strm0_cntl          ( std__pe22__lane6_strm0_cntl       ),      
               .std__pe22__lane6_strm0_data          ( std__pe22__lane6_strm0_data       ),      
               .std__pe22__lane6_strm0_data_valid    ( std__pe22__lane6_strm0_data_valid ),      
               .std__pe22__lane6_strm0_data_mask     ( std__pe22__lane6_strm0_data_mask  ),      

               .pe22__std__lane6_strm1_ready         ( pe22__std__lane6_strm1_ready      ),      
               .std__pe22__lane6_strm1_cntl          ( std__pe22__lane6_strm1_cntl       ),      
               .std__pe22__lane6_strm1_data          ( std__pe22__lane6_strm1_data       ),      
               .std__pe22__lane6_strm1_data_valid    ( std__pe22__lane6_strm1_data_valid ),      
               .std__pe22__lane6_strm1_data_mask     ( std__pe22__lane6_strm1_data_mask  ),      

               // PE 22, Lane 7                 
               .pe22__std__lane7_strm0_ready         ( pe22__std__lane7_strm0_ready      ),      
               .std__pe22__lane7_strm0_cntl          ( std__pe22__lane7_strm0_cntl       ),      
               .std__pe22__lane7_strm0_data          ( std__pe22__lane7_strm0_data       ),      
               .std__pe22__lane7_strm0_data_valid    ( std__pe22__lane7_strm0_data_valid ),      
               .std__pe22__lane7_strm0_data_mask     ( std__pe22__lane7_strm0_data_mask  ),      

               .pe22__std__lane7_strm1_ready         ( pe22__std__lane7_strm1_ready      ),      
               .std__pe22__lane7_strm1_cntl          ( std__pe22__lane7_strm1_cntl       ),      
               .std__pe22__lane7_strm1_data          ( std__pe22__lane7_strm1_data       ),      
               .std__pe22__lane7_strm1_data_valid    ( std__pe22__lane7_strm1_data_valid ),      
               .std__pe22__lane7_strm1_data_mask     ( std__pe22__lane7_strm1_data_mask  ),      

               // PE 22, Lane 8                 
               .pe22__std__lane8_strm0_ready         ( pe22__std__lane8_strm0_ready      ),      
               .std__pe22__lane8_strm0_cntl          ( std__pe22__lane8_strm0_cntl       ),      
               .std__pe22__lane8_strm0_data          ( std__pe22__lane8_strm0_data       ),      
               .std__pe22__lane8_strm0_data_valid    ( std__pe22__lane8_strm0_data_valid ),      
               .std__pe22__lane8_strm0_data_mask     ( std__pe22__lane8_strm0_data_mask  ),      

               .pe22__std__lane8_strm1_ready         ( pe22__std__lane8_strm1_ready      ),      
               .std__pe22__lane8_strm1_cntl          ( std__pe22__lane8_strm1_cntl       ),      
               .std__pe22__lane8_strm1_data          ( std__pe22__lane8_strm1_data       ),      
               .std__pe22__lane8_strm1_data_valid    ( std__pe22__lane8_strm1_data_valid ),      
               .std__pe22__lane8_strm1_data_mask     ( std__pe22__lane8_strm1_data_mask  ),      

               // PE 22, Lane 9                 
               .pe22__std__lane9_strm0_ready         ( pe22__std__lane9_strm0_ready      ),      
               .std__pe22__lane9_strm0_cntl          ( std__pe22__lane9_strm0_cntl       ),      
               .std__pe22__lane9_strm0_data          ( std__pe22__lane9_strm0_data       ),      
               .std__pe22__lane9_strm0_data_valid    ( std__pe22__lane9_strm0_data_valid ),      
               .std__pe22__lane9_strm0_data_mask     ( std__pe22__lane9_strm0_data_mask  ),      

               .pe22__std__lane9_strm1_ready         ( pe22__std__lane9_strm1_ready      ),      
               .std__pe22__lane9_strm1_cntl          ( std__pe22__lane9_strm1_cntl       ),      
               .std__pe22__lane9_strm1_data          ( std__pe22__lane9_strm1_data       ),      
               .std__pe22__lane9_strm1_data_valid    ( std__pe22__lane9_strm1_data_valid ),      
               .std__pe22__lane9_strm1_data_mask     ( std__pe22__lane9_strm1_data_mask  ),      

               // PE 22, Lane 10                 
               .pe22__std__lane10_strm0_ready         ( pe22__std__lane10_strm0_ready      ),      
               .std__pe22__lane10_strm0_cntl          ( std__pe22__lane10_strm0_cntl       ),      
               .std__pe22__lane10_strm0_data          ( std__pe22__lane10_strm0_data       ),      
               .std__pe22__lane10_strm0_data_valid    ( std__pe22__lane10_strm0_data_valid ),      
               .std__pe22__lane10_strm0_data_mask     ( std__pe22__lane10_strm0_data_mask  ),      

               .pe22__std__lane10_strm1_ready         ( pe22__std__lane10_strm1_ready      ),      
               .std__pe22__lane10_strm1_cntl          ( std__pe22__lane10_strm1_cntl       ),      
               .std__pe22__lane10_strm1_data          ( std__pe22__lane10_strm1_data       ),      
               .std__pe22__lane10_strm1_data_valid    ( std__pe22__lane10_strm1_data_valid ),      
               .std__pe22__lane10_strm1_data_mask     ( std__pe22__lane10_strm1_data_mask  ),      

               // PE 22, Lane 11                 
               .pe22__std__lane11_strm0_ready         ( pe22__std__lane11_strm0_ready      ),      
               .std__pe22__lane11_strm0_cntl          ( std__pe22__lane11_strm0_cntl       ),      
               .std__pe22__lane11_strm0_data          ( std__pe22__lane11_strm0_data       ),      
               .std__pe22__lane11_strm0_data_valid    ( std__pe22__lane11_strm0_data_valid ),      
               .std__pe22__lane11_strm0_data_mask     ( std__pe22__lane11_strm0_data_mask  ),      

               .pe22__std__lane11_strm1_ready         ( pe22__std__lane11_strm1_ready      ),      
               .std__pe22__lane11_strm1_cntl          ( std__pe22__lane11_strm1_cntl       ),      
               .std__pe22__lane11_strm1_data          ( std__pe22__lane11_strm1_data       ),      
               .std__pe22__lane11_strm1_data_valid    ( std__pe22__lane11_strm1_data_valid ),      
               .std__pe22__lane11_strm1_data_mask     ( std__pe22__lane11_strm1_data_mask  ),      

               // PE 22, Lane 12                 
               .pe22__std__lane12_strm0_ready         ( pe22__std__lane12_strm0_ready      ),      
               .std__pe22__lane12_strm0_cntl          ( std__pe22__lane12_strm0_cntl       ),      
               .std__pe22__lane12_strm0_data          ( std__pe22__lane12_strm0_data       ),      
               .std__pe22__lane12_strm0_data_valid    ( std__pe22__lane12_strm0_data_valid ),      
               .std__pe22__lane12_strm0_data_mask     ( std__pe22__lane12_strm0_data_mask  ),      

               .pe22__std__lane12_strm1_ready         ( pe22__std__lane12_strm1_ready      ),      
               .std__pe22__lane12_strm1_cntl          ( std__pe22__lane12_strm1_cntl       ),      
               .std__pe22__lane12_strm1_data          ( std__pe22__lane12_strm1_data       ),      
               .std__pe22__lane12_strm1_data_valid    ( std__pe22__lane12_strm1_data_valid ),      
               .std__pe22__lane12_strm1_data_mask     ( std__pe22__lane12_strm1_data_mask  ),      

               // PE 22, Lane 13                 
               .pe22__std__lane13_strm0_ready         ( pe22__std__lane13_strm0_ready      ),      
               .std__pe22__lane13_strm0_cntl          ( std__pe22__lane13_strm0_cntl       ),      
               .std__pe22__lane13_strm0_data          ( std__pe22__lane13_strm0_data       ),      
               .std__pe22__lane13_strm0_data_valid    ( std__pe22__lane13_strm0_data_valid ),      
               .std__pe22__lane13_strm0_data_mask     ( std__pe22__lane13_strm0_data_mask  ),      

               .pe22__std__lane13_strm1_ready         ( pe22__std__lane13_strm1_ready      ),      
               .std__pe22__lane13_strm1_cntl          ( std__pe22__lane13_strm1_cntl       ),      
               .std__pe22__lane13_strm1_data          ( std__pe22__lane13_strm1_data       ),      
               .std__pe22__lane13_strm1_data_valid    ( std__pe22__lane13_strm1_data_valid ),      
               .std__pe22__lane13_strm1_data_mask     ( std__pe22__lane13_strm1_data_mask  ),      

               // PE 22, Lane 14                 
               .pe22__std__lane14_strm0_ready         ( pe22__std__lane14_strm0_ready      ),      
               .std__pe22__lane14_strm0_cntl          ( std__pe22__lane14_strm0_cntl       ),      
               .std__pe22__lane14_strm0_data          ( std__pe22__lane14_strm0_data       ),      
               .std__pe22__lane14_strm0_data_valid    ( std__pe22__lane14_strm0_data_valid ),      
               .std__pe22__lane14_strm0_data_mask     ( std__pe22__lane14_strm0_data_mask  ),      

               .pe22__std__lane14_strm1_ready         ( pe22__std__lane14_strm1_ready      ),      
               .std__pe22__lane14_strm1_cntl          ( std__pe22__lane14_strm1_cntl       ),      
               .std__pe22__lane14_strm1_data          ( std__pe22__lane14_strm1_data       ),      
               .std__pe22__lane14_strm1_data_valid    ( std__pe22__lane14_strm1_data_valid ),      
               .std__pe22__lane14_strm1_data_mask     ( std__pe22__lane14_strm1_data_mask  ),      

               // PE 22, Lane 15                 
               .pe22__std__lane15_strm0_ready         ( pe22__std__lane15_strm0_ready      ),      
               .std__pe22__lane15_strm0_cntl          ( std__pe22__lane15_strm0_cntl       ),      
               .std__pe22__lane15_strm0_data          ( std__pe22__lane15_strm0_data       ),      
               .std__pe22__lane15_strm0_data_valid    ( std__pe22__lane15_strm0_data_valid ),      
               .std__pe22__lane15_strm0_data_mask     ( std__pe22__lane15_strm0_data_mask  ),      

               .pe22__std__lane15_strm1_ready         ( pe22__std__lane15_strm1_ready      ),      
               .std__pe22__lane15_strm1_cntl          ( std__pe22__lane15_strm1_cntl       ),      
               .std__pe22__lane15_strm1_data          ( std__pe22__lane15_strm1_data       ),      
               .std__pe22__lane15_strm1_data_valid    ( std__pe22__lane15_strm1_data_valid ),      
               .std__pe22__lane15_strm1_data_mask     ( std__pe22__lane15_strm1_data_mask  ),      

               // PE 22, Lane 16                 
               .pe22__std__lane16_strm0_ready         ( pe22__std__lane16_strm0_ready      ),      
               .std__pe22__lane16_strm0_cntl          ( std__pe22__lane16_strm0_cntl       ),      
               .std__pe22__lane16_strm0_data          ( std__pe22__lane16_strm0_data       ),      
               .std__pe22__lane16_strm0_data_valid    ( std__pe22__lane16_strm0_data_valid ),      
               .std__pe22__lane16_strm0_data_mask     ( std__pe22__lane16_strm0_data_mask  ),      

               .pe22__std__lane16_strm1_ready         ( pe22__std__lane16_strm1_ready      ),      
               .std__pe22__lane16_strm1_cntl          ( std__pe22__lane16_strm1_cntl       ),      
               .std__pe22__lane16_strm1_data          ( std__pe22__lane16_strm1_data       ),      
               .std__pe22__lane16_strm1_data_valid    ( std__pe22__lane16_strm1_data_valid ),      
               .std__pe22__lane16_strm1_data_mask     ( std__pe22__lane16_strm1_data_mask  ),      

               // PE 22, Lane 17                 
               .pe22__std__lane17_strm0_ready         ( pe22__std__lane17_strm0_ready      ),      
               .std__pe22__lane17_strm0_cntl          ( std__pe22__lane17_strm0_cntl       ),      
               .std__pe22__lane17_strm0_data          ( std__pe22__lane17_strm0_data       ),      
               .std__pe22__lane17_strm0_data_valid    ( std__pe22__lane17_strm0_data_valid ),      
               .std__pe22__lane17_strm0_data_mask     ( std__pe22__lane17_strm0_data_mask  ),      

               .pe22__std__lane17_strm1_ready         ( pe22__std__lane17_strm1_ready      ),      
               .std__pe22__lane17_strm1_cntl          ( std__pe22__lane17_strm1_cntl       ),      
               .std__pe22__lane17_strm1_data          ( std__pe22__lane17_strm1_data       ),      
               .std__pe22__lane17_strm1_data_valid    ( std__pe22__lane17_strm1_data_valid ),      
               .std__pe22__lane17_strm1_data_mask     ( std__pe22__lane17_strm1_data_mask  ),      

               // PE 22, Lane 18                 
               .pe22__std__lane18_strm0_ready         ( pe22__std__lane18_strm0_ready      ),      
               .std__pe22__lane18_strm0_cntl          ( std__pe22__lane18_strm0_cntl       ),      
               .std__pe22__lane18_strm0_data          ( std__pe22__lane18_strm0_data       ),      
               .std__pe22__lane18_strm0_data_valid    ( std__pe22__lane18_strm0_data_valid ),      
               .std__pe22__lane18_strm0_data_mask     ( std__pe22__lane18_strm0_data_mask  ),      

               .pe22__std__lane18_strm1_ready         ( pe22__std__lane18_strm1_ready      ),      
               .std__pe22__lane18_strm1_cntl          ( std__pe22__lane18_strm1_cntl       ),      
               .std__pe22__lane18_strm1_data          ( std__pe22__lane18_strm1_data       ),      
               .std__pe22__lane18_strm1_data_valid    ( std__pe22__lane18_strm1_data_valid ),      
               .std__pe22__lane18_strm1_data_mask     ( std__pe22__lane18_strm1_data_mask  ),      

               // PE 22, Lane 19                 
               .pe22__std__lane19_strm0_ready         ( pe22__std__lane19_strm0_ready      ),      
               .std__pe22__lane19_strm0_cntl          ( std__pe22__lane19_strm0_cntl       ),      
               .std__pe22__lane19_strm0_data          ( std__pe22__lane19_strm0_data       ),      
               .std__pe22__lane19_strm0_data_valid    ( std__pe22__lane19_strm0_data_valid ),      
               .std__pe22__lane19_strm0_data_mask     ( std__pe22__lane19_strm0_data_mask  ),      

               .pe22__std__lane19_strm1_ready         ( pe22__std__lane19_strm1_ready      ),      
               .std__pe22__lane19_strm1_cntl          ( std__pe22__lane19_strm1_cntl       ),      
               .std__pe22__lane19_strm1_data          ( std__pe22__lane19_strm1_data       ),      
               .std__pe22__lane19_strm1_data_valid    ( std__pe22__lane19_strm1_data_valid ),      
               .std__pe22__lane19_strm1_data_mask     ( std__pe22__lane19_strm1_data_mask  ),      

               // PE 22, Lane 20                 
               .pe22__std__lane20_strm0_ready         ( pe22__std__lane20_strm0_ready      ),      
               .std__pe22__lane20_strm0_cntl          ( std__pe22__lane20_strm0_cntl       ),      
               .std__pe22__lane20_strm0_data          ( std__pe22__lane20_strm0_data       ),      
               .std__pe22__lane20_strm0_data_valid    ( std__pe22__lane20_strm0_data_valid ),      
               .std__pe22__lane20_strm0_data_mask     ( std__pe22__lane20_strm0_data_mask  ),      

               .pe22__std__lane20_strm1_ready         ( pe22__std__lane20_strm1_ready      ),      
               .std__pe22__lane20_strm1_cntl          ( std__pe22__lane20_strm1_cntl       ),      
               .std__pe22__lane20_strm1_data          ( std__pe22__lane20_strm1_data       ),      
               .std__pe22__lane20_strm1_data_valid    ( std__pe22__lane20_strm1_data_valid ),      
               .std__pe22__lane20_strm1_data_mask     ( std__pe22__lane20_strm1_data_mask  ),      

               // PE 22, Lane 21                 
               .pe22__std__lane21_strm0_ready         ( pe22__std__lane21_strm0_ready      ),      
               .std__pe22__lane21_strm0_cntl          ( std__pe22__lane21_strm0_cntl       ),      
               .std__pe22__lane21_strm0_data          ( std__pe22__lane21_strm0_data       ),      
               .std__pe22__lane21_strm0_data_valid    ( std__pe22__lane21_strm0_data_valid ),      
               .std__pe22__lane21_strm0_data_mask     ( std__pe22__lane21_strm0_data_mask  ),      

               .pe22__std__lane21_strm1_ready         ( pe22__std__lane21_strm1_ready      ),      
               .std__pe22__lane21_strm1_cntl          ( std__pe22__lane21_strm1_cntl       ),      
               .std__pe22__lane21_strm1_data          ( std__pe22__lane21_strm1_data       ),      
               .std__pe22__lane21_strm1_data_valid    ( std__pe22__lane21_strm1_data_valid ),      
               .std__pe22__lane21_strm1_data_mask     ( std__pe22__lane21_strm1_data_mask  ),      

               // PE 22, Lane 22                 
               .pe22__std__lane22_strm0_ready         ( pe22__std__lane22_strm0_ready      ),      
               .std__pe22__lane22_strm0_cntl          ( std__pe22__lane22_strm0_cntl       ),      
               .std__pe22__lane22_strm0_data          ( std__pe22__lane22_strm0_data       ),      
               .std__pe22__lane22_strm0_data_valid    ( std__pe22__lane22_strm0_data_valid ),      
               .std__pe22__lane22_strm0_data_mask     ( std__pe22__lane22_strm0_data_mask  ),      

               .pe22__std__lane22_strm1_ready         ( pe22__std__lane22_strm1_ready      ),      
               .std__pe22__lane22_strm1_cntl          ( std__pe22__lane22_strm1_cntl       ),      
               .std__pe22__lane22_strm1_data          ( std__pe22__lane22_strm1_data       ),      
               .std__pe22__lane22_strm1_data_valid    ( std__pe22__lane22_strm1_data_valid ),      
               .std__pe22__lane22_strm1_data_mask     ( std__pe22__lane22_strm1_data_mask  ),      

               // PE 22, Lane 23                 
               .pe22__std__lane23_strm0_ready         ( pe22__std__lane23_strm0_ready      ),      
               .std__pe22__lane23_strm0_cntl          ( std__pe22__lane23_strm0_cntl       ),      
               .std__pe22__lane23_strm0_data          ( std__pe22__lane23_strm0_data       ),      
               .std__pe22__lane23_strm0_data_valid    ( std__pe22__lane23_strm0_data_valid ),      
               .std__pe22__lane23_strm0_data_mask     ( std__pe22__lane23_strm0_data_mask  ),      

               .pe22__std__lane23_strm1_ready         ( pe22__std__lane23_strm1_ready      ),      
               .std__pe22__lane23_strm1_cntl          ( std__pe22__lane23_strm1_cntl       ),      
               .std__pe22__lane23_strm1_data          ( std__pe22__lane23_strm1_data       ),      
               .std__pe22__lane23_strm1_data_valid    ( std__pe22__lane23_strm1_data_valid ),      
               .std__pe22__lane23_strm1_data_mask     ( std__pe22__lane23_strm1_data_mask  ),      

               // PE 22, Lane 24                 
               .pe22__std__lane24_strm0_ready         ( pe22__std__lane24_strm0_ready      ),      
               .std__pe22__lane24_strm0_cntl          ( std__pe22__lane24_strm0_cntl       ),      
               .std__pe22__lane24_strm0_data          ( std__pe22__lane24_strm0_data       ),      
               .std__pe22__lane24_strm0_data_valid    ( std__pe22__lane24_strm0_data_valid ),      
               .std__pe22__lane24_strm0_data_mask     ( std__pe22__lane24_strm0_data_mask  ),      

               .pe22__std__lane24_strm1_ready         ( pe22__std__lane24_strm1_ready      ),      
               .std__pe22__lane24_strm1_cntl          ( std__pe22__lane24_strm1_cntl       ),      
               .std__pe22__lane24_strm1_data          ( std__pe22__lane24_strm1_data       ),      
               .std__pe22__lane24_strm1_data_valid    ( std__pe22__lane24_strm1_data_valid ),      
               .std__pe22__lane24_strm1_data_mask     ( std__pe22__lane24_strm1_data_mask  ),      

               // PE 22, Lane 25                 
               .pe22__std__lane25_strm0_ready         ( pe22__std__lane25_strm0_ready      ),      
               .std__pe22__lane25_strm0_cntl          ( std__pe22__lane25_strm0_cntl       ),      
               .std__pe22__lane25_strm0_data          ( std__pe22__lane25_strm0_data       ),      
               .std__pe22__lane25_strm0_data_valid    ( std__pe22__lane25_strm0_data_valid ),      
               .std__pe22__lane25_strm0_data_mask     ( std__pe22__lane25_strm0_data_mask  ),      

               .pe22__std__lane25_strm1_ready         ( pe22__std__lane25_strm1_ready      ),      
               .std__pe22__lane25_strm1_cntl          ( std__pe22__lane25_strm1_cntl       ),      
               .std__pe22__lane25_strm1_data          ( std__pe22__lane25_strm1_data       ),      
               .std__pe22__lane25_strm1_data_valid    ( std__pe22__lane25_strm1_data_valid ),      
               .std__pe22__lane25_strm1_data_mask     ( std__pe22__lane25_strm1_data_mask  ),      

               // PE 22, Lane 26                 
               .pe22__std__lane26_strm0_ready         ( pe22__std__lane26_strm0_ready      ),      
               .std__pe22__lane26_strm0_cntl          ( std__pe22__lane26_strm0_cntl       ),      
               .std__pe22__lane26_strm0_data          ( std__pe22__lane26_strm0_data       ),      
               .std__pe22__lane26_strm0_data_valid    ( std__pe22__lane26_strm0_data_valid ),      
               .std__pe22__lane26_strm0_data_mask     ( std__pe22__lane26_strm0_data_mask  ),      

               .pe22__std__lane26_strm1_ready         ( pe22__std__lane26_strm1_ready      ),      
               .std__pe22__lane26_strm1_cntl          ( std__pe22__lane26_strm1_cntl       ),      
               .std__pe22__lane26_strm1_data          ( std__pe22__lane26_strm1_data       ),      
               .std__pe22__lane26_strm1_data_valid    ( std__pe22__lane26_strm1_data_valid ),      
               .std__pe22__lane26_strm1_data_mask     ( std__pe22__lane26_strm1_data_mask  ),      

               // PE 22, Lane 27                 
               .pe22__std__lane27_strm0_ready         ( pe22__std__lane27_strm0_ready      ),      
               .std__pe22__lane27_strm0_cntl          ( std__pe22__lane27_strm0_cntl       ),      
               .std__pe22__lane27_strm0_data          ( std__pe22__lane27_strm0_data       ),      
               .std__pe22__lane27_strm0_data_valid    ( std__pe22__lane27_strm0_data_valid ),      
               .std__pe22__lane27_strm0_data_mask     ( std__pe22__lane27_strm0_data_mask  ),      

               .pe22__std__lane27_strm1_ready         ( pe22__std__lane27_strm1_ready      ),      
               .std__pe22__lane27_strm1_cntl          ( std__pe22__lane27_strm1_cntl       ),      
               .std__pe22__lane27_strm1_data          ( std__pe22__lane27_strm1_data       ),      
               .std__pe22__lane27_strm1_data_valid    ( std__pe22__lane27_strm1_data_valid ),      
               .std__pe22__lane27_strm1_data_mask     ( std__pe22__lane27_strm1_data_mask  ),      

               // PE 22, Lane 28                 
               .pe22__std__lane28_strm0_ready         ( pe22__std__lane28_strm0_ready      ),      
               .std__pe22__lane28_strm0_cntl          ( std__pe22__lane28_strm0_cntl       ),      
               .std__pe22__lane28_strm0_data          ( std__pe22__lane28_strm0_data       ),      
               .std__pe22__lane28_strm0_data_valid    ( std__pe22__lane28_strm0_data_valid ),      
               .std__pe22__lane28_strm0_data_mask     ( std__pe22__lane28_strm0_data_mask  ),      

               .pe22__std__lane28_strm1_ready         ( pe22__std__lane28_strm1_ready      ),      
               .std__pe22__lane28_strm1_cntl          ( std__pe22__lane28_strm1_cntl       ),      
               .std__pe22__lane28_strm1_data          ( std__pe22__lane28_strm1_data       ),      
               .std__pe22__lane28_strm1_data_valid    ( std__pe22__lane28_strm1_data_valid ),      
               .std__pe22__lane28_strm1_data_mask     ( std__pe22__lane28_strm1_data_mask  ),      

               // PE 22, Lane 29                 
               .pe22__std__lane29_strm0_ready         ( pe22__std__lane29_strm0_ready      ),      
               .std__pe22__lane29_strm0_cntl          ( std__pe22__lane29_strm0_cntl       ),      
               .std__pe22__lane29_strm0_data          ( std__pe22__lane29_strm0_data       ),      
               .std__pe22__lane29_strm0_data_valid    ( std__pe22__lane29_strm0_data_valid ),      
               .std__pe22__lane29_strm0_data_mask     ( std__pe22__lane29_strm0_data_mask  ),      

               .pe22__std__lane29_strm1_ready         ( pe22__std__lane29_strm1_ready      ),      
               .std__pe22__lane29_strm1_cntl          ( std__pe22__lane29_strm1_cntl       ),      
               .std__pe22__lane29_strm1_data          ( std__pe22__lane29_strm1_data       ),      
               .std__pe22__lane29_strm1_data_valid    ( std__pe22__lane29_strm1_data_valid ),      
               .std__pe22__lane29_strm1_data_mask     ( std__pe22__lane29_strm1_data_mask  ),      

               // PE 22, Lane 30                 
               .pe22__std__lane30_strm0_ready         ( pe22__std__lane30_strm0_ready      ),      
               .std__pe22__lane30_strm0_cntl          ( std__pe22__lane30_strm0_cntl       ),      
               .std__pe22__lane30_strm0_data          ( std__pe22__lane30_strm0_data       ),      
               .std__pe22__lane30_strm0_data_valid    ( std__pe22__lane30_strm0_data_valid ),      
               .std__pe22__lane30_strm0_data_mask     ( std__pe22__lane30_strm0_data_mask  ),      

               .pe22__std__lane30_strm1_ready         ( pe22__std__lane30_strm1_ready      ),      
               .std__pe22__lane30_strm1_cntl          ( std__pe22__lane30_strm1_cntl       ),      
               .std__pe22__lane30_strm1_data          ( std__pe22__lane30_strm1_data       ),      
               .std__pe22__lane30_strm1_data_valid    ( std__pe22__lane30_strm1_data_valid ),      
               .std__pe22__lane30_strm1_data_mask     ( std__pe22__lane30_strm1_data_mask  ),      

               // PE 22, Lane 31                 
               .pe22__std__lane31_strm0_ready         ( pe22__std__lane31_strm0_ready      ),      
               .std__pe22__lane31_strm0_cntl          ( std__pe22__lane31_strm0_cntl       ),      
               .std__pe22__lane31_strm0_data          ( std__pe22__lane31_strm0_data       ),      
               .std__pe22__lane31_strm0_data_valid    ( std__pe22__lane31_strm0_data_valid ),      
               .std__pe22__lane31_strm0_data_mask     ( std__pe22__lane31_strm0_data_mask  ),      

               .pe22__std__lane31_strm1_ready         ( pe22__std__lane31_strm1_ready      ),      
               .std__pe22__lane31_strm1_cntl          ( std__pe22__lane31_strm1_cntl       ),      
               .std__pe22__lane31_strm1_data          ( std__pe22__lane31_strm1_data       ),      
               .std__pe22__lane31_strm1_data_valid    ( std__pe22__lane31_strm1_data_valid ),      
               .std__pe22__lane31_strm1_data_mask     ( std__pe22__lane31_strm1_data_mask  ),      

               // PE 23, Lane 0                 
               .pe23__std__lane0_strm0_ready         ( pe23__std__lane0_strm0_ready      ),      
               .std__pe23__lane0_strm0_cntl          ( std__pe23__lane0_strm0_cntl       ),      
               .std__pe23__lane0_strm0_data          ( std__pe23__lane0_strm0_data       ),      
               .std__pe23__lane0_strm0_data_valid    ( std__pe23__lane0_strm0_data_valid ),      
               .std__pe23__lane0_strm0_data_mask     ( std__pe23__lane0_strm0_data_mask  ),      

               .pe23__std__lane0_strm1_ready         ( pe23__std__lane0_strm1_ready      ),      
               .std__pe23__lane0_strm1_cntl          ( std__pe23__lane0_strm1_cntl       ),      
               .std__pe23__lane0_strm1_data          ( std__pe23__lane0_strm1_data       ),      
               .std__pe23__lane0_strm1_data_valid    ( std__pe23__lane0_strm1_data_valid ),      
               .std__pe23__lane0_strm1_data_mask     ( std__pe23__lane0_strm1_data_mask  ),      

               // PE 23, Lane 1                 
               .pe23__std__lane1_strm0_ready         ( pe23__std__lane1_strm0_ready      ),      
               .std__pe23__lane1_strm0_cntl          ( std__pe23__lane1_strm0_cntl       ),      
               .std__pe23__lane1_strm0_data          ( std__pe23__lane1_strm0_data       ),      
               .std__pe23__lane1_strm0_data_valid    ( std__pe23__lane1_strm0_data_valid ),      
               .std__pe23__lane1_strm0_data_mask     ( std__pe23__lane1_strm0_data_mask  ),      

               .pe23__std__lane1_strm1_ready         ( pe23__std__lane1_strm1_ready      ),      
               .std__pe23__lane1_strm1_cntl          ( std__pe23__lane1_strm1_cntl       ),      
               .std__pe23__lane1_strm1_data          ( std__pe23__lane1_strm1_data       ),      
               .std__pe23__lane1_strm1_data_valid    ( std__pe23__lane1_strm1_data_valid ),      
               .std__pe23__lane1_strm1_data_mask     ( std__pe23__lane1_strm1_data_mask  ),      

               // PE 23, Lane 2                 
               .pe23__std__lane2_strm0_ready         ( pe23__std__lane2_strm0_ready      ),      
               .std__pe23__lane2_strm0_cntl          ( std__pe23__lane2_strm0_cntl       ),      
               .std__pe23__lane2_strm0_data          ( std__pe23__lane2_strm0_data       ),      
               .std__pe23__lane2_strm0_data_valid    ( std__pe23__lane2_strm0_data_valid ),      
               .std__pe23__lane2_strm0_data_mask     ( std__pe23__lane2_strm0_data_mask  ),      

               .pe23__std__lane2_strm1_ready         ( pe23__std__lane2_strm1_ready      ),      
               .std__pe23__lane2_strm1_cntl          ( std__pe23__lane2_strm1_cntl       ),      
               .std__pe23__lane2_strm1_data          ( std__pe23__lane2_strm1_data       ),      
               .std__pe23__lane2_strm1_data_valid    ( std__pe23__lane2_strm1_data_valid ),      
               .std__pe23__lane2_strm1_data_mask     ( std__pe23__lane2_strm1_data_mask  ),      

               // PE 23, Lane 3                 
               .pe23__std__lane3_strm0_ready         ( pe23__std__lane3_strm0_ready      ),      
               .std__pe23__lane3_strm0_cntl          ( std__pe23__lane3_strm0_cntl       ),      
               .std__pe23__lane3_strm0_data          ( std__pe23__lane3_strm0_data       ),      
               .std__pe23__lane3_strm0_data_valid    ( std__pe23__lane3_strm0_data_valid ),      
               .std__pe23__lane3_strm0_data_mask     ( std__pe23__lane3_strm0_data_mask  ),      

               .pe23__std__lane3_strm1_ready         ( pe23__std__lane3_strm1_ready      ),      
               .std__pe23__lane3_strm1_cntl          ( std__pe23__lane3_strm1_cntl       ),      
               .std__pe23__lane3_strm1_data          ( std__pe23__lane3_strm1_data       ),      
               .std__pe23__lane3_strm1_data_valid    ( std__pe23__lane3_strm1_data_valid ),      
               .std__pe23__lane3_strm1_data_mask     ( std__pe23__lane3_strm1_data_mask  ),      

               // PE 23, Lane 4                 
               .pe23__std__lane4_strm0_ready         ( pe23__std__lane4_strm0_ready      ),      
               .std__pe23__lane4_strm0_cntl          ( std__pe23__lane4_strm0_cntl       ),      
               .std__pe23__lane4_strm0_data          ( std__pe23__lane4_strm0_data       ),      
               .std__pe23__lane4_strm0_data_valid    ( std__pe23__lane4_strm0_data_valid ),      
               .std__pe23__lane4_strm0_data_mask     ( std__pe23__lane4_strm0_data_mask  ),      

               .pe23__std__lane4_strm1_ready         ( pe23__std__lane4_strm1_ready      ),      
               .std__pe23__lane4_strm1_cntl          ( std__pe23__lane4_strm1_cntl       ),      
               .std__pe23__lane4_strm1_data          ( std__pe23__lane4_strm1_data       ),      
               .std__pe23__lane4_strm1_data_valid    ( std__pe23__lane4_strm1_data_valid ),      
               .std__pe23__lane4_strm1_data_mask     ( std__pe23__lane4_strm1_data_mask  ),      

               // PE 23, Lane 5                 
               .pe23__std__lane5_strm0_ready         ( pe23__std__lane5_strm0_ready      ),      
               .std__pe23__lane5_strm0_cntl          ( std__pe23__lane5_strm0_cntl       ),      
               .std__pe23__lane5_strm0_data          ( std__pe23__lane5_strm0_data       ),      
               .std__pe23__lane5_strm0_data_valid    ( std__pe23__lane5_strm0_data_valid ),      
               .std__pe23__lane5_strm0_data_mask     ( std__pe23__lane5_strm0_data_mask  ),      

               .pe23__std__lane5_strm1_ready         ( pe23__std__lane5_strm1_ready      ),      
               .std__pe23__lane5_strm1_cntl          ( std__pe23__lane5_strm1_cntl       ),      
               .std__pe23__lane5_strm1_data          ( std__pe23__lane5_strm1_data       ),      
               .std__pe23__lane5_strm1_data_valid    ( std__pe23__lane5_strm1_data_valid ),      
               .std__pe23__lane5_strm1_data_mask     ( std__pe23__lane5_strm1_data_mask  ),      

               // PE 23, Lane 6                 
               .pe23__std__lane6_strm0_ready         ( pe23__std__lane6_strm0_ready      ),      
               .std__pe23__lane6_strm0_cntl          ( std__pe23__lane6_strm0_cntl       ),      
               .std__pe23__lane6_strm0_data          ( std__pe23__lane6_strm0_data       ),      
               .std__pe23__lane6_strm0_data_valid    ( std__pe23__lane6_strm0_data_valid ),      
               .std__pe23__lane6_strm0_data_mask     ( std__pe23__lane6_strm0_data_mask  ),      

               .pe23__std__lane6_strm1_ready         ( pe23__std__lane6_strm1_ready      ),      
               .std__pe23__lane6_strm1_cntl          ( std__pe23__lane6_strm1_cntl       ),      
               .std__pe23__lane6_strm1_data          ( std__pe23__lane6_strm1_data       ),      
               .std__pe23__lane6_strm1_data_valid    ( std__pe23__lane6_strm1_data_valid ),      
               .std__pe23__lane6_strm1_data_mask     ( std__pe23__lane6_strm1_data_mask  ),      

               // PE 23, Lane 7                 
               .pe23__std__lane7_strm0_ready         ( pe23__std__lane7_strm0_ready      ),      
               .std__pe23__lane7_strm0_cntl          ( std__pe23__lane7_strm0_cntl       ),      
               .std__pe23__lane7_strm0_data          ( std__pe23__lane7_strm0_data       ),      
               .std__pe23__lane7_strm0_data_valid    ( std__pe23__lane7_strm0_data_valid ),      
               .std__pe23__lane7_strm0_data_mask     ( std__pe23__lane7_strm0_data_mask  ),      

               .pe23__std__lane7_strm1_ready         ( pe23__std__lane7_strm1_ready      ),      
               .std__pe23__lane7_strm1_cntl          ( std__pe23__lane7_strm1_cntl       ),      
               .std__pe23__lane7_strm1_data          ( std__pe23__lane7_strm1_data       ),      
               .std__pe23__lane7_strm1_data_valid    ( std__pe23__lane7_strm1_data_valid ),      
               .std__pe23__lane7_strm1_data_mask     ( std__pe23__lane7_strm1_data_mask  ),      

               // PE 23, Lane 8                 
               .pe23__std__lane8_strm0_ready         ( pe23__std__lane8_strm0_ready      ),      
               .std__pe23__lane8_strm0_cntl          ( std__pe23__lane8_strm0_cntl       ),      
               .std__pe23__lane8_strm0_data          ( std__pe23__lane8_strm0_data       ),      
               .std__pe23__lane8_strm0_data_valid    ( std__pe23__lane8_strm0_data_valid ),      
               .std__pe23__lane8_strm0_data_mask     ( std__pe23__lane8_strm0_data_mask  ),      

               .pe23__std__lane8_strm1_ready         ( pe23__std__lane8_strm1_ready      ),      
               .std__pe23__lane8_strm1_cntl          ( std__pe23__lane8_strm1_cntl       ),      
               .std__pe23__lane8_strm1_data          ( std__pe23__lane8_strm1_data       ),      
               .std__pe23__lane8_strm1_data_valid    ( std__pe23__lane8_strm1_data_valid ),      
               .std__pe23__lane8_strm1_data_mask     ( std__pe23__lane8_strm1_data_mask  ),      

               // PE 23, Lane 9                 
               .pe23__std__lane9_strm0_ready         ( pe23__std__lane9_strm0_ready      ),      
               .std__pe23__lane9_strm0_cntl          ( std__pe23__lane9_strm0_cntl       ),      
               .std__pe23__lane9_strm0_data          ( std__pe23__lane9_strm0_data       ),      
               .std__pe23__lane9_strm0_data_valid    ( std__pe23__lane9_strm0_data_valid ),      
               .std__pe23__lane9_strm0_data_mask     ( std__pe23__lane9_strm0_data_mask  ),      

               .pe23__std__lane9_strm1_ready         ( pe23__std__lane9_strm1_ready      ),      
               .std__pe23__lane9_strm1_cntl          ( std__pe23__lane9_strm1_cntl       ),      
               .std__pe23__lane9_strm1_data          ( std__pe23__lane9_strm1_data       ),      
               .std__pe23__lane9_strm1_data_valid    ( std__pe23__lane9_strm1_data_valid ),      
               .std__pe23__lane9_strm1_data_mask     ( std__pe23__lane9_strm1_data_mask  ),      

               // PE 23, Lane 10                 
               .pe23__std__lane10_strm0_ready         ( pe23__std__lane10_strm0_ready      ),      
               .std__pe23__lane10_strm0_cntl          ( std__pe23__lane10_strm0_cntl       ),      
               .std__pe23__lane10_strm0_data          ( std__pe23__lane10_strm0_data       ),      
               .std__pe23__lane10_strm0_data_valid    ( std__pe23__lane10_strm0_data_valid ),      
               .std__pe23__lane10_strm0_data_mask     ( std__pe23__lane10_strm0_data_mask  ),      

               .pe23__std__lane10_strm1_ready         ( pe23__std__lane10_strm1_ready      ),      
               .std__pe23__lane10_strm1_cntl          ( std__pe23__lane10_strm1_cntl       ),      
               .std__pe23__lane10_strm1_data          ( std__pe23__lane10_strm1_data       ),      
               .std__pe23__lane10_strm1_data_valid    ( std__pe23__lane10_strm1_data_valid ),      
               .std__pe23__lane10_strm1_data_mask     ( std__pe23__lane10_strm1_data_mask  ),      

               // PE 23, Lane 11                 
               .pe23__std__lane11_strm0_ready         ( pe23__std__lane11_strm0_ready      ),      
               .std__pe23__lane11_strm0_cntl          ( std__pe23__lane11_strm0_cntl       ),      
               .std__pe23__lane11_strm0_data          ( std__pe23__lane11_strm0_data       ),      
               .std__pe23__lane11_strm0_data_valid    ( std__pe23__lane11_strm0_data_valid ),      
               .std__pe23__lane11_strm0_data_mask     ( std__pe23__lane11_strm0_data_mask  ),      

               .pe23__std__lane11_strm1_ready         ( pe23__std__lane11_strm1_ready      ),      
               .std__pe23__lane11_strm1_cntl          ( std__pe23__lane11_strm1_cntl       ),      
               .std__pe23__lane11_strm1_data          ( std__pe23__lane11_strm1_data       ),      
               .std__pe23__lane11_strm1_data_valid    ( std__pe23__lane11_strm1_data_valid ),      
               .std__pe23__lane11_strm1_data_mask     ( std__pe23__lane11_strm1_data_mask  ),      

               // PE 23, Lane 12                 
               .pe23__std__lane12_strm0_ready         ( pe23__std__lane12_strm0_ready      ),      
               .std__pe23__lane12_strm0_cntl          ( std__pe23__lane12_strm0_cntl       ),      
               .std__pe23__lane12_strm0_data          ( std__pe23__lane12_strm0_data       ),      
               .std__pe23__lane12_strm0_data_valid    ( std__pe23__lane12_strm0_data_valid ),      
               .std__pe23__lane12_strm0_data_mask     ( std__pe23__lane12_strm0_data_mask  ),      

               .pe23__std__lane12_strm1_ready         ( pe23__std__lane12_strm1_ready      ),      
               .std__pe23__lane12_strm1_cntl          ( std__pe23__lane12_strm1_cntl       ),      
               .std__pe23__lane12_strm1_data          ( std__pe23__lane12_strm1_data       ),      
               .std__pe23__lane12_strm1_data_valid    ( std__pe23__lane12_strm1_data_valid ),      
               .std__pe23__lane12_strm1_data_mask     ( std__pe23__lane12_strm1_data_mask  ),      

               // PE 23, Lane 13                 
               .pe23__std__lane13_strm0_ready         ( pe23__std__lane13_strm0_ready      ),      
               .std__pe23__lane13_strm0_cntl          ( std__pe23__lane13_strm0_cntl       ),      
               .std__pe23__lane13_strm0_data          ( std__pe23__lane13_strm0_data       ),      
               .std__pe23__lane13_strm0_data_valid    ( std__pe23__lane13_strm0_data_valid ),      
               .std__pe23__lane13_strm0_data_mask     ( std__pe23__lane13_strm0_data_mask  ),      

               .pe23__std__lane13_strm1_ready         ( pe23__std__lane13_strm1_ready      ),      
               .std__pe23__lane13_strm1_cntl          ( std__pe23__lane13_strm1_cntl       ),      
               .std__pe23__lane13_strm1_data          ( std__pe23__lane13_strm1_data       ),      
               .std__pe23__lane13_strm1_data_valid    ( std__pe23__lane13_strm1_data_valid ),      
               .std__pe23__lane13_strm1_data_mask     ( std__pe23__lane13_strm1_data_mask  ),      

               // PE 23, Lane 14                 
               .pe23__std__lane14_strm0_ready         ( pe23__std__lane14_strm0_ready      ),      
               .std__pe23__lane14_strm0_cntl          ( std__pe23__lane14_strm0_cntl       ),      
               .std__pe23__lane14_strm0_data          ( std__pe23__lane14_strm0_data       ),      
               .std__pe23__lane14_strm0_data_valid    ( std__pe23__lane14_strm0_data_valid ),      
               .std__pe23__lane14_strm0_data_mask     ( std__pe23__lane14_strm0_data_mask  ),      

               .pe23__std__lane14_strm1_ready         ( pe23__std__lane14_strm1_ready      ),      
               .std__pe23__lane14_strm1_cntl          ( std__pe23__lane14_strm1_cntl       ),      
               .std__pe23__lane14_strm1_data          ( std__pe23__lane14_strm1_data       ),      
               .std__pe23__lane14_strm1_data_valid    ( std__pe23__lane14_strm1_data_valid ),      
               .std__pe23__lane14_strm1_data_mask     ( std__pe23__lane14_strm1_data_mask  ),      

               // PE 23, Lane 15                 
               .pe23__std__lane15_strm0_ready         ( pe23__std__lane15_strm0_ready      ),      
               .std__pe23__lane15_strm0_cntl          ( std__pe23__lane15_strm0_cntl       ),      
               .std__pe23__lane15_strm0_data          ( std__pe23__lane15_strm0_data       ),      
               .std__pe23__lane15_strm0_data_valid    ( std__pe23__lane15_strm0_data_valid ),      
               .std__pe23__lane15_strm0_data_mask     ( std__pe23__lane15_strm0_data_mask  ),      

               .pe23__std__lane15_strm1_ready         ( pe23__std__lane15_strm1_ready      ),      
               .std__pe23__lane15_strm1_cntl          ( std__pe23__lane15_strm1_cntl       ),      
               .std__pe23__lane15_strm1_data          ( std__pe23__lane15_strm1_data       ),      
               .std__pe23__lane15_strm1_data_valid    ( std__pe23__lane15_strm1_data_valid ),      
               .std__pe23__lane15_strm1_data_mask     ( std__pe23__lane15_strm1_data_mask  ),      

               // PE 23, Lane 16                 
               .pe23__std__lane16_strm0_ready         ( pe23__std__lane16_strm0_ready      ),      
               .std__pe23__lane16_strm0_cntl          ( std__pe23__lane16_strm0_cntl       ),      
               .std__pe23__lane16_strm0_data          ( std__pe23__lane16_strm0_data       ),      
               .std__pe23__lane16_strm0_data_valid    ( std__pe23__lane16_strm0_data_valid ),      
               .std__pe23__lane16_strm0_data_mask     ( std__pe23__lane16_strm0_data_mask  ),      

               .pe23__std__lane16_strm1_ready         ( pe23__std__lane16_strm1_ready      ),      
               .std__pe23__lane16_strm1_cntl          ( std__pe23__lane16_strm1_cntl       ),      
               .std__pe23__lane16_strm1_data          ( std__pe23__lane16_strm1_data       ),      
               .std__pe23__lane16_strm1_data_valid    ( std__pe23__lane16_strm1_data_valid ),      
               .std__pe23__lane16_strm1_data_mask     ( std__pe23__lane16_strm1_data_mask  ),      

               // PE 23, Lane 17                 
               .pe23__std__lane17_strm0_ready         ( pe23__std__lane17_strm0_ready      ),      
               .std__pe23__lane17_strm0_cntl          ( std__pe23__lane17_strm0_cntl       ),      
               .std__pe23__lane17_strm0_data          ( std__pe23__lane17_strm0_data       ),      
               .std__pe23__lane17_strm0_data_valid    ( std__pe23__lane17_strm0_data_valid ),      
               .std__pe23__lane17_strm0_data_mask     ( std__pe23__lane17_strm0_data_mask  ),      

               .pe23__std__lane17_strm1_ready         ( pe23__std__lane17_strm1_ready      ),      
               .std__pe23__lane17_strm1_cntl          ( std__pe23__lane17_strm1_cntl       ),      
               .std__pe23__lane17_strm1_data          ( std__pe23__lane17_strm1_data       ),      
               .std__pe23__lane17_strm1_data_valid    ( std__pe23__lane17_strm1_data_valid ),      
               .std__pe23__lane17_strm1_data_mask     ( std__pe23__lane17_strm1_data_mask  ),      

               // PE 23, Lane 18                 
               .pe23__std__lane18_strm0_ready         ( pe23__std__lane18_strm0_ready      ),      
               .std__pe23__lane18_strm0_cntl          ( std__pe23__lane18_strm0_cntl       ),      
               .std__pe23__lane18_strm0_data          ( std__pe23__lane18_strm0_data       ),      
               .std__pe23__lane18_strm0_data_valid    ( std__pe23__lane18_strm0_data_valid ),      
               .std__pe23__lane18_strm0_data_mask     ( std__pe23__lane18_strm0_data_mask  ),      

               .pe23__std__lane18_strm1_ready         ( pe23__std__lane18_strm1_ready      ),      
               .std__pe23__lane18_strm1_cntl          ( std__pe23__lane18_strm1_cntl       ),      
               .std__pe23__lane18_strm1_data          ( std__pe23__lane18_strm1_data       ),      
               .std__pe23__lane18_strm1_data_valid    ( std__pe23__lane18_strm1_data_valid ),      
               .std__pe23__lane18_strm1_data_mask     ( std__pe23__lane18_strm1_data_mask  ),      

               // PE 23, Lane 19                 
               .pe23__std__lane19_strm0_ready         ( pe23__std__lane19_strm0_ready      ),      
               .std__pe23__lane19_strm0_cntl          ( std__pe23__lane19_strm0_cntl       ),      
               .std__pe23__lane19_strm0_data          ( std__pe23__lane19_strm0_data       ),      
               .std__pe23__lane19_strm0_data_valid    ( std__pe23__lane19_strm0_data_valid ),      
               .std__pe23__lane19_strm0_data_mask     ( std__pe23__lane19_strm0_data_mask  ),      

               .pe23__std__lane19_strm1_ready         ( pe23__std__lane19_strm1_ready      ),      
               .std__pe23__lane19_strm1_cntl          ( std__pe23__lane19_strm1_cntl       ),      
               .std__pe23__lane19_strm1_data          ( std__pe23__lane19_strm1_data       ),      
               .std__pe23__lane19_strm1_data_valid    ( std__pe23__lane19_strm1_data_valid ),      
               .std__pe23__lane19_strm1_data_mask     ( std__pe23__lane19_strm1_data_mask  ),      

               // PE 23, Lane 20                 
               .pe23__std__lane20_strm0_ready         ( pe23__std__lane20_strm0_ready      ),      
               .std__pe23__lane20_strm0_cntl          ( std__pe23__lane20_strm0_cntl       ),      
               .std__pe23__lane20_strm0_data          ( std__pe23__lane20_strm0_data       ),      
               .std__pe23__lane20_strm0_data_valid    ( std__pe23__lane20_strm0_data_valid ),      
               .std__pe23__lane20_strm0_data_mask     ( std__pe23__lane20_strm0_data_mask  ),      

               .pe23__std__lane20_strm1_ready         ( pe23__std__lane20_strm1_ready      ),      
               .std__pe23__lane20_strm1_cntl          ( std__pe23__lane20_strm1_cntl       ),      
               .std__pe23__lane20_strm1_data          ( std__pe23__lane20_strm1_data       ),      
               .std__pe23__lane20_strm1_data_valid    ( std__pe23__lane20_strm1_data_valid ),      
               .std__pe23__lane20_strm1_data_mask     ( std__pe23__lane20_strm1_data_mask  ),      

               // PE 23, Lane 21                 
               .pe23__std__lane21_strm0_ready         ( pe23__std__lane21_strm0_ready      ),      
               .std__pe23__lane21_strm0_cntl          ( std__pe23__lane21_strm0_cntl       ),      
               .std__pe23__lane21_strm0_data          ( std__pe23__lane21_strm0_data       ),      
               .std__pe23__lane21_strm0_data_valid    ( std__pe23__lane21_strm0_data_valid ),      
               .std__pe23__lane21_strm0_data_mask     ( std__pe23__lane21_strm0_data_mask  ),      

               .pe23__std__lane21_strm1_ready         ( pe23__std__lane21_strm1_ready      ),      
               .std__pe23__lane21_strm1_cntl          ( std__pe23__lane21_strm1_cntl       ),      
               .std__pe23__lane21_strm1_data          ( std__pe23__lane21_strm1_data       ),      
               .std__pe23__lane21_strm1_data_valid    ( std__pe23__lane21_strm1_data_valid ),      
               .std__pe23__lane21_strm1_data_mask     ( std__pe23__lane21_strm1_data_mask  ),      

               // PE 23, Lane 22                 
               .pe23__std__lane22_strm0_ready         ( pe23__std__lane22_strm0_ready      ),      
               .std__pe23__lane22_strm0_cntl          ( std__pe23__lane22_strm0_cntl       ),      
               .std__pe23__lane22_strm0_data          ( std__pe23__lane22_strm0_data       ),      
               .std__pe23__lane22_strm0_data_valid    ( std__pe23__lane22_strm0_data_valid ),      
               .std__pe23__lane22_strm0_data_mask     ( std__pe23__lane22_strm0_data_mask  ),      

               .pe23__std__lane22_strm1_ready         ( pe23__std__lane22_strm1_ready      ),      
               .std__pe23__lane22_strm1_cntl          ( std__pe23__lane22_strm1_cntl       ),      
               .std__pe23__lane22_strm1_data          ( std__pe23__lane22_strm1_data       ),      
               .std__pe23__lane22_strm1_data_valid    ( std__pe23__lane22_strm1_data_valid ),      
               .std__pe23__lane22_strm1_data_mask     ( std__pe23__lane22_strm1_data_mask  ),      

               // PE 23, Lane 23                 
               .pe23__std__lane23_strm0_ready         ( pe23__std__lane23_strm0_ready      ),      
               .std__pe23__lane23_strm0_cntl          ( std__pe23__lane23_strm0_cntl       ),      
               .std__pe23__lane23_strm0_data          ( std__pe23__lane23_strm0_data       ),      
               .std__pe23__lane23_strm0_data_valid    ( std__pe23__lane23_strm0_data_valid ),      
               .std__pe23__lane23_strm0_data_mask     ( std__pe23__lane23_strm0_data_mask  ),      

               .pe23__std__lane23_strm1_ready         ( pe23__std__lane23_strm1_ready      ),      
               .std__pe23__lane23_strm1_cntl          ( std__pe23__lane23_strm1_cntl       ),      
               .std__pe23__lane23_strm1_data          ( std__pe23__lane23_strm1_data       ),      
               .std__pe23__lane23_strm1_data_valid    ( std__pe23__lane23_strm1_data_valid ),      
               .std__pe23__lane23_strm1_data_mask     ( std__pe23__lane23_strm1_data_mask  ),      

               // PE 23, Lane 24                 
               .pe23__std__lane24_strm0_ready         ( pe23__std__lane24_strm0_ready      ),      
               .std__pe23__lane24_strm0_cntl          ( std__pe23__lane24_strm0_cntl       ),      
               .std__pe23__lane24_strm0_data          ( std__pe23__lane24_strm0_data       ),      
               .std__pe23__lane24_strm0_data_valid    ( std__pe23__lane24_strm0_data_valid ),      
               .std__pe23__lane24_strm0_data_mask     ( std__pe23__lane24_strm0_data_mask  ),      

               .pe23__std__lane24_strm1_ready         ( pe23__std__lane24_strm1_ready      ),      
               .std__pe23__lane24_strm1_cntl          ( std__pe23__lane24_strm1_cntl       ),      
               .std__pe23__lane24_strm1_data          ( std__pe23__lane24_strm1_data       ),      
               .std__pe23__lane24_strm1_data_valid    ( std__pe23__lane24_strm1_data_valid ),      
               .std__pe23__lane24_strm1_data_mask     ( std__pe23__lane24_strm1_data_mask  ),      

               // PE 23, Lane 25                 
               .pe23__std__lane25_strm0_ready         ( pe23__std__lane25_strm0_ready      ),      
               .std__pe23__lane25_strm0_cntl          ( std__pe23__lane25_strm0_cntl       ),      
               .std__pe23__lane25_strm0_data          ( std__pe23__lane25_strm0_data       ),      
               .std__pe23__lane25_strm0_data_valid    ( std__pe23__lane25_strm0_data_valid ),      
               .std__pe23__lane25_strm0_data_mask     ( std__pe23__lane25_strm0_data_mask  ),      

               .pe23__std__lane25_strm1_ready         ( pe23__std__lane25_strm1_ready      ),      
               .std__pe23__lane25_strm1_cntl          ( std__pe23__lane25_strm1_cntl       ),      
               .std__pe23__lane25_strm1_data          ( std__pe23__lane25_strm1_data       ),      
               .std__pe23__lane25_strm1_data_valid    ( std__pe23__lane25_strm1_data_valid ),      
               .std__pe23__lane25_strm1_data_mask     ( std__pe23__lane25_strm1_data_mask  ),      

               // PE 23, Lane 26                 
               .pe23__std__lane26_strm0_ready         ( pe23__std__lane26_strm0_ready      ),      
               .std__pe23__lane26_strm0_cntl          ( std__pe23__lane26_strm0_cntl       ),      
               .std__pe23__lane26_strm0_data          ( std__pe23__lane26_strm0_data       ),      
               .std__pe23__lane26_strm0_data_valid    ( std__pe23__lane26_strm0_data_valid ),      
               .std__pe23__lane26_strm0_data_mask     ( std__pe23__lane26_strm0_data_mask  ),      

               .pe23__std__lane26_strm1_ready         ( pe23__std__lane26_strm1_ready      ),      
               .std__pe23__lane26_strm1_cntl          ( std__pe23__lane26_strm1_cntl       ),      
               .std__pe23__lane26_strm1_data          ( std__pe23__lane26_strm1_data       ),      
               .std__pe23__lane26_strm1_data_valid    ( std__pe23__lane26_strm1_data_valid ),      
               .std__pe23__lane26_strm1_data_mask     ( std__pe23__lane26_strm1_data_mask  ),      

               // PE 23, Lane 27                 
               .pe23__std__lane27_strm0_ready         ( pe23__std__lane27_strm0_ready      ),      
               .std__pe23__lane27_strm0_cntl          ( std__pe23__lane27_strm0_cntl       ),      
               .std__pe23__lane27_strm0_data          ( std__pe23__lane27_strm0_data       ),      
               .std__pe23__lane27_strm0_data_valid    ( std__pe23__lane27_strm0_data_valid ),      
               .std__pe23__lane27_strm0_data_mask     ( std__pe23__lane27_strm0_data_mask  ),      

               .pe23__std__lane27_strm1_ready         ( pe23__std__lane27_strm1_ready      ),      
               .std__pe23__lane27_strm1_cntl          ( std__pe23__lane27_strm1_cntl       ),      
               .std__pe23__lane27_strm1_data          ( std__pe23__lane27_strm1_data       ),      
               .std__pe23__lane27_strm1_data_valid    ( std__pe23__lane27_strm1_data_valid ),      
               .std__pe23__lane27_strm1_data_mask     ( std__pe23__lane27_strm1_data_mask  ),      

               // PE 23, Lane 28                 
               .pe23__std__lane28_strm0_ready         ( pe23__std__lane28_strm0_ready      ),      
               .std__pe23__lane28_strm0_cntl          ( std__pe23__lane28_strm0_cntl       ),      
               .std__pe23__lane28_strm0_data          ( std__pe23__lane28_strm0_data       ),      
               .std__pe23__lane28_strm0_data_valid    ( std__pe23__lane28_strm0_data_valid ),      
               .std__pe23__lane28_strm0_data_mask     ( std__pe23__lane28_strm0_data_mask  ),      

               .pe23__std__lane28_strm1_ready         ( pe23__std__lane28_strm1_ready      ),      
               .std__pe23__lane28_strm1_cntl          ( std__pe23__lane28_strm1_cntl       ),      
               .std__pe23__lane28_strm1_data          ( std__pe23__lane28_strm1_data       ),      
               .std__pe23__lane28_strm1_data_valid    ( std__pe23__lane28_strm1_data_valid ),      
               .std__pe23__lane28_strm1_data_mask     ( std__pe23__lane28_strm1_data_mask  ),      

               // PE 23, Lane 29                 
               .pe23__std__lane29_strm0_ready         ( pe23__std__lane29_strm0_ready      ),      
               .std__pe23__lane29_strm0_cntl          ( std__pe23__lane29_strm0_cntl       ),      
               .std__pe23__lane29_strm0_data          ( std__pe23__lane29_strm0_data       ),      
               .std__pe23__lane29_strm0_data_valid    ( std__pe23__lane29_strm0_data_valid ),      
               .std__pe23__lane29_strm0_data_mask     ( std__pe23__lane29_strm0_data_mask  ),      

               .pe23__std__lane29_strm1_ready         ( pe23__std__lane29_strm1_ready      ),      
               .std__pe23__lane29_strm1_cntl          ( std__pe23__lane29_strm1_cntl       ),      
               .std__pe23__lane29_strm1_data          ( std__pe23__lane29_strm1_data       ),      
               .std__pe23__lane29_strm1_data_valid    ( std__pe23__lane29_strm1_data_valid ),      
               .std__pe23__lane29_strm1_data_mask     ( std__pe23__lane29_strm1_data_mask  ),      

               // PE 23, Lane 30                 
               .pe23__std__lane30_strm0_ready         ( pe23__std__lane30_strm0_ready      ),      
               .std__pe23__lane30_strm0_cntl          ( std__pe23__lane30_strm0_cntl       ),      
               .std__pe23__lane30_strm0_data          ( std__pe23__lane30_strm0_data       ),      
               .std__pe23__lane30_strm0_data_valid    ( std__pe23__lane30_strm0_data_valid ),      
               .std__pe23__lane30_strm0_data_mask     ( std__pe23__lane30_strm0_data_mask  ),      

               .pe23__std__lane30_strm1_ready         ( pe23__std__lane30_strm1_ready      ),      
               .std__pe23__lane30_strm1_cntl          ( std__pe23__lane30_strm1_cntl       ),      
               .std__pe23__lane30_strm1_data          ( std__pe23__lane30_strm1_data       ),      
               .std__pe23__lane30_strm1_data_valid    ( std__pe23__lane30_strm1_data_valid ),      
               .std__pe23__lane30_strm1_data_mask     ( std__pe23__lane30_strm1_data_mask  ),      

               // PE 23, Lane 31                 
               .pe23__std__lane31_strm0_ready         ( pe23__std__lane31_strm0_ready      ),      
               .std__pe23__lane31_strm0_cntl          ( std__pe23__lane31_strm0_cntl       ),      
               .std__pe23__lane31_strm0_data          ( std__pe23__lane31_strm0_data       ),      
               .std__pe23__lane31_strm0_data_valid    ( std__pe23__lane31_strm0_data_valid ),      
               .std__pe23__lane31_strm0_data_mask     ( std__pe23__lane31_strm0_data_mask  ),      

               .pe23__std__lane31_strm1_ready         ( pe23__std__lane31_strm1_ready      ),      
               .std__pe23__lane31_strm1_cntl          ( std__pe23__lane31_strm1_cntl       ),      
               .std__pe23__lane31_strm1_data          ( std__pe23__lane31_strm1_data       ),      
               .std__pe23__lane31_strm1_data_valid    ( std__pe23__lane31_strm1_data_valid ),      
               .std__pe23__lane31_strm1_data_mask     ( std__pe23__lane31_strm1_data_mask  ),      

               // PE 24, Lane 0                 
               .pe24__std__lane0_strm0_ready         ( pe24__std__lane0_strm0_ready      ),      
               .std__pe24__lane0_strm0_cntl          ( std__pe24__lane0_strm0_cntl       ),      
               .std__pe24__lane0_strm0_data          ( std__pe24__lane0_strm0_data       ),      
               .std__pe24__lane0_strm0_data_valid    ( std__pe24__lane0_strm0_data_valid ),      
               .std__pe24__lane0_strm0_data_mask     ( std__pe24__lane0_strm0_data_mask  ),      

               .pe24__std__lane0_strm1_ready         ( pe24__std__lane0_strm1_ready      ),      
               .std__pe24__lane0_strm1_cntl          ( std__pe24__lane0_strm1_cntl       ),      
               .std__pe24__lane0_strm1_data          ( std__pe24__lane0_strm1_data       ),      
               .std__pe24__lane0_strm1_data_valid    ( std__pe24__lane0_strm1_data_valid ),      
               .std__pe24__lane0_strm1_data_mask     ( std__pe24__lane0_strm1_data_mask  ),      

               // PE 24, Lane 1                 
               .pe24__std__lane1_strm0_ready         ( pe24__std__lane1_strm0_ready      ),      
               .std__pe24__lane1_strm0_cntl          ( std__pe24__lane1_strm0_cntl       ),      
               .std__pe24__lane1_strm0_data          ( std__pe24__lane1_strm0_data       ),      
               .std__pe24__lane1_strm0_data_valid    ( std__pe24__lane1_strm0_data_valid ),      
               .std__pe24__lane1_strm0_data_mask     ( std__pe24__lane1_strm0_data_mask  ),      

               .pe24__std__lane1_strm1_ready         ( pe24__std__lane1_strm1_ready      ),      
               .std__pe24__lane1_strm1_cntl          ( std__pe24__lane1_strm1_cntl       ),      
               .std__pe24__lane1_strm1_data          ( std__pe24__lane1_strm1_data       ),      
               .std__pe24__lane1_strm1_data_valid    ( std__pe24__lane1_strm1_data_valid ),      
               .std__pe24__lane1_strm1_data_mask     ( std__pe24__lane1_strm1_data_mask  ),      

               // PE 24, Lane 2                 
               .pe24__std__lane2_strm0_ready         ( pe24__std__lane2_strm0_ready      ),      
               .std__pe24__lane2_strm0_cntl          ( std__pe24__lane2_strm0_cntl       ),      
               .std__pe24__lane2_strm0_data          ( std__pe24__lane2_strm0_data       ),      
               .std__pe24__lane2_strm0_data_valid    ( std__pe24__lane2_strm0_data_valid ),      
               .std__pe24__lane2_strm0_data_mask     ( std__pe24__lane2_strm0_data_mask  ),      

               .pe24__std__lane2_strm1_ready         ( pe24__std__lane2_strm1_ready      ),      
               .std__pe24__lane2_strm1_cntl          ( std__pe24__lane2_strm1_cntl       ),      
               .std__pe24__lane2_strm1_data          ( std__pe24__lane2_strm1_data       ),      
               .std__pe24__lane2_strm1_data_valid    ( std__pe24__lane2_strm1_data_valid ),      
               .std__pe24__lane2_strm1_data_mask     ( std__pe24__lane2_strm1_data_mask  ),      

               // PE 24, Lane 3                 
               .pe24__std__lane3_strm0_ready         ( pe24__std__lane3_strm0_ready      ),      
               .std__pe24__lane3_strm0_cntl          ( std__pe24__lane3_strm0_cntl       ),      
               .std__pe24__lane3_strm0_data          ( std__pe24__lane3_strm0_data       ),      
               .std__pe24__lane3_strm0_data_valid    ( std__pe24__lane3_strm0_data_valid ),      
               .std__pe24__lane3_strm0_data_mask     ( std__pe24__lane3_strm0_data_mask  ),      

               .pe24__std__lane3_strm1_ready         ( pe24__std__lane3_strm1_ready      ),      
               .std__pe24__lane3_strm1_cntl          ( std__pe24__lane3_strm1_cntl       ),      
               .std__pe24__lane3_strm1_data          ( std__pe24__lane3_strm1_data       ),      
               .std__pe24__lane3_strm1_data_valid    ( std__pe24__lane3_strm1_data_valid ),      
               .std__pe24__lane3_strm1_data_mask     ( std__pe24__lane3_strm1_data_mask  ),      

               // PE 24, Lane 4                 
               .pe24__std__lane4_strm0_ready         ( pe24__std__lane4_strm0_ready      ),      
               .std__pe24__lane4_strm0_cntl          ( std__pe24__lane4_strm0_cntl       ),      
               .std__pe24__lane4_strm0_data          ( std__pe24__lane4_strm0_data       ),      
               .std__pe24__lane4_strm0_data_valid    ( std__pe24__lane4_strm0_data_valid ),      
               .std__pe24__lane4_strm0_data_mask     ( std__pe24__lane4_strm0_data_mask  ),      

               .pe24__std__lane4_strm1_ready         ( pe24__std__lane4_strm1_ready      ),      
               .std__pe24__lane4_strm1_cntl          ( std__pe24__lane4_strm1_cntl       ),      
               .std__pe24__lane4_strm1_data          ( std__pe24__lane4_strm1_data       ),      
               .std__pe24__lane4_strm1_data_valid    ( std__pe24__lane4_strm1_data_valid ),      
               .std__pe24__lane4_strm1_data_mask     ( std__pe24__lane4_strm1_data_mask  ),      

               // PE 24, Lane 5                 
               .pe24__std__lane5_strm0_ready         ( pe24__std__lane5_strm0_ready      ),      
               .std__pe24__lane5_strm0_cntl          ( std__pe24__lane5_strm0_cntl       ),      
               .std__pe24__lane5_strm0_data          ( std__pe24__lane5_strm0_data       ),      
               .std__pe24__lane5_strm0_data_valid    ( std__pe24__lane5_strm0_data_valid ),      
               .std__pe24__lane5_strm0_data_mask     ( std__pe24__lane5_strm0_data_mask  ),      

               .pe24__std__lane5_strm1_ready         ( pe24__std__lane5_strm1_ready      ),      
               .std__pe24__lane5_strm1_cntl          ( std__pe24__lane5_strm1_cntl       ),      
               .std__pe24__lane5_strm1_data          ( std__pe24__lane5_strm1_data       ),      
               .std__pe24__lane5_strm1_data_valid    ( std__pe24__lane5_strm1_data_valid ),      
               .std__pe24__lane5_strm1_data_mask     ( std__pe24__lane5_strm1_data_mask  ),      

               // PE 24, Lane 6                 
               .pe24__std__lane6_strm0_ready         ( pe24__std__lane6_strm0_ready      ),      
               .std__pe24__lane6_strm0_cntl          ( std__pe24__lane6_strm0_cntl       ),      
               .std__pe24__lane6_strm0_data          ( std__pe24__lane6_strm0_data       ),      
               .std__pe24__lane6_strm0_data_valid    ( std__pe24__lane6_strm0_data_valid ),      
               .std__pe24__lane6_strm0_data_mask     ( std__pe24__lane6_strm0_data_mask  ),      

               .pe24__std__lane6_strm1_ready         ( pe24__std__lane6_strm1_ready      ),      
               .std__pe24__lane6_strm1_cntl          ( std__pe24__lane6_strm1_cntl       ),      
               .std__pe24__lane6_strm1_data          ( std__pe24__lane6_strm1_data       ),      
               .std__pe24__lane6_strm1_data_valid    ( std__pe24__lane6_strm1_data_valid ),      
               .std__pe24__lane6_strm1_data_mask     ( std__pe24__lane6_strm1_data_mask  ),      

               // PE 24, Lane 7                 
               .pe24__std__lane7_strm0_ready         ( pe24__std__lane7_strm0_ready      ),      
               .std__pe24__lane7_strm0_cntl          ( std__pe24__lane7_strm0_cntl       ),      
               .std__pe24__lane7_strm0_data          ( std__pe24__lane7_strm0_data       ),      
               .std__pe24__lane7_strm0_data_valid    ( std__pe24__lane7_strm0_data_valid ),      
               .std__pe24__lane7_strm0_data_mask     ( std__pe24__lane7_strm0_data_mask  ),      

               .pe24__std__lane7_strm1_ready         ( pe24__std__lane7_strm1_ready      ),      
               .std__pe24__lane7_strm1_cntl          ( std__pe24__lane7_strm1_cntl       ),      
               .std__pe24__lane7_strm1_data          ( std__pe24__lane7_strm1_data       ),      
               .std__pe24__lane7_strm1_data_valid    ( std__pe24__lane7_strm1_data_valid ),      
               .std__pe24__lane7_strm1_data_mask     ( std__pe24__lane7_strm1_data_mask  ),      

               // PE 24, Lane 8                 
               .pe24__std__lane8_strm0_ready         ( pe24__std__lane8_strm0_ready      ),      
               .std__pe24__lane8_strm0_cntl          ( std__pe24__lane8_strm0_cntl       ),      
               .std__pe24__lane8_strm0_data          ( std__pe24__lane8_strm0_data       ),      
               .std__pe24__lane8_strm0_data_valid    ( std__pe24__lane8_strm0_data_valid ),      
               .std__pe24__lane8_strm0_data_mask     ( std__pe24__lane8_strm0_data_mask  ),      

               .pe24__std__lane8_strm1_ready         ( pe24__std__lane8_strm1_ready      ),      
               .std__pe24__lane8_strm1_cntl          ( std__pe24__lane8_strm1_cntl       ),      
               .std__pe24__lane8_strm1_data          ( std__pe24__lane8_strm1_data       ),      
               .std__pe24__lane8_strm1_data_valid    ( std__pe24__lane8_strm1_data_valid ),      
               .std__pe24__lane8_strm1_data_mask     ( std__pe24__lane8_strm1_data_mask  ),      

               // PE 24, Lane 9                 
               .pe24__std__lane9_strm0_ready         ( pe24__std__lane9_strm0_ready      ),      
               .std__pe24__lane9_strm0_cntl          ( std__pe24__lane9_strm0_cntl       ),      
               .std__pe24__lane9_strm0_data          ( std__pe24__lane9_strm0_data       ),      
               .std__pe24__lane9_strm0_data_valid    ( std__pe24__lane9_strm0_data_valid ),      
               .std__pe24__lane9_strm0_data_mask     ( std__pe24__lane9_strm0_data_mask  ),      

               .pe24__std__lane9_strm1_ready         ( pe24__std__lane9_strm1_ready      ),      
               .std__pe24__lane9_strm1_cntl          ( std__pe24__lane9_strm1_cntl       ),      
               .std__pe24__lane9_strm1_data          ( std__pe24__lane9_strm1_data       ),      
               .std__pe24__lane9_strm1_data_valid    ( std__pe24__lane9_strm1_data_valid ),      
               .std__pe24__lane9_strm1_data_mask     ( std__pe24__lane9_strm1_data_mask  ),      

               // PE 24, Lane 10                 
               .pe24__std__lane10_strm0_ready         ( pe24__std__lane10_strm0_ready      ),      
               .std__pe24__lane10_strm0_cntl          ( std__pe24__lane10_strm0_cntl       ),      
               .std__pe24__lane10_strm0_data          ( std__pe24__lane10_strm0_data       ),      
               .std__pe24__lane10_strm0_data_valid    ( std__pe24__lane10_strm0_data_valid ),      
               .std__pe24__lane10_strm0_data_mask     ( std__pe24__lane10_strm0_data_mask  ),      

               .pe24__std__lane10_strm1_ready         ( pe24__std__lane10_strm1_ready      ),      
               .std__pe24__lane10_strm1_cntl          ( std__pe24__lane10_strm1_cntl       ),      
               .std__pe24__lane10_strm1_data          ( std__pe24__lane10_strm1_data       ),      
               .std__pe24__lane10_strm1_data_valid    ( std__pe24__lane10_strm1_data_valid ),      
               .std__pe24__lane10_strm1_data_mask     ( std__pe24__lane10_strm1_data_mask  ),      

               // PE 24, Lane 11                 
               .pe24__std__lane11_strm0_ready         ( pe24__std__lane11_strm0_ready      ),      
               .std__pe24__lane11_strm0_cntl          ( std__pe24__lane11_strm0_cntl       ),      
               .std__pe24__lane11_strm0_data          ( std__pe24__lane11_strm0_data       ),      
               .std__pe24__lane11_strm0_data_valid    ( std__pe24__lane11_strm0_data_valid ),      
               .std__pe24__lane11_strm0_data_mask     ( std__pe24__lane11_strm0_data_mask  ),      

               .pe24__std__lane11_strm1_ready         ( pe24__std__lane11_strm1_ready      ),      
               .std__pe24__lane11_strm1_cntl          ( std__pe24__lane11_strm1_cntl       ),      
               .std__pe24__lane11_strm1_data          ( std__pe24__lane11_strm1_data       ),      
               .std__pe24__lane11_strm1_data_valid    ( std__pe24__lane11_strm1_data_valid ),      
               .std__pe24__lane11_strm1_data_mask     ( std__pe24__lane11_strm1_data_mask  ),      

               // PE 24, Lane 12                 
               .pe24__std__lane12_strm0_ready         ( pe24__std__lane12_strm0_ready      ),      
               .std__pe24__lane12_strm0_cntl          ( std__pe24__lane12_strm0_cntl       ),      
               .std__pe24__lane12_strm0_data          ( std__pe24__lane12_strm0_data       ),      
               .std__pe24__lane12_strm0_data_valid    ( std__pe24__lane12_strm0_data_valid ),      
               .std__pe24__lane12_strm0_data_mask     ( std__pe24__lane12_strm0_data_mask  ),      

               .pe24__std__lane12_strm1_ready         ( pe24__std__lane12_strm1_ready      ),      
               .std__pe24__lane12_strm1_cntl          ( std__pe24__lane12_strm1_cntl       ),      
               .std__pe24__lane12_strm1_data          ( std__pe24__lane12_strm1_data       ),      
               .std__pe24__lane12_strm1_data_valid    ( std__pe24__lane12_strm1_data_valid ),      
               .std__pe24__lane12_strm1_data_mask     ( std__pe24__lane12_strm1_data_mask  ),      

               // PE 24, Lane 13                 
               .pe24__std__lane13_strm0_ready         ( pe24__std__lane13_strm0_ready      ),      
               .std__pe24__lane13_strm0_cntl          ( std__pe24__lane13_strm0_cntl       ),      
               .std__pe24__lane13_strm0_data          ( std__pe24__lane13_strm0_data       ),      
               .std__pe24__lane13_strm0_data_valid    ( std__pe24__lane13_strm0_data_valid ),      
               .std__pe24__lane13_strm0_data_mask     ( std__pe24__lane13_strm0_data_mask  ),      

               .pe24__std__lane13_strm1_ready         ( pe24__std__lane13_strm1_ready      ),      
               .std__pe24__lane13_strm1_cntl          ( std__pe24__lane13_strm1_cntl       ),      
               .std__pe24__lane13_strm1_data          ( std__pe24__lane13_strm1_data       ),      
               .std__pe24__lane13_strm1_data_valid    ( std__pe24__lane13_strm1_data_valid ),      
               .std__pe24__lane13_strm1_data_mask     ( std__pe24__lane13_strm1_data_mask  ),      

               // PE 24, Lane 14                 
               .pe24__std__lane14_strm0_ready         ( pe24__std__lane14_strm0_ready      ),      
               .std__pe24__lane14_strm0_cntl          ( std__pe24__lane14_strm0_cntl       ),      
               .std__pe24__lane14_strm0_data          ( std__pe24__lane14_strm0_data       ),      
               .std__pe24__lane14_strm0_data_valid    ( std__pe24__lane14_strm0_data_valid ),      
               .std__pe24__lane14_strm0_data_mask     ( std__pe24__lane14_strm0_data_mask  ),      

               .pe24__std__lane14_strm1_ready         ( pe24__std__lane14_strm1_ready      ),      
               .std__pe24__lane14_strm1_cntl          ( std__pe24__lane14_strm1_cntl       ),      
               .std__pe24__lane14_strm1_data          ( std__pe24__lane14_strm1_data       ),      
               .std__pe24__lane14_strm1_data_valid    ( std__pe24__lane14_strm1_data_valid ),      
               .std__pe24__lane14_strm1_data_mask     ( std__pe24__lane14_strm1_data_mask  ),      

               // PE 24, Lane 15                 
               .pe24__std__lane15_strm0_ready         ( pe24__std__lane15_strm0_ready      ),      
               .std__pe24__lane15_strm0_cntl          ( std__pe24__lane15_strm0_cntl       ),      
               .std__pe24__lane15_strm0_data          ( std__pe24__lane15_strm0_data       ),      
               .std__pe24__lane15_strm0_data_valid    ( std__pe24__lane15_strm0_data_valid ),      
               .std__pe24__lane15_strm0_data_mask     ( std__pe24__lane15_strm0_data_mask  ),      

               .pe24__std__lane15_strm1_ready         ( pe24__std__lane15_strm1_ready      ),      
               .std__pe24__lane15_strm1_cntl          ( std__pe24__lane15_strm1_cntl       ),      
               .std__pe24__lane15_strm1_data          ( std__pe24__lane15_strm1_data       ),      
               .std__pe24__lane15_strm1_data_valid    ( std__pe24__lane15_strm1_data_valid ),      
               .std__pe24__lane15_strm1_data_mask     ( std__pe24__lane15_strm1_data_mask  ),      

               // PE 24, Lane 16                 
               .pe24__std__lane16_strm0_ready         ( pe24__std__lane16_strm0_ready      ),      
               .std__pe24__lane16_strm0_cntl          ( std__pe24__lane16_strm0_cntl       ),      
               .std__pe24__lane16_strm0_data          ( std__pe24__lane16_strm0_data       ),      
               .std__pe24__lane16_strm0_data_valid    ( std__pe24__lane16_strm0_data_valid ),      
               .std__pe24__lane16_strm0_data_mask     ( std__pe24__lane16_strm0_data_mask  ),      

               .pe24__std__lane16_strm1_ready         ( pe24__std__lane16_strm1_ready      ),      
               .std__pe24__lane16_strm1_cntl          ( std__pe24__lane16_strm1_cntl       ),      
               .std__pe24__lane16_strm1_data          ( std__pe24__lane16_strm1_data       ),      
               .std__pe24__lane16_strm1_data_valid    ( std__pe24__lane16_strm1_data_valid ),      
               .std__pe24__lane16_strm1_data_mask     ( std__pe24__lane16_strm1_data_mask  ),      

               // PE 24, Lane 17                 
               .pe24__std__lane17_strm0_ready         ( pe24__std__lane17_strm0_ready      ),      
               .std__pe24__lane17_strm0_cntl          ( std__pe24__lane17_strm0_cntl       ),      
               .std__pe24__lane17_strm0_data          ( std__pe24__lane17_strm0_data       ),      
               .std__pe24__lane17_strm0_data_valid    ( std__pe24__lane17_strm0_data_valid ),      
               .std__pe24__lane17_strm0_data_mask     ( std__pe24__lane17_strm0_data_mask  ),      

               .pe24__std__lane17_strm1_ready         ( pe24__std__lane17_strm1_ready      ),      
               .std__pe24__lane17_strm1_cntl          ( std__pe24__lane17_strm1_cntl       ),      
               .std__pe24__lane17_strm1_data          ( std__pe24__lane17_strm1_data       ),      
               .std__pe24__lane17_strm1_data_valid    ( std__pe24__lane17_strm1_data_valid ),      
               .std__pe24__lane17_strm1_data_mask     ( std__pe24__lane17_strm1_data_mask  ),      

               // PE 24, Lane 18                 
               .pe24__std__lane18_strm0_ready         ( pe24__std__lane18_strm0_ready      ),      
               .std__pe24__lane18_strm0_cntl          ( std__pe24__lane18_strm0_cntl       ),      
               .std__pe24__lane18_strm0_data          ( std__pe24__lane18_strm0_data       ),      
               .std__pe24__lane18_strm0_data_valid    ( std__pe24__lane18_strm0_data_valid ),      
               .std__pe24__lane18_strm0_data_mask     ( std__pe24__lane18_strm0_data_mask  ),      

               .pe24__std__lane18_strm1_ready         ( pe24__std__lane18_strm1_ready      ),      
               .std__pe24__lane18_strm1_cntl          ( std__pe24__lane18_strm1_cntl       ),      
               .std__pe24__lane18_strm1_data          ( std__pe24__lane18_strm1_data       ),      
               .std__pe24__lane18_strm1_data_valid    ( std__pe24__lane18_strm1_data_valid ),      
               .std__pe24__lane18_strm1_data_mask     ( std__pe24__lane18_strm1_data_mask  ),      

               // PE 24, Lane 19                 
               .pe24__std__lane19_strm0_ready         ( pe24__std__lane19_strm0_ready      ),      
               .std__pe24__lane19_strm0_cntl          ( std__pe24__lane19_strm0_cntl       ),      
               .std__pe24__lane19_strm0_data          ( std__pe24__lane19_strm0_data       ),      
               .std__pe24__lane19_strm0_data_valid    ( std__pe24__lane19_strm0_data_valid ),      
               .std__pe24__lane19_strm0_data_mask     ( std__pe24__lane19_strm0_data_mask  ),      

               .pe24__std__lane19_strm1_ready         ( pe24__std__lane19_strm1_ready      ),      
               .std__pe24__lane19_strm1_cntl          ( std__pe24__lane19_strm1_cntl       ),      
               .std__pe24__lane19_strm1_data          ( std__pe24__lane19_strm1_data       ),      
               .std__pe24__lane19_strm1_data_valid    ( std__pe24__lane19_strm1_data_valid ),      
               .std__pe24__lane19_strm1_data_mask     ( std__pe24__lane19_strm1_data_mask  ),      

               // PE 24, Lane 20                 
               .pe24__std__lane20_strm0_ready         ( pe24__std__lane20_strm0_ready      ),      
               .std__pe24__lane20_strm0_cntl          ( std__pe24__lane20_strm0_cntl       ),      
               .std__pe24__lane20_strm0_data          ( std__pe24__lane20_strm0_data       ),      
               .std__pe24__lane20_strm0_data_valid    ( std__pe24__lane20_strm0_data_valid ),      
               .std__pe24__lane20_strm0_data_mask     ( std__pe24__lane20_strm0_data_mask  ),      

               .pe24__std__lane20_strm1_ready         ( pe24__std__lane20_strm1_ready      ),      
               .std__pe24__lane20_strm1_cntl          ( std__pe24__lane20_strm1_cntl       ),      
               .std__pe24__lane20_strm1_data          ( std__pe24__lane20_strm1_data       ),      
               .std__pe24__lane20_strm1_data_valid    ( std__pe24__lane20_strm1_data_valid ),      
               .std__pe24__lane20_strm1_data_mask     ( std__pe24__lane20_strm1_data_mask  ),      

               // PE 24, Lane 21                 
               .pe24__std__lane21_strm0_ready         ( pe24__std__lane21_strm0_ready      ),      
               .std__pe24__lane21_strm0_cntl          ( std__pe24__lane21_strm0_cntl       ),      
               .std__pe24__lane21_strm0_data          ( std__pe24__lane21_strm0_data       ),      
               .std__pe24__lane21_strm0_data_valid    ( std__pe24__lane21_strm0_data_valid ),      
               .std__pe24__lane21_strm0_data_mask     ( std__pe24__lane21_strm0_data_mask  ),      

               .pe24__std__lane21_strm1_ready         ( pe24__std__lane21_strm1_ready      ),      
               .std__pe24__lane21_strm1_cntl          ( std__pe24__lane21_strm1_cntl       ),      
               .std__pe24__lane21_strm1_data          ( std__pe24__lane21_strm1_data       ),      
               .std__pe24__lane21_strm1_data_valid    ( std__pe24__lane21_strm1_data_valid ),      
               .std__pe24__lane21_strm1_data_mask     ( std__pe24__lane21_strm1_data_mask  ),      

               // PE 24, Lane 22                 
               .pe24__std__lane22_strm0_ready         ( pe24__std__lane22_strm0_ready      ),      
               .std__pe24__lane22_strm0_cntl          ( std__pe24__lane22_strm0_cntl       ),      
               .std__pe24__lane22_strm0_data          ( std__pe24__lane22_strm0_data       ),      
               .std__pe24__lane22_strm0_data_valid    ( std__pe24__lane22_strm0_data_valid ),      
               .std__pe24__lane22_strm0_data_mask     ( std__pe24__lane22_strm0_data_mask  ),      

               .pe24__std__lane22_strm1_ready         ( pe24__std__lane22_strm1_ready      ),      
               .std__pe24__lane22_strm1_cntl          ( std__pe24__lane22_strm1_cntl       ),      
               .std__pe24__lane22_strm1_data          ( std__pe24__lane22_strm1_data       ),      
               .std__pe24__lane22_strm1_data_valid    ( std__pe24__lane22_strm1_data_valid ),      
               .std__pe24__lane22_strm1_data_mask     ( std__pe24__lane22_strm1_data_mask  ),      

               // PE 24, Lane 23                 
               .pe24__std__lane23_strm0_ready         ( pe24__std__lane23_strm0_ready      ),      
               .std__pe24__lane23_strm0_cntl          ( std__pe24__lane23_strm0_cntl       ),      
               .std__pe24__lane23_strm0_data          ( std__pe24__lane23_strm0_data       ),      
               .std__pe24__lane23_strm0_data_valid    ( std__pe24__lane23_strm0_data_valid ),      
               .std__pe24__lane23_strm0_data_mask     ( std__pe24__lane23_strm0_data_mask  ),      

               .pe24__std__lane23_strm1_ready         ( pe24__std__lane23_strm1_ready      ),      
               .std__pe24__lane23_strm1_cntl          ( std__pe24__lane23_strm1_cntl       ),      
               .std__pe24__lane23_strm1_data          ( std__pe24__lane23_strm1_data       ),      
               .std__pe24__lane23_strm1_data_valid    ( std__pe24__lane23_strm1_data_valid ),      
               .std__pe24__lane23_strm1_data_mask     ( std__pe24__lane23_strm1_data_mask  ),      

               // PE 24, Lane 24                 
               .pe24__std__lane24_strm0_ready         ( pe24__std__lane24_strm0_ready      ),      
               .std__pe24__lane24_strm0_cntl          ( std__pe24__lane24_strm0_cntl       ),      
               .std__pe24__lane24_strm0_data          ( std__pe24__lane24_strm0_data       ),      
               .std__pe24__lane24_strm0_data_valid    ( std__pe24__lane24_strm0_data_valid ),      
               .std__pe24__lane24_strm0_data_mask     ( std__pe24__lane24_strm0_data_mask  ),      

               .pe24__std__lane24_strm1_ready         ( pe24__std__lane24_strm1_ready      ),      
               .std__pe24__lane24_strm1_cntl          ( std__pe24__lane24_strm1_cntl       ),      
               .std__pe24__lane24_strm1_data          ( std__pe24__lane24_strm1_data       ),      
               .std__pe24__lane24_strm1_data_valid    ( std__pe24__lane24_strm1_data_valid ),      
               .std__pe24__lane24_strm1_data_mask     ( std__pe24__lane24_strm1_data_mask  ),      

               // PE 24, Lane 25                 
               .pe24__std__lane25_strm0_ready         ( pe24__std__lane25_strm0_ready      ),      
               .std__pe24__lane25_strm0_cntl          ( std__pe24__lane25_strm0_cntl       ),      
               .std__pe24__lane25_strm0_data          ( std__pe24__lane25_strm0_data       ),      
               .std__pe24__lane25_strm0_data_valid    ( std__pe24__lane25_strm0_data_valid ),      
               .std__pe24__lane25_strm0_data_mask     ( std__pe24__lane25_strm0_data_mask  ),      

               .pe24__std__lane25_strm1_ready         ( pe24__std__lane25_strm1_ready      ),      
               .std__pe24__lane25_strm1_cntl          ( std__pe24__lane25_strm1_cntl       ),      
               .std__pe24__lane25_strm1_data          ( std__pe24__lane25_strm1_data       ),      
               .std__pe24__lane25_strm1_data_valid    ( std__pe24__lane25_strm1_data_valid ),      
               .std__pe24__lane25_strm1_data_mask     ( std__pe24__lane25_strm1_data_mask  ),      

               // PE 24, Lane 26                 
               .pe24__std__lane26_strm0_ready         ( pe24__std__lane26_strm0_ready      ),      
               .std__pe24__lane26_strm0_cntl          ( std__pe24__lane26_strm0_cntl       ),      
               .std__pe24__lane26_strm0_data          ( std__pe24__lane26_strm0_data       ),      
               .std__pe24__lane26_strm0_data_valid    ( std__pe24__lane26_strm0_data_valid ),      
               .std__pe24__lane26_strm0_data_mask     ( std__pe24__lane26_strm0_data_mask  ),      

               .pe24__std__lane26_strm1_ready         ( pe24__std__lane26_strm1_ready      ),      
               .std__pe24__lane26_strm1_cntl          ( std__pe24__lane26_strm1_cntl       ),      
               .std__pe24__lane26_strm1_data          ( std__pe24__lane26_strm1_data       ),      
               .std__pe24__lane26_strm1_data_valid    ( std__pe24__lane26_strm1_data_valid ),      
               .std__pe24__lane26_strm1_data_mask     ( std__pe24__lane26_strm1_data_mask  ),      

               // PE 24, Lane 27                 
               .pe24__std__lane27_strm0_ready         ( pe24__std__lane27_strm0_ready      ),      
               .std__pe24__lane27_strm0_cntl          ( std__pe24__lane27_strm0_cntl       ),      
               .std__pe24__lane27_strm0_data          ( std__pe24__lane27_strm0_data       ),      
               .std__pe24__lane27_strm0_data_valid    ( std__pe24__lane27_strm0_data_valid ),      
               .std__pe24__lane27_strm0_data_mask     ( std__pe24__lane27_strm0_data_mask  ),      

               .pe24__std__lane27_strm1_ready         ( pe24__std__lane27_strm1_ready      ),      
               .std__pe24__lane27_strm1_cntl          ( std__pe24__lane27_strm1_cntl       ),      
               .std__pe24__lane27_strm1_data          ( std__pe24__lane27_strm1_data       ),      
               .std__pe24__lane27_strm1_data_valid    ( std__pe24__lane27_strm1_data_valid ),      
               .std__pe24__lane27_strm1_data_mask     ( std__pe24__lane27_strm1_data_mask  ),      

               // PE 24, Lane 28                 
               .pe24__std__lane28_strm0_ready         ( pe24__std__lane28_strm0_ready      ),      
               .std__pe24__lane28_strm0_cntl          ( std__pe24__lane28_strm0_cntl       ),      
               .std__pe24__lane28_strm0_data          ( std__pe24__lane28_strm0_data       ),      
               .std__pe24__lane28_strm0_data_valid    ( std__pe24__lane28_strm0_data_valid ),      
               .std__pe24__lane28_strm0_data_mask     ( std__pe24__lane28_strm0_data_mask  ),      

               .pe24__std__lane28_strm1_ready         ( pe24__std__lane28_strm1_ready      ),      
               .std__pe24__lane28_strm1_cntl          ( std__pe24__lane28_strm1_cntl       ),      
               .std__pe24__lane28_strm1_data          ( std__pe24__lane28_strm1_data       ),      
               .std__pe24__lane28_strm1_data_valid    ( std__pe24__lane28_strm1_data_valid ),      
               .std__pe24__lane28_strm1_data_mask     ( std__pe24__lane28_strm1_data_mask  ),      

               // PE 24, Lane 29                 
               .pe24__std__lane29_strm0_ready         ( pe24__std__lane29_strm0_ready      ),      
               .std__pe24__lane29_strm0_cntl          ( std__pe24__lane29_strm0_cntl       ),      
               .std__pe24__lane29_strm0_data          ( std__pe24__lane29_strm0_data       ),      
               .std__pe24__lane29_strm0_data_valid    ( std__pe24__lane29_strm0_data_valid ),      
               .std__pe24__lane29_strm0_data_mask     ( std__pe24__lane29_strm0_data_mask  ),      

               .pe24__std__lane29_strm1_ready         ( pe24__std__lane29_strm1_ready      ),      
               .std__pe24__lane29_strm1_cntl          ( std__pe24__lane29_strm1_cntl       ),      
               .std__pe24__lane29_strm1_data          ( std__pe24__lane29_strm1_data       ),      
               .std__pe24__lane29_strm1_data_valid    ( std__pe24__lane29_strm1_data_valid ),      
               .std__pe24__lane29_strm1_data_mask     ( std__pe24__lane29_strm1_data_mask  ),      

               // PE 24, Lane 30                 
               .pe24__std__lane30_strm0_ready         ( pe24__std__lane30_strm0_ready      ),      
               .std__pe24__lane30_strm0_cntl          ( std__pe24__lane30_strm0_cntl       ),      
               .std__pe24__lane30_strm0_data          ( std__pe24__lane30_strm0_data       ),      
               .std__pe24__lane30_strm0_data_valid    ( std__pe24__lane30_strm0_data_valid ),      
               .std__pe24__lane30_strm0_data_mask     ( std__pe24__lane30_strm0_data_mask  ),      

               .pe24__std__lane30_strm1_ready         ( pe24__std__lane30_strm1_ready      ),      
               .std__pe24__lane30_strm1_cntl          ( std__pe24__lane30_strm1_cntl       ),      
               .std__pe24__lane30_strm1_data          ( std__pe24__lane30_strm1_data       ),      
               .std__pe24__lane30_strm1_data_valid    ( std__pe24__lane30_strm1_data_valid ),      
               .std__pe24__lane30_strm1_data_mask     ( std__pe24__lane30_strm1_data_mask  ),      

               // PE 24, Lane 31                 
               .pe24__std__lane31_strm0_ready         ( pe24__std__lane31_strm0_ready      ),      
               .std__pe24__lane31_strm0_cntl          ( std__pe24__lane31_strm0_cntl       ),      
               .std__pe24__lane31_strm0_data          ( std__pe24__lane31_strm0_data       ),      
               .std__pe24__lane31_strm0_data_valid    ( std__pe24__lane31_strm0_data_valid ),      
               .std__pe24__lane31_strm0_data_mask     ( std__pe24__lane31_strm0_data_mask  ),      

               .pe24__std__lane31_strm1_ready         ( pe24__std__lane31_strm1_ready      ),      
               .std__pe24__lane31_strm1_cntl          ( std__pe24__lane31_strm1_cntl       ),      
               .std__pe24__lane31_strm1_data          ( std__pe24__lane31_strm1_data       ),      
               .std__pe24__lane31_strm1_data_valid    ( std__pe24__lane31_strm1_data_valid ),      
               .std__pe24__lane31_strm1_data_mask     ( std__pe24__lane31_strm1_data_mask  ),      

               // PE 25, Lane 0                 
               .pe25__std__lane0_strm0_ready         ( pe25__std__lane0_strm0_ready      ),      
               .std__pe25__lane0_strm0_cntl          ( std__pe25__lane0_strm0_cntl       ),      
               .std__pe25__lane0_strm0_data          ( std__pe25__lane0_strm0_data       ),      
               .std__pe25__lane0_strm0_data_valid    ( std__pe25__lane0_strm0_data_valid ),      
               .std__pe25__lane0_strm0_data_mask     ( std__pe25__lane0_strm0_data_mask  ),      

               .pe25__std__lane0_strm1_ready         ( pe25__std__lane0_strm1_ready      ),      
               .std__pe25__lane0_strm1_cntl          ( std__pe25__lane0_strm1_cntl       ),      
               .std__pe25__lane0_strm1_data          ( std__pe25__lane0_strm1_data       ),      
               .std__pe25__lane0_strm1_data_valid    ( std__pe25__lane0_strm1_data_valid ),      
               .std__pe25__lane0_strm1_data_mask     ( std__pe25__lane0_strm1_data_mask  ),      

               // PE 25, Lane 1                 
               .pe25__std__lane1_strm0_ready         ( pe25__std__lane1_strm0_ready      ),      
               .std__pe25__lane1_strm0_cntl          ( std__pe25__lane1_strm0_cntl       ),      
               .std__pe25__lane1_strm0_data          ( std__pe25__lane1_strm0_data       ),      
               .std__pe25__lane1_strm0_data_valid    ( std__pe25__lane1_strm0_data_valid ),      
               .std__pe25__lane1_strm0_data_mask     ( std__pe25__lane1_strm0_data_mask  ),      

               .pe25__std__lane1_strm1_ready         ( pe25__std__lane1_strm1_ready      ),      
               .std__pe25__lane1_strm1_cntl          ( std__pe25__lane1_strm1_cntl       ),      
               .std__pe25__lane1_strm1_data          ( std__pe25__lane1_strm1_data       ),      
               .std__pe25__lane1_strm1_data_valid    ( std__pe25__lane1_strm1_data_valid ),      
               .std__pe25__lane1_strm1_data_mask     ( std__pe25__lane1_strm1_data_mask  ),      

               // PE 25, Lane 2                 
               .pe25__std__lane2_strm0_ready         ( pe25__std__lane2_strm0_ready      ),      
               .std__pe25__lane2_strm0_cntl          ( std__pe25__lane2_strm0_cntl       ),      
               .std__pe25__lane2_strm0_data          ( std__pe25__lane2_strm0_data       ),      
               .std__pe25__lane2_strm0_data_valid    ( std__pe25__lane2_strm0_data_valid ),      
               .std__pe25__lane2_strm0_data_mask     ( std__pe25__lane2_strm0_data_mask  ),      

               .pe25__std__lane2_strm1_ready         ( pe25__std__lane2_strm1_ready      ),      
               .std__pe25__lane2_strm1_cntl          ( std__pe25__lane2_strm1_cntl       ),      
               .std__pe25__lane2_strm1_data          ( std__pe25__lane2_strm1_data       ),      
               .std__pe25__lane2_strm1_data_valid    ( std__pe25__lane2_strm1_data_valid ),      
               .std__pe25__lane2_strm1_data_mask     ( std__pe25__lane2_strm1_data_mask  ),      

               // PE 25, Lane 3                 
               .pe25__std__lane3_strm0_ready         ( pe25__std__lane3_strm0_ready      ),      
               .std__pe25__lane3_strm0_cntl          ( std__pe25__lane3_strm0_cntl       ),      
               .std__pe25__lane3_strm0_data          ( std__pe25__lane3_strm0_data       ),      
               .std__pe25__lane3_strm0_data_valid    ( std__pe25__lane3_strm0_data_valid ),      
               .std__pe25__lane3_strm0_data_mask     ( std__pe25__lane3_strm0_data_mask  ),      

               .pe25__std__lane3_strm1_ready         ( pe25__std__lane3_strm1_ready      ),      
               .std__pe25__lane3_strm1_cntl          ( std__pe25__lane3_strm1_cntl       ),      
               .std__pe25__lane3_strm1_data          ( std__pe25__lane3_strm1_data       ),      
               .std__pe25__lane3_strm1_data_valid    ( std__pe25__lane3_strm1_data_valid ),      
               .std__pe25__lane3_strm1_data_mask     ( std__pe25__lane3_strm1_data_mask  ),      

               // PE 25, Lane 4                 
               .pe25__std__lane4_strm0_ready         ( pe25__std__lane4_strm0_ready      ),      
               .std__pe25__lane4_strm0_cntl          ( std__pe25__lane4_strm0_cntl       ),      
               .std__pe25__lane4_strm0_data          ( std__pe25__lane4_strm0_data       ),      
               .std__pe25__lane4_strm0_data_valid    ( std__pe25__lane4_strm0_data_valid ),      
               .std__pe25__lane4_strm0_data_mask     ( std__pe25__lane4_strm0_data_mask  ),      

               .pe25__std__lane4_strm1_ready         ( pe25__std__lane4_strm1_ready      ),      
               .std__pe25__lane4_strm1_cntl          ( std__pe25__lane4_strm1_cntl       ),      
               .std__pe25__lane4_strm1_data          ( std__pe25__lane4_strm1_data       ),      
               .std__pe25__lane4_strm1_data_valid    ( std__pe25__lane4_strm1_data_valid ),      
               .std__pe25__lane4_strm1_data_mask     ( std__pe25__lane4_strm1_data_mask  ),      

               // PE 25, Lane 5                 
               .pe25__std__lane5_strm0_ready         ( pe25__std__lane5_strm0_ready      ),      
               .std__pe25__lane5_strm0_cntl          ( std__pe25__lane5_strm0_cntl       ),      
               .std__pe25__lane5_strm0_data          ( std__pe25__lane5_strm0_data       ),      
               .std__pe25__lane5_strm0_data_valid    ( std__pe25__lane5_strm0_data_valid ),      
               .std__pe25__lane5_strm0_data_mask     ( std__pe25__lane5_strm0_data_mask  ),      

               .pe25__std__lane5_strm1_ready         ( pe25__std__lane5_strm1_ready      ),      
               .std__pe25__lane5_strm1_cntl          ( std__pe25__lane5_strm1_cntl       ),      
               .std__pe25__lane5_strm1_data          ( std__pe25__lane5_strm1_data       ),      
               .std__pe25__lane5_strm1_data_valid    ( std__pe25__lane5_strm1_data_valid ),      
               .std__pe25__lane5_strm1_data_mask     ( std__pe25__lane5_strm1_data_mask  ),      

               // PE 25, Lane 6                 
               .pe25__std__lane6_strm0_ready         ( pe25__std__lane6_strm0_ready      ),      
               .std__pe25__lane6_strm0_cntl          ( std__pe25__lane6_strm0_cntl       ),      
               .std__pe25__lane6_strm0_data          ( std__pe25__lane6_strm0_data       ),      
               .std__pe25__lane6_strm0_data_valid    ( std__pe25__lane6_strm0_data_valid ),      
               .std__pe25__lane6_strm0_data_mask     ( std__pe25__lane6_strm0_data_mask  ),      

               .pe25__std__lane6_strm1_ready         ( pe25__std__lane6_strm1_ready      ),      
               .std__pe25__lane6_strm1_cntl          ( std__pe25__lane6_strm1_cntl       ),      
               .std__pe25__lane6_strm1_data          ( std__pe25__lane6_strm1_data       ),      
               .std__pe25__lane6_strm1_data_valid    ( std__pe25__lane6_strm1_data_valid ),      
               .std__pe25__lane6_strm1_data_mask     ( std__pe25__lane6_strm1_data_mask  ),      

               // PE 25, Lane 7                 
               .pe25__std__lane7_strm0_ready         ( pe25__std__lane7_strm0_ready      ),      
               .std__pe25__lane7_strm0_cntl          ( std__pe25__lane7_strm0_cntl       ),      
               .std__pe25__lane7_strm0_data          ( std__pe25__lane7_strm0_data       ),      
               .std__pe25__lane7_strm0_data_valid    ( std__pe25__lane7_strm0_data_valid ),      
               .std__pe25__lane7_strm0_data_mask     ( std__pe25__lane7_strm0_data_mask  ),      

               .pe25__std__lane7_strm1_ready         ( pe25__std__lane7_strm1_ready      ),      
               .std__pe25__lane7_strm1_cntl          ( std__pe25__lane7_strm1_cntl       ),      
               .std__pe25__lane7_strm1_data          ( std__pe25__lane7_strm1_data       ),      
               .std__pe25__lane7_strm1_data_valid    ( std__pe25__lane7_strm1_data_valid ),      
               .std__pe25__lane7_strm1_data_mask     ( std__pe25__lane7_strm1_data_mask  ),      

               // PE 25, Lane 8                 
               .pe25__std__lane8_strm0_ready         ( pe25__std__lane8_strm0_ready      ),      
               .std__pe25__lane8_strm0_cntl          ( std__pe25__lane8_strm0_cntl       ),      
               .std__pe25__lane8_strm0_data          ( std__pe25__lane8_strm0_data       ),      
               .std__pe25__lane8_strm0_data_valid    ( std__pe25__lane8_strm0_data_valid ),      
               .std__pe25__lane8_strm0_data_mask     ( std__pe25__lane8_strm0_data_mask  ),      

               .pe25__std__lane8_strm1_ready         ( pe25__std__lane8_strm1_ready      ),      
               .std__pe25__lane8_strm1_cntl          ( std__pe25__lane8_strm1_cntl       ),      
               .std__pe25__lane8_strm1_data          ( std__pe25__lane8_strm1_data       ),      
               .std__pe25__lane8_strm1_data_valid    ( std__pe25__lane8_strm1_data_valid ),      
               .std__pe25__lane8_strm1_data_mask     ( std__pe25__lane8_strm1_data_mask  ),      

               // PE 25, Lane 9                 
               .pe25__std__lane9_strm0_ready         ( pe25__std__lane9_strm0_ready      ),      
               .std__pe25__lane9_strm0_cntl          ( std__pe25__lane9_strm0_cntl       ),      
               .std__pe25__lane9_strm0_data          ( std__pe25__lane9_strm0_data       ),      
               .std__pe25__lane9_strm0_data_valid    ( std__pe25__lane9_strm0_data_valid ),      
               .std__pe25__lane9_strm0_data_mask     ( std__pe25__lane9_strm0_data_mask  ),      

               .pe25__std__lane9_strm1_ready         ( pe25__std__lane9_strm1_ready      ),      
               .std__pe25__lane9_strm1_cntl          ( std__pe25__lane9_strm1_cntl       ),      
               .std__pe25__lane9_strm1_data          ( std__pe25__lane9_strm1_data       ),      
               .std__pe25__lane9_strm1_data_valid    ( std__pe25__lane9_strm1_data_valid ),      
               .std__pe25__lane9_strm1_data_mask     ( std__pe25__lane9_strm1_data_mask  ),      

               // PE 25, Lane 10                 
               .pe25__std__lane10_strm0_ready         ( pe25__std__lane10_strm0_ready      ),      
               .std__pe25__lane10_strm0_cntl          ( std__pe25__lane10_strm0_cntl       ),      
               .std__pe25__lane10_strm0_data          ( std__pe25__lane10_strm0_data       ),      
               .std__pe25__lane10_strm0_data_valid    ( std__pe25__lane10_strm0_data_valid ),      
               .std__pe25__lane10_strm0_data_mask     ( std__pe25__lane10_strm0_data_mask  ),      

               .pe25__std__lane10_strm1_ready         ( pe25__std__lane10_strm1_ready      ),      
               .std__pe25__lane10_strm1_cntl          ( std__pe25__lane10_strm1_cntl       ),      
               .std__pe25__lane10_strm1_data          ( std__pe25__lane10_strm1_data       ),      
               .std__pe25__lane10_strm1_data_valid    ( std__pe25__lane10_strm1_data_valid ),      
               .std__pe25__lane10_strm1_data_mask     ( std__pe25__lane10_strm1_data_mask  ),      

               // PE 25, Lane 11                 
               .pe25__std__lane11_strm0_ready         ( pe25__std__lane11_strm0_ready      ),      
               .std__pe25__lane11_strm0_cntl          ( std__pe25__lane11_strm0_cntl       ),      
               .std__pe25__lane11_strm0_data          ( std__pe25__lane11_strm0_data       ),      
               .std__pe25__lane11_strm0_data_valid    ( std__pe25__lane11_strm0_data_valid ),      
               .std__pe25__lane11_strm0_data_mask     ( std__pe25__lane11_strm0_data_mask  ),      

               .pe25__std__lane11_strm1_ready         ( pe25__std__lane11_strm1_ready      ),      
               .std__pe25__lane11_strm1_cntl          ( std__pe25__lane11_strm1_cntl       ),      
               .std__pe25__lane11_strm1_data          ( std__pe25__lane11_strm1_data       ),      
               .std__pe25__lane11_strm1_data_valid    ( std__pe25__lane11_strm1_data_valid ),      
               .std__pe25__lane11_strm1_data_mask     ( std__pe25__lane11_strm1_data_mask  ),      

               // PE 25, Lane 12                 
               .pe25__std__lane12_strm0_ready         ( pe25__std__lane12_strm0_ready      ),      
               .std__pe25__lane12_strm0_cntl          ( std__pe25__lane12_strm0_cntl       ),      
               .std__pe25__lane12_strm0_data          ( std__pe25__lane12_strm0_data       ),      
               .std__pe25__lane12_strm0_data_valid    ( std__pe25__lane12_strm0_data_valid ),      
               .std__pe25__lane12_strm0_data_mask     ( std__pe25__lane12_strm0_data_mask  ),      

               .pe25__std__lane12_strm1_ready         ( pe25__std__lane12_strm1_ready      ),      
               .std__pe25__lane12_strm1_cntl          ( std__pe25__lane12_strm1_cntl       ),      
               .std__pe25__lane12_strm1_data          ( std__pe25__lane12_strm1_data       ),      
               .std__pe25__lane12_strm1_data_valid    ( std__pe25__lane12_strm1_data_valid ),      
               .std__pe25__lane12_strm1_data_mask     ( std__pe25__lane12_strm1_data_mask  ),      

               // PE 25, Lane 13                 
               .pe25__std__lane13_strm0_ready         ( pe25__std__lane13_strm0_ready      ),      
               .std__pe25__lane13_strm0_cntl          ( std__pe25__lane13_strm0_cntl       ),      
               .std__pe25__lane13_strm0_data          ( std__pe25__lane13_strm0_data       ),      
               .std__pe25__lane13_strm0_data_valid    ( std__pe25__lane13_strm0_data_valid ),      
               .std__pe25__lane13_strm0_data_mask     ( std__pe25__lane13_strm0_data_mask  ),      

               .pe25__std__lane13_strm1_ready         ( pe25__std__lane13_strm1_ready      ),      
               .std__pe25__lane13_strm1_cntl          ( std__pe25__lane13_strm1_cntl       ),      
               .std__pe25__lane13_strm1_data          ( std__pe25__lane13_strm1_data       ),      
               .std__pe25__lane13_strm1_data_valid    ( std__pe25__lane13_strm1_data_valid ),      
               .std__pe25__lane13_strm1_data_mask     ( std__pe25__lane13_strm1_data_mask  ),      

               // PE 25, Lane 14                 
               .pe25__std__lane14_strm0_ready         ( pe25__std__lane14_strm0_ready      ),      
               .std__pe25__lane14_strm0_cntl          ( std__pe25__lane14_strm0_cntl       ),      
               .std__pe25__lane14_strm0_data          ( std__pe25__lane14_strm0_data       ),      
               .std__pe25__lane14_strm0_data_valid    ( std__pe25__lane14_strm0_data_valid ),      
               .std__pe25__lane14_strm0_data_mask     ( std__pe25__lane14_strm0_data_mask  ),      

               .pe25__std__lane14_strm1_ready         ( pe25__std__lane14_strm1_ready      ),      
               .std__pe25__lane14_strm1_cntl          ( std__pe25__lane14_strm1_cntl       ),      
               .std__pe25__lane14_strm1_data          ( std__pe25__lane14_strm1_data       ),      
               .std__pe25__lane14_strm1_data_valid    ( std__pe25__lane14_strm1_data_valid ),      
               .std__pe25__lane14_strm1_data_mask     ( std__pe25__lane14_strm1_data_mask  ),      

               // PE 25, Lane 15                 
               .pe25__std__lane15_strm0_ready         ( pe25__std__lane15_strm0_ready      ),      
               .std__pe25__lane15_strm0_cntl          ( std__pe25__lane15_strm0_cntl       ),      
               .std__pe25__lane15_strm0_data          ( std__pe25__lane15_strm0_data       ),      
               .std__pe25__lane15_strm0_data_valid    ( std__pe25__lane15_strm0_data_valid ),      
               .std__pe25__lane15_strm0_data_mask     ( std__pe25__lane15_strm0_data_mask  ),      

               .pe25__std__lane15_strm1_ready         ( pe25__std__lane15_strm1_ready      ),      
               .std__pe25__lane15_strm1_cntl          ( std__pe25__lane15_strm1_cntl       ),      
               .std__pe25__lane15_strm1_data          ( std__pe25__lane15_strm1_data       ),      
               .std__pe25__lane15_strm1_data_valid    ( std__pe25__lane15_strm1_data_valid ),      
               .std__pe25__lane15_strm1_data_mask     ( std__pe25__lane15_strm1_data_mask  ),      

               // PE 25, Lane 16                 
               .pe25__std__lane16_strm0_ready         ( pe25__std__lane16_strm0_ready      ),      
               .std__pe25__lane16_strm0_cntl          ( std__pe25__lane16_strm0_cntl       ),      
               .std__pe25__lane16_strm0_data          ( std__pe25__lane16_strm0_data       ),      
               .std__pe25__lane16_strm0_data_valid    ( std__pe25__lane16_strm0_data_valid ),      
               .std__pe25__lane16_strm0_data_mask     ( std__pe25__lane16_strm0_data_mask  ),      

               .pe25__std__lane16_strm1_ready         ( pe25__std__lane16_strm1_ready      ),      
               .std__pe25__lane16_strm1_cntl          ( std__pe25__lane16_strm1_cntl       ),      
               .std__pe25__lane16_strm1_data          ( std__pe25__lane16_strm1_data       ),      
               .std__pe25__lane16_strm1_data_valid    ( std__pe25__lane16_strm1_data_valid ),      
               .std__pe25__lane16_strm1_data_mask     ( std__pe25__lane16_strm1_data_mask  ),      

               // PE 25, Lane 17                 
               .pe25__std__lane17_strm0_ready         ( pe25__std__lane17_strm0_ready      ),      
               .std__pe25__lane17_strm0_cntl          ( std__pe25__lane17_strm0_cntl       ),      
               .std__pe25__lane17_strm0_data          ( std__pe25__lane17_strm0_data       ),      
               .std__pe25__lane17_strm0_data_valid    ( std__pe25__lane17_strm0_data_valid ),      
               .std__pe25__lane17_strm0_data_mask     ( std__pe25__lane17_strm0_data_mask  ),      

               .pe25__std__lane17_strm1_ready         ( pe25__std__lane17_strm1_ready      ),      
               .std__pe25__lane17_strm1_cntl          ( std__pe25__lane17_strm1_cntl       ),      
               .std__pe25__lane17_strm1_data          ( std__pe25__lane17_strm1_data       ),      
               .std__pe25__lane17_strm1_data_valid    ( std__pe25__lane17_strm1_data_valid ),      
               .std__pe25__lane17_strm1_data_mask     ( std__pe25__lane17_strm1_data_mask  ),      

               // PE 25, Lane 18                 
               .pe25__std__lane18_strm0_ready         ( pe25__std__lane18_strm0_ready      ),      
               .std__pe25__lane18_strm0_cntl          ( std__pe25__lane18_strm0_cntl       ),      
               .std__pe25__lane18_strm0_data          ( std__pe25__lane18_strm0_data       ),      
               .std__pe25__lane18_strm0_data_valid    ( std__pe25__lane18_strm0_data_valid ),      
               .std__pe25__lane18_strm0_data_mask     ( std__pe25__lane18_strm0_data_mask  ),      

               .pe25__std__lane18_strm1_ready         ( pe25__std__lane18_strm1_ready      ),      
               .std__pe25__lane18_strm1_cntl          ( std__pe25__lane18_strm1_cntl       ),      
               .std__pe25__lane18_strm1_data          ( std__pe25__lane18_strm1_data       ),      
               .std__pe25__lane18_strm1_data_valid    ( std__pe25__lane18_strm1_data_valid ),      
               .std__pe25__lane18_strm1_data_mask     ( std__pe25__lane18_strm1_data_mask  ),      

               // PE 25, Lane 19                 
               .pe25__std__lane19_strm0_ready         ( pe25__std__lane19_strm0_ready      ),      
               .std__pe25__lane19_strm0_cntl          ( std__pe25__lane19_strm0_cntl       ),      
               .std__pe25__lane19_strm0_data          ( std__pe25__lane19_strm0_data       ),      
               .std__pe25__lane19_strm0_data_valid    ( std__pe25__lane19_strm0_data_valid ),      
               .std__pe25__lane19_strm0_data_mask     ( std__pe25__lane19_strm0_data_mask  ),      

               .pe25__std__lane19_strm1_ready         ( pe25__std__lane19_strm1_ready      ),      
               .std__pe25__lane19_strm1_cntl          ( std__pe25__lane19_strm1_cntl       ),      
               .std__pe25__lane19_strm1_data          ( std__pe25__lane19_strm1_data       ),      
               .std__pe25__lane19_strm1_data_valid    ( std__pe25__lane19_strm1_data_valid ),      
               .std__pe25__lane19_strm1_data_mask     ( std__pe25__lane19_strm1_data_mask  ),      

               // PE 25, Lane 20                 
               .pe25__std__lane20_strm0_ready         ( pe25__std__lane20_strm0_ready      ),      
               .std__pe25__lane20_strm0_cntl          ( std__pe25__lane20_strm0_cntl       ),      
               .std__pe25__lane20_strm0_data          ( std__pe25__lane20_strm0_data       ),      
               .std__pe25__lane20_strm0_data_valid    ( std__pe25__lane20_strm0_data_valid ),      
               .std__pe25__lane20_strm0_data_mask     ( std__pe25__lane20_strm0_data_mask  ),      

               .pe25__std__lane20_strm1_ready         ( pe25__std__lane20_strm1_ready      ),      
               .std__pe25__lane20_strm1_cntl          ( std__pe25__lane20_strm1_cntl       ),      
               .std__pe25__lane20_strm1_data          ( std__pe25__lane20_strm1_data       ),      
               .std__pe25__lane20_strm1_data_valid    ( std__pe25__lane20_strm1_data_valid ),      
               .std__pe25__lane20_strm1_data_mask     ( std__pe25__lane20_strm1_data_mask  ),      

               // PE 25, Lane 21                 
               .pe25__std__lane21_strm0_ready         ( pe25__std__lane21_strm0_ready      ),      
               .std__pe25__lane21_strm0_cntl          ( std__pe25__lane21_strm0_cntl       ),      
               .std__pe25__lane21_strm0_data          ( std__pe25__lane21_strm0_data       ),      
               .std__pe25__lane21_strm0_data_valid    ( std__pe25__lane21_strm0_data_valid ),      
               .std__pe25__lane21_strm0_data_mask     ( std__pe25__lane21_strm0_data_mask  ),      

               .pe25__std__lane21_strm1_ready         ( pe25__std__lane21_strm1_ready      ),      
               .std__pe25__lane21_strm1_cntl          ( std__pe25__lane21_strm1_cntl       ),      
               .std__pe25__lane21_strm1_data          ( std__pe25__lane21_strm1_data       ),      
               .std__pe25__lane21_strm1_data_valid    ( std__pe25__lane21_strm1_data_valid ),      
               .std__pe25__lane21_strm1_data_mask     ( std__pe25__lane21_strm1_data_mask  ),      

               // PE 25, Lane 22                 
               .pe25__std__lane22_strm0_ready         ( pe25__std__lane22_strm0_ready      ),      
               .std__pe25__lane22_strm0_cntl          ( std__pe25__lane22_strm0_cntl       ),      
               .std__pe25__lane22_strm0_data          ( std__pe25__lane22_strm0_data       ),      
               .std__pe25__lane22_strm0_data_valid    ( std__pe25__lane22_strm0_data_valid ),      
               .std__pe25__lane22_strm0_data_mask     ( std__pe25__lane22_strm0_data_mask  ),      

               .pe25__std__lane22_strm1_ready         ( pe25__std__lane22_strm1_ready      ),      
               .std__pe25__lane22_strm1_cntl          ( std__pe25__lane22_strm1_cntl       ),      
               .std__pe25__lane22_strm1_data          ( std__pe25__lane22_strm1_data       ),      
               .std__pe25__lane22_strm1_data_valid    ( std__pe25__lane22_strm1_data_valid ),      
               .std__pe25__lane22_strm1_data_mask     ( std__pe25__lane22_strm1_data_mask  ),      

               // PE 25, Lane 23                 
               .pe25__std__lane23_strm0_ready         ( pe25__std__lane23_strm0_ready      ),      
               .std__pe25__lane23_strm0_cntl          ( std__pe25__lane23_strm0_cntl       ),      
               .std__pe25__lane23_strm0_data          ( std__pe25__lane23_strm0_data       ),      
               .std__pe25__lane23_strm0_data_valid    ( std__pe25__lane23_strm0_data_valid ),      
               .std__pe25__lane23_strm0_data_mask     ( std__pe25__lane23_strm0_data_mask  ),      

               .pe25__std__lane23_strm1_ready         ( pe25__std__lane23_strm1_ready      ),      
               .std__pe25__lane23_strm1_cntl          ( std__pe25__lane23_strm1_cntl       ),      
               .std__pe25__lane23_strm1_data          ( std__pe25__lane23_strm1_data       ),      
               .std__pe25__lane23_strm1_data_valid    ( std__pe25__lane23_strm1_data_valid ),      
               .std__pe25__lane23_strm1_data_mask     ( std__pe25__lane23_strm1_data_mask  ),      

               // PE 25, Lane 24                 
               .pe25__std__lane24_strm0_ready         ( pe25__std__lane24_strm0_ready      ),      
               .std__pe25__lane24_strm0_cntl          ( std__pe25__lane24_strm0_cntl       ),      
               .std__pe25__lane24_strm0_data          ( std__pe25__lane24_strm0_data       ),      
               .std__pe25__lane24_strm0_data_valid    ( std__pe25__lane24_strm0_data_valid ),      
               .std__pe25__lane24_strm0_data_mask     ( std__pe25__lane24_strm0_data_mask  ),      

               .pe25__std__lane24_strm1_ready         ( pe25__std__lane24_strm1_ready      ),      
               .std__pe25__lane24_strm1_cntl          ( std__pe25__lane24_strm1_cntl       ),      
               .std__pe25__lane24_strm1_data          ( std__pe25__lane24_strm1_data       ),      
               .std__pe25__lane24_strm1_data_valid    ( std__pe25__lane24_strm1_data_valid ),      
               .std__pe25__lane24_strm1_data_mask     ( std__pe25__lane24_strm1_data_mask  ),      

               // PE 25, Lane 25                 
               .pe25__std__lane25_strm0_ready         ( pe25__std__lane25_strm0_ready      ),      
               .std__pe25__lane25_strm0_cntl          ( std__pe25__lane25_strm0_cntl       ),      
               .std__pe25__lane25_strm0_data          ( std__pe25__lane25_strm0_data       ),      
               .std__pe25__lane25_strm0_data_valid    ( std__pe25__lane25_strm0_data_valid ),      
               .std__pe25__lane25_strm0_data_mask     ( std__pe25__lane25_strm0_data_mask  ),      

               .pe25__std__lane25_strm1_ready         ( pe25__std__lane25_strm1_ready      ),      
               .std__pe25__lane25_strm1_cntl          ( std__pe25__lane25_strm1_cntl       ),      
               .std__pe25__lane25_strm1_data          ( std__pe25__lane25_strm1_data       ),      
               .std__pe25__lane25_strm1_data_valid    ( std__pe25__lane25_strm1_data_valid ),      
               .std__pe25__lane25_strm1_data_mask     ( std__pe25__lane25_strm1_data_mask  ),      

               // PE 25, Lane 26                 
               .pe25__std__lane26_strm0_ready         ( pe25__std__lane26_strm0_ready      ),      
               .std__pe25__lane26_strm0_cntl          ( std__pe25__lane26_strm0_cntl       ),      
               .std__pe25__lane26_strm0_data          ( std__pe25__lane26_strm0_data       ),      
               .std__pe25__lane26_strm0_data_valid    ( std__pe25__lane26_strm0_data_valid ),      
               .std__pe25__lane26_strm0_data_mask     ( std__pe25__lane26_strm0_data_mask  ),      

               .pe25__std__lane26_strm1_ready         ( pe25__std__lane26_strm1_ready      ),      
               .std__pe25__lane26_strm1_cntl          ( std__pe25__lane26_strm1_cntl       ),      
               .std__pe25__lane26_strm1_data          ( std__pe25__lane26_strm1_data       ),      
               .std__pe25__lane26_strm1_data_valid    ( std__pe25__lane26_strm1_data_valid ),      
               .std__pe25__lane26_strm1_data_mask     ( std__pe25__lane26_strm1_data_mask  ),      

               // PE 25, Lane 27                 
               .pe25__std__lane27_strm0_ready         ( pe25__std__lane27_strm0_ready      ),      
               .std__pe25__lane27_strm0_cntl          ( std__pe25__lane27_strm0_cntl       ),      
               .std__pe25__lane27_strm0_data          ( std__pe25__lane27_strm0_data       ),      
               .std__pe25__lane27_strm0_data_valid    ( std__pe25__lane27_strm0_data_valid ),      
               .std__pe25__lane27_strm0_data_mask     ( std__pe25__lane27_strm0_data_mask  ),      

               .pe25__std__lane27_strm1_ready         ( pe25__std__lane27_strm1_ready      ),      
               .std__pe25__lane27_strm1_cntl          ( std__pe25__lane27_strm1_cntl       ),      
               .std__pe25__lane27_strm1_data          ( std__pe25__lane27_strm1_data       ),      
               .std__pe25__lane27_strm1_data_valid    ( std__pe25__lane27_strm1_data_valid ),      
               .std__pe25__lane27_strm1_data_mask     ( std__pe25__lane27_strm1_data_mask  ),      

               // PE 25, Lane 28                 
               .pe25__std__lane28_strm0_ready         ( pe25__std__lane28_strm0_ready      ),      
               .std__pe25__lane28_strm0_cntl          ( std__pe25__lane28_strm0_cntl       ),      
               .std__pe25__lane28_strm0_data          ( std__pe25__lane28_strm0_data       ),      
               .std__pe25__lane28_strm0_data_valid    ( std__pe25__lane28_strm0_data_valid ),      
               .std__pe25__lane28_strm0_data_mask     ( std__pe25__lane28_strm0_data_mask  ),      

               .pe25__std__lane28_strm1_ready         ( pe25__std__lane28_strm1_ready      ),      
               .std__pe25__lane28_strm1_cntl          ( std__pe25__lane28_strm1_cntl       ),      
               .std__pe25__lane28_strm1_data          ( std__pe25__lane28_strm1_data       ),      
               .std__pe25__lane28_strm1_data_valid    ( std__pe25__lane28_strm1_data_valid ),      
               .std__pe25__lane28_strm1_data_mask     ( std__pe25__lane28_strm1_data_mask  ),      

               // PE 25, Lane 29                 
               .pe25__std__lane29_strm0_ready         ( pe25__std__lane29_strm0_ready      ),      
               .std__pe25__lane29_strm0_cntl          ( std__pe25__lane29_strm0_cntl       ),      
               .std__pe25__lane29_strm0_data          ( std__pe25__lane29_strm0_data       ),      
               .std__pe25__lane29_strm0_data_valid    ( std__pe25__lane29_strm0_data_valid ),      
               .std__pe25__lane29_strm0_data_mask     ( std__pe25__lane29_strm0_data_mask  ),      

               .pe25__std__lane29_strm1_ready         ( pe25__std__lane29_strm1_ready      ),      
               .std__pe25__lane29_strm1_cntl          ( std__pe25__lane29_strm1_cntl       ),      
               .std__pe25__lane29_strm1_data          ( std__pe25__lane29_strm1_data       ),      
               .std__pe25__lane29_strm1_data_valid    ( std__pe25__lane29_strm1_data_valid ),      
               .std__pe25__lane29_strm1_data_mask     ( std__pe25__lane29_strm1_data_mask  ),      

               // PE 25, Lane 30                 
               .pe25__std__lane30_strm0_ready         ( pe25__std__lane30_strm0_ready      ),      
               .std__pe25__lane30_strm0_cntl          ( std__pe25__lane30_strm0_cntl       ),      
               .std__pe25__lane30_strm0_data          ( std__pe25__lane30_strm0_data       ),      
               .std__pe25__lane30_strm0_data_valid    ( std__pe25__lane30_strm0_data_valid ),      
               .std__pe25__lane30_strm0_data_mask     ( std__pe25__lane30_strm0_data_mask  ),      

               .pe25__std__lane30_strm1_ready         ( pe25__std__lane30_strm1_ready      ),      
               .std__pe25__lane30_strm1_cntl          ( std__pe25__lane30_strm1_cntl       ),      
               .std__pe25__lane30_strm1_data          ( std__pe25__lane30_strm1_data       ),      
               .std__pe25__lane30_strm1_data_valid    ( std__pe25__lane30_strm1_data_valid ),      
               .std__pe25__lane30_strm1_data_mask     ( std__pe25__lane30_strm1_data_mask  ),      

               // PE 25, Lane 31                 
               .pe25__std__lane31_strm0_ready         ( pe25__std__lane31_strm0_ready      ),      
               .std__pe25__lane31_strm0_cntl          ( std__pe25__lane31_strm0_cntl       ),      
               .std__pe25__lane31_strm0_data          ( std__pe25__lane31_strm0_data       ),      
               .std__pe25__lane31_strm0_data_valid    ( std__pe25__lane31_strm0_data_valid ),      
               .std__pe25__lane31_strm0_data_mask     ( std__pe25__lane31_strm0_data_mask  ),      

               .pe25__std__lane31_strm1_ready         ( pe25__std__lane31_strm1_ready      ),      
               .std__pe25__lane31_strm1_cntl          ( std__pe25__lane31_strm1_cntl       ),      
               .std__pe25__lane31_strm1_data          ( std__pe25__lane31_strm1_data       ),      
               .std__pe25__lane31_strm1_data_valid    ( std__pe25__lane31_strm1_data_valid ),      
               .std__pe25__lane31_strm1_data_mask     ( std__pe25__lane31_strm1_data_mask  ),      

               // PE 26, Lane 0                 
               .pe26__std__lane0_strm0_ready         ( pe26__std__lane0_strm0_ready      ),      
               .std__pe26__lane0_strm0_cntl          ( std__pe26__lane0_strm0_cntl       ),      
               .std__pe26__lane0_strm0_data          ( std__pe26__lane0_strm0_data       ),      
               .std__pe26__lane0_strm0_data_valid    ( std__pe26__lane0_strm0_data_valid ),      
               .std__pe26__lane0_strm0_data_mask     ( std__pe26__lane0_strm0_data_mask  ),      

               .pe26__std__lane0_strm1_ready         ( pe26__std__lane0_strm1_ready      ),      
               .std__pe26__lane0_strm1_cntl          ( std__pe26__lane0_strm1_cntl       ),      
               .std__pe26__lane0_strm1_data          ( std__pe26__lane0_strm1_data       ),      
               .std__pe26__lane0_strm1_data_valid    ( std__pe26__lane0_strm1_data_valid ),      
               .std__pe26__lane0_strm1_data_mask     ( std__pe26__lane0_strm1_data_mask  ),      

               // PE 26, Lane 1                 
               .pe26__std__lane1_strm0_ready         ( pe26__std__lane1_strm0_ready      ),      
               .std__pe26__lane1_strm0_cntl          ( std__pe26__lane1_strm0_cntl       ),      
               .std__pe26__lane1_strm0_data          ( std__pe26__lane1_strm0_data       ),      
               .std__pe26__lane1_strm0_data_valid    ( std__pe26__lane1_strm0_data_valid ),      
               .std__pe26__lane1_strm0_data_mask     ( std__pe26__lane1_strm0_data_mask  ),      

               .pe26__std__lane1_strm1_ready         ( pe26__std__lane1_strm1_ready      ),      
               .std__pe26__lane1_strm1_cntl          ( std__pe26__lane1_strm1_cntl       ),      
               .std__pe26__lane1_strm1_data          ( std__pe26__lane1_strm1_data       ),      
               .std__pe26__lane1_strm1_data_valid    ( std__pe26__lane1_strm1_data_valid ),      
               .std__pe26__lane1_strm1_data_mask     ( std__pe26__lane1_strm1_data_mask  ),      

               // PE 26, Lane 2                 
               .pe26__std__lane2_strm0_ready         ( pe26__std__lane2_strm0_ready      ),      
               .std__pe26__lane2_strm0_cntl          ( std__pe26__lane2_strm0_cntl       ),      
               .std__pe26__lane2_strm0_data          ( std__pe26__lane2_strm0_data       ),      
               .std__pe26__lane2_strm0_data_valid    ( std__pe26__lane2_strm0_data_valid ),      
               .std__pe26__lane2_strm0_data_mask     ( std__pe26__lane2_strm0_data_mask  ),      

               .pe26__std__lane2_strm1_ready         ( pe26__std__lane2_strm1_ready      ),      
               .std__pe26__lane2_strm1_cntl          ( std__pe26__lane2_strm1_cntl       ),      
               .std__pe26__lane2_strm1_data          ( std__pe26__lane2_strm1_data       ),      
               .std__pe26__lane2_strm1_data_valid    ( std__pe26__lane2_strm1_data_valid ),      
               .std__pe26__lane2_strm1_data_mask     ( std__pe26__lane2_strm1_data_mask  ),      

               // PE 26, Lane 3                 
               .pe26__std__lane3_strm0_ready         ( pe26__std__lane3_strm0_ready      ),      
               .std__pe26__lane3_strm0_cntl          ( std__pe26__lane3_strm0_cntl       ),      
               .std__pe26__lane3_strm0_data          ( std__pe26__lane3_strm0_data       ),      
               .std__pe26__lane3_strm0_data_valid    ( std__pe26__lane3_strm0_data_valid ),      
               .std__pe26__lane3_strm0_data_mask     ( std__pe26__lane3_strm0_data_mask  ),      

               .pe26__std__lane3_strm1_ready         ( pe26__std__lane3_strm1_ready      ),      
               .std__pe26__lane3_strm1_cntl          ( std__pe26__lane3_strm1_cntl       ),      
               .std__pe26__lane3_strm1_data          ( std__pe26__lane3_strm1_data       ),      
               .std__pe26__lane3_strm1_data_valid    ( std__pe26__lane3_strm1_data_valid ),      
               .std__pe26__lane3_strm1_data_mask     ( std__pe26__lane3_strm1_data_mask  ),      

               // PE 26, Lane 4                 
               .pe26__std__lane4_strm0_ready         ( pe26__std__lane4_strm0_ready      ),      
               .std__pe26__lane4_strm0_cntl          ( std__pe26__lane4_strm0_cntl       ),      
               .std__pe26__lane4_strm0_data          ( std__pe26__lane4_strm0_data       ),      
               .std__pe26__lane4_strm0_data_valid    ( std__pe26__lane4_strm0_data_valid ),      
               .std__pe26__lane4_strm0_data_mask     ( std__pe26__lane4_strm0_data_mask  ),      

               .pe26__std__lane4_strm1_ready         ( pe26__std__lane4_strm1_ready      ),      
               .std__pe26__lane4_strm1_cntl          ( std__pe26__lane4_strm1_cntl       ),      
               .std__pe26__lane4_strm1_data          ( std__pe26__lane4_strm1_data       ),      
               .std__pe26__lane4_strm1_data_valid    ( std__pe26__lane4_strm1_data_valid ),      
               .std__pe26__lane4_strm1_data_mask     ( std__pe26__lane4_strm1_data_mask  ),      

               // PE 26, Lane 5                 
               .pe26__std__lane5_strm0_ready         ( pe26__std__lane5_strm0_ready      ),      
               .std__pe26__lane5_strm0_cntl          ( std__pe26__lane5_strm0_cntl       ),      
               .std__pe26__lane5_strm0_data          ( std__pe26__lane5_strm0_data       ),      
               .std__pe26__lane5_strm0_data_valid    ( std__pe26__lane5_strm0_data_valid ),      
               .std__pe26__lane5_strm0_data_mask     ( std__pe26__lane5_strm0_data_mask  ),      

               .pe26__std__lane5_strm1_ready         ( pe26__std__lane5_strm1_ready      ),      
               .std__pe26__lane5_strm1_cntl          ( std__pe26__lane5_strm1_cntl       ),      
               .std__pe26__lane5_strm1_data          ( std__pe26__lane5_strm1_data       ),      
               .std__pe26__lane5_strm1_data_valid    ( std__pe26__lane5_strm1_data_valid ),      
               .std__pe26__lane5_strm1_data_mask     ( std__pe26__lane5_strm1_data_mask  ),      

               // PE 26, Lane 6                 
               .pe26__std__lane6_strm0_ready         ( pe26__std__lane6_strm0_ready      ),      
               .std__pe26__lane6_strm0_cntl          ( std__pe26__lane6_strm0_cntl       ),      
               .std__pe26__lane6_strm0_data          ( std__pe26__lane6_strm0_data       ),      
               .std__pe26__lane6_strm0_data_valid    ( std__pe26__lane6_strm0_data_valid ),      
               .std__pe26__lane6_strm0_data_mask     ( std__pe26__lane6_strm0_data_mask  ),      

               .pe26__std__lane6_strm1_ready         ( pe26__std__lane6_strm1_ready      ),      
               .std__pe26__lane6_strm1_cntl          ( std__pe26__lane6_strm1_cntl       ),      
               .std__pe26__lane6_strm1_data          ( std__pe26__lane6_strm1_data       ),      
               .std__pe26__lane6_strm1_data_valid    ( std__pe26__lane6_strm1_data_valid ),      
               .std__pe26__lane6_strm1_data_mask     ( std__pe26__lane6_strm1_data_mask  ),      

               // PE 26, Lane 7                 
               .pe26__std__lane7_strm0_ready         ( pe26__std__lane7_strm0_ready      ),      
               .std__pe26__lane7_strm0_cntl          ( std__pe26__lane7_strm0_cntl       ),      
               .std__pe26__lane7_strm0_data          ( std__pe26__lane7_strm0_data       ),      
               .std__pe26__lane7_strm0_data_valid    ( std__pe26__lane7_strm0_data_valid ),      
               .std__pe26__lane7_strm0_data_mask     ( std__pe26__lane7_strm0_data_mask  ),      

               .pe26__std__lane7_strm1_ready         ( pe26__std__lane7_strm1_ready      ),      
               .std__pe26__lane7_strm1_cntl          ( std__pe26__lane7_strm1_cntl       ),      
               .std__pe26__lane7_strm1_data          ( std__pe26__lane7_strm1_data       ),      
               .std__pe26__lane7_strm1_data_valid    ( std__pe26__lane7_strm1_data_valid ),      
               .std__pe26__lane7_strm1_data_mask     ( std__pe26__lane7_strm1_data_mask  ),      

               // PE 26, Lane 8                 
               .pe26__std__lane8_strm0_ready         ( pe26__std__lane8_strm0_ready      ),      
               .std__pe26__lane8_strm0_cntl          ( std__pe26__lane8_strm0_cntl       ),      
               .std__pe26__lane8_strm0_data          ( std__pe26__lane8_strm0_data       ),      
               .std__pe26__lane8_strm0_data_valid    ( std__pe26__lane8_strm0_data_valid ),      
               .std__pe26__lane8_strm0_data_mask     ( std__pe26__lane8_strm0_data_mask  ),      

               .pe26__std__lane8_strm1_ready         ( pe26__std__lane8_strm1_ready      ),      
               .std__pe26__lane8_strm1_cntl          ( std__pe26__lane8_strm1_cntl       ),      
               .std__pe26__lane8_strm1_data          ( std__pe26__lane8_strm1_data       ),      
               .std__pe26__lane8_strm1_data_valid    ( std__pe26__lane8_strm1_data_valid ),      
               .std__pe26__lane8_strm1_data_mask     ( std__pe26__lane8_strm1_data_mask  ),      

               // PE 26, Lane 9                 
               .pe26__std__lane9_strm0_ready         ( pe26__std__lane9_strm0_ready      ),      
               .std__pe26__lane9_strm0_cntl          ( std__pe26__lane9_strm0_cntl       ),      
               .std__pe26__lane9_strm0_data          ( std__pe26__lane9_strm0_data       ),      
               .std__pe26__lane9_strm0_data_valid    ( std__pe26__lane9_strm0_data_valid ),      
               .std__pe26__lane9_strm0_data_mask     ( std__pe26__lane9_strm0_data_mask  ),      

               .pe26__std__lane9_strm1_ready         ( pe26__std__lane9_strm1_ready      ),      
               .std__pe26__lane9_strm1_cntl          ( std__pe26__lane9_strm1_cntl       ),      
               .std__pe26__lane9_strm1_data          ( std__pe26__lane9_strm1_data       ),      
               .std__pe26__lane9_strm1_data_valid    ( std__pe26__lane9_strm1_data_valid ),      
               .std__pe26__lane9_strm1_data_mask     ( std__pe26__lane9_strm1_data_mask  ),      

               // PE 26, Lane 10                 
               .pe26__std__lane10_strm0_ready         ( pe26__std__lane10_strm0_ready      ),      
               .std__pe26__lane10_strm0_cntl          ( std__pe26__lane10_strm0_cntl       ),      
               .std__pe26__lane10_strm0_data          ( std__pe26__lane10_strm0_data       ),      
               .std__pe26__lane10_strm0_data_valid    ( std__pe26__lane10_strm0_data_valid ),      
               .std__pe26__lane10_strm0_data_mask     ( std__pe26__lane10_strm0_data_mask  ),      

               .pe26__std__lane10_strm1_ready         ( pe26__std__lane10_strm1_ready      ),      
               .std__pe26__lane10_strm1_cntl          ( std__pe26__lane10_strm1_cntl       ),      
               .std__pe26__lane10_strm1_data          ( std__pe26__lane10_strm1_data       ),      
               .std__pe26__lane10_strm1_data_valid    ( std__pe26__lane10_strm1_data_valid ),      
               .std__pe26__lane10_strm1_data_mask     ( std__pe26__lane10_strm1_data_mask  ),      

               // PE 26, Lane 11                 
               .pe26__std__lane11_strm0_ready         ( pe26__std__lane11_strm0_ready      ),      
               .std__pe26__lane11_strm0_cntl          ( std__pe26__lane11_strm0_cntl       ),      
               .std__pe26__lane11_strm0_data          ( std__pe26__lane11_strm0_data       ),      
               .std__pe26__lane11_strm0_data_valid    ( std__pe26__lane11_strm0_data_valid ),      
               .std__pe26__lane11_strm0_data_mask     ( std__pe26__lane11_strm0_data_mask  ),      

               .pe26__std__lane11_strm1_ready         ( pe26__std__lane11_strm1_ready      ),      
               .std__pe26__lane11_strm1_cntl          ( std__pe26__lane11_strm1_cntl       ),      
               .std__pe26__lane11_strm1_data          ( std__pe26__lane11_strm1_data       ),      
               .std__pe26__lane11_strm1_data_valid    ( std__pe26__lane11_strm1_data_valid ),      
               .std__pe26__lane11_strm1_data_mask     ( std__pe26__lane11_strm1_data_mask  ),      

               // PE 26, Lane 12                 
               .pe26__std__lane12_strm0_ready         ( pe26__std__lane12_strm0_ready      ),      
               .std__pe26__lane12_strm0_cntl          ( std__pe26__lane12_strm0_cntl       ),      
               .std__pe26__lane12_strm0_data          ( std__pe26__lane12_strm0_data       ),      
               .std__pe26__lane12_strm0_data_valid    ( std__pe26__lane12_strm0_data_valid ),      
               .std__pe26__lane12_strm0_data_mask     ( std__pe26__lane12_strm0_data_mask  ),      

               .pe26__std__lane12_strm1_ready         ( pe26__std__lane12_strm1_ready      ),      
               .std__pe26__lane12_strm1_cntl          ( std__pe26__lane12_strm1_cntl       ),      
               .std__pe26__lane12_strm1_data          ( std__pe26__lane12_strm1_data       ),      
               .std__pe26__lane12_strm1_data_valid    ( std__pe26__lane12_strm1_data_valid ),      
               .std__pe26__lane12_strm1_data_mask     ( std__pe26__lane12_strm1_data_mask  ),      

               // PE 26, Lane 13                 
               .pe26__std__lane13_strm0_ready         ( pe26__std__lane13_strm0_ready      ),      
               .std__pe26__lane13_strm0_cntl          ( std__pe26__lane13_strm0_cntl       ),      
               .std__pe26__lane13_strm0_data          ( std__pe26__lane13_strm0_data       ),      
               .std__pe26__lane13_strm0_data_valid    ( std__pe26__lane13_strm0_data_valid ),      
               .std__pe26__lane13_strm0_data_mask     ( std__pe26__lane13_strm0_data_mask  ),      

               .pe26__std__lane13_strm1_ready         ( pe26__std__lane13_strm1_ready      ),      
               .std__pe26__lane13_strm1_cntl          ( std__pe26__lane13_strm1_cntl       ),      
               .std__pe26__lane13_strm1_data          ( std__pe26__lane13_strm1_data       ),      
               .std__pe26__lane13_strm1_data_valid    ( std__pe26__lane13_strm1_data_valid ),      
               .std__pe26__lane13_strm1_data_mask     ( std__pe26__lane13_strm1_data_mask  ),      

               // PE 26, Lane 14                 
               .pe26__std__lane14_strm0_ready         ( pe26__std__lane14_strm0_ready      ),      
               .std__pe26__lane14_strm0_cntl          ( std__pe26__lane14_strm0_cntl       ),      
               .std__pe26__lane14_strm0_data          ( std__pe26__lane14_strm0_data       ),      
               .std__pe26__lane14_strm0_data_valid    ( std__pe26__lane14_strm0_data_valid ),      
               .std__pe26__lane14_strm0_data_mask     ( std__pe26__lane14_strm0_data_mask  ),      

               .pe26__std__lane14_strm1_ready         ( pe26__std__lane14_strm1_ready      ),      
               .std__pe26__lane14_strm1_cntl          ( std__pe26__lane14_strm1_cntl       ),      
               .std__pe26__lane14_strm1_data          ( std__pe26__lane14_strm1_data       ),      
               .std__pe26__lane14_strm1_data_valid    ( std__pe26__lane14_strm1_data_valid ),      
               .std__pe26__lane14_strm1_data_mask     ( std__pe26__lane14_strm1_data_mask  ),      

               // PE 26, Lane 15                 
               .pe26__std__lane15_strm0_ready         ( pe26__std__lane15_strm0_ready      ),      
               .std__pe26__lane15_strm0_cntl          ( std__pe26__lane15_strm0_cntl       ),      
               .std__pe26__lane15_strm0_data          ( std__pe26__lane15_strm0_data       ),      
               .std__pe26__lane15_strm0_data_valid    ( std__pe26__lane15_strm0_data_valid ),      
               .std__pe26__lane15_strm0_data_mask     ( std__pe26__lane15_strm0_data_mask  ),      

               .pe26__std__lane15_strm1_ready         ( pe26__std__lane15_strm1_ready      ),      
               .std__pe26__lane15_strm1_cntl          ( std__pe26__lane15_strm1_cntl       ),      
               .std__pe26__lane15_strm1_data          ( std__pe26__lane15_strm1_data       ),      
               .std__pe26__lane15_strm1_data_valid    ( std__pe26__lane15_strm1_data_valid ),      
               .std__pe26__lane15_strm1_data_mask     ( std__pe26__lane15_strm1_data_mask  ),      

               // PE 26, Lane 16                 
               .pe26__std__lane16_strm0_ready         ( pe26__std__lane16_strm0_ready      ),      
               .std__pe26__lane16_strm0_cntl          ( std__pe26__lane16_strm0_cntl       ),      
               .std__pe26__lane16_strm0_data          ( std__pe26__lane16_strm0_data       ),      
               .std__pe26__lane16_strm0_data_valid    ( std__pe26__lane16_strm0_data_valid ),      
               .std__pe26__lane16_strm0_data_mask     ( std__pe26__lane16_strm0_data_mask  ),      

               .pe26__std__lane16_strm1_ready         ( pe26__std__lane16_strm1_ready      ),      
               .std__pe26__lane16_strm1_cntl          ( std__pe26__lane16_strm1_cntl       ),      
               .std__pe26__lane16_strm1_data          ( std__pe26__lane16_strm1_data       ),      
               .std__pe26__lane16_strm1_data_valid    ( std__pe26__lane16_strm1_data_valid ),      
               .std__pe26__lane16_strm1_data_mask     ( std__pe26__lane16_strm1_data_mask  ),      

               // PE 26, Lane 17                 
               .pe26__std__lane17_strm0_ready         ( pe26__std__lane17_strm0_ready      ),      
               .std__pe26__lane17_strm0_cntl          ( std__pe26__lane17_strm0_cntl       ),      
               .std__pe26__lane17_strm0_data          ( std__pe26__lane17_strm0_data       ),      
               .std__pe26__lane17_strm0_data_valid    ( std__pe26__lane17_strm0_data_valid ),      
               .std__pe26__lane17_strm0_data_mask     ( std__pe26__lane17_strm0_data_mask  ),      

               .pe26__std__lane17_strm1_ready         ( pe26__std__lane17_strm1_ready      ),      
               .std__pe26__lane17_strm1_cntl          ( std__pe26__lane17_strm1_cntl       ),      
               .std__pe26__lane17_strm1_data          ( std__pe26__lane17_strm1_data       ),      
               .std__pe26__lane17_strm1_data_valid    ( std__pe26__lane17_strm1_data_valid ),      
               .std__pe26__lane17_strm1_data_mask     ( std__pe26__lane17_strm1_data_mask  ),      

               // PE 26, Lane 18                 
               .pe26__std__lane18_strm0_ready         ( pe26__std__lane18_strm0_ready      ),      
               .std__pe26__lane18_strm0_cntl          ( std__pe26__lane18_strm0_cntl       ),      
               .std__pe26__lane18_strm0_data          ( std__pe26__lane18_strm0_data       ),      
               .std__pe26__lane18_strm0_data_valid    ( std__pe26__lane18_strm0_data_valid ),      
               .std__pe26__lane18_strm0_data_mask     ( std__pe26__lane18_strm0_data_mask  ),      

               .pe26__std__lane18_strm1_ready         ( pe26__std__lane18_strm1_ready      ),      
               .std__pe26__lane18_strm1_cntl          ( std__pe26__lane18_strm1_cntl       ),      
               .std__pe26__lane18_strm1_data          ( std__pe26__lane18_strm1_data       ),      
               .std__pe26__lane18_strm1_data_valid    ( std__pe26__lane18_strm1_data_valid ),      
               .std__pe26__lane18_strm1_data_mask     ( std__pe26__lane18_strm1_data_mask  ),      

               // PE 26, Lane 19                 
               .pe26__std__lane19_strm0_ready         ( pe26__std__lane19_strm0_ready      ),      
               .std__pe26__lane19_strm0_cntl          ( std__pe26__lane19_strm0_cntl       ),      
               .std__pe26__lane19_strm0_data          ( std__pe26__lane19_strm0_data       ),      
               .std__pe26__lane19_strm0_data_valid    ( std__pe26__lane19_strm0_data_valid ),      
               .std__pe26__lane19_strm0_data_mask     ( std__pe26__lane19_strm0_data_mask  ),      

               .pe26__std__lane19_strm1_ready         ( pe26__std__lane19_strm1_ready      ),      
               .std__pe26__lane19_strm1_cntl          ( std__pe26__lane19_strm1_cntl       ),      
               .std__pe26__lane19_strm1_data          ( std__pe26__lane19_strm1_data       ),      
               .std__pe26__lane19_strm1_data_valid    ( std__pe26__lane19_strm1_data_valid ),      
               .std__pe26__lane19_strm1_data_mask     ( std__pe26__lane19_strm1_data_mask  ),      

               // PE 26, Lane 20                 
               .pe26__std__lane20_strm0_ready         ( pe26__std__lane20_strm0_ready      ),      
               .std__pe26__lane20_strm0_cntl          ( std__pe26__lane20_strm0_cntl       ),      
               .std__pe26__lane20_strm0_data          ( std__pe26__lane20_strm0_data       ),      
               .std__pe26__lane20_strm0_data_valid    ( std__pe26__lane20_strm0_data_valid ),      
               .std__pe26__lane20_strm0_data_mask     ( std__pe26__lane20_strm0_data_mask  ),      

               .pe26__std__lane20_strm1_ready         ( pe26__std__lane20_strm1_ready      ),      
               .std__pe26__lane20_strm1_cntl          ( std__pe26__lane20_strm1_cntl       ),      
               .std__pe26__lane20_strm1_data          ( std__pe26__lane20_strm1_data       ),      
               .std__pe26__lane20_strm1_data_valid    ( std__pe26__lane20_strm1_data_valid ),      
               .std__pe26__lane20_strm1_data_mask     ( std__pe26__lane20_strm1_data_mask  ),      

               // PE 26, Lane 21                 
               .pe26__std__lane21_strm0_ready         ( pe26__std__lane21_strm0_ready      ),      
               .std__pe26__lane21_strm0_cntl          ( std__pe26__lane21_strm0_cntl       ),      
               .std__pe26__lane21_strm0_data          ( std__pe26__lane21_strm0_data       ),      
               .std__pe26__lane21_strm0_data_valid    ( std__pe26__lane21_strm0_data_valid ),      
               .std__pe26__lane21_strm0_data_mask     ( std__pe26__lane21_strm0_data_mask  ),      

               .pe26__std__lane21_strm1_ready         ( pe26__std__lane21_strm1_ready      ),      
               .std__pe26__lane21_strm1_cntl          ( std__pe26__lane21_strm1_cntl       ),      
               .std__pe26__lane21_strm1_data          ( std__pe26__lane21_strm1_data       ),      
               .std__pe26__lane21_strm1_data_valid    ( std__pe26__lane21_strm1_data_valid ),      
               .std__pe26__lane21_strm1_data_mask     ( std__pe26__lane21_strm1_data_mask  ),      

               // PE 26, Lane 22                 
               .pe26__std__lane22_strm0_ready         ( pe26__std__lane22_strm0_ready      ),      
               .std__pe26__lane22_strm0_cntl          ( std__pe26__lane22_strm0_cntl       ),      
               .std__pe26__lane22_strm0_data          ( std__pe26__lane22_strm0_data       ),      
               .std__pe26__lane22_strm0_data_valid    ( std__pe26__lane22_strm0_data_valid ),      
               .std__pe26__lane22_strm0_data_mask     ( std__pe26__lane22_strm0_data_mask  ),      

               .pe26__std__lane22_strm1_ready         ( pe26__std__lane22_strm1_ready      ),      
               .std__pe26__lane22_strm1_cntl          ( std__pe26__lane22_strm1_cntl       ),      
               .std__pe26__lane22_strm1_data          ( std__pe26__lane22_strm1_data       ),      
               .std__pe26__lane22_strm1_data_valid    ( std__pe26__lane22_strm1_data_valid ),      
               .std__pe26__lane22_strm1_data_mask     ( std__pe26__lane22_strm1_data_mask  ),      

               // PE 26, Lane 23                 
               .pe26__std__lane23_strm0_ready         ( pe26__std__lane23_strm0_ready      ),      
               .std__pe26__lane23_strm0_cntl          ( std__pe26__lane23_strm0_cntl       ),      
               .std__pe26__lane23_strm0_data          ( std__pe26__lane23_strm0_data       ),      
               .std__pe26__lane23_strm0_data_valid    ( std__pe26__lane23_strm0_data_valid ),      
               .std__pe26__lane23_strm0_data_mask     ( std__pe26__lane23_strm0_data_mask  ),      

               .pe26__std__lane23_strm1_ready         ( pe26__std__lane23_strm1_ready      ),      
               .std__pe26__lane23_strm1_cntl          ( std__pe26__lane23_strm1_cntl       ),      
               .std__pe26__lane23_strm1_data          ( std__pe26__lane23_strm1_data       ),      
               .std__pe26__lane23_strm1_data_valid    ( std__pe26__lane23_strm1_data_valid ),      
               .std__pe26__lane23_strm1_data_mask     ( std__pe26__lane23_strm1_data_mask  ),      

               // PE 26, Lane 24                 
               .pe26__std__lane24_strm0_ready         ( pe26__std__lane24_strm0_ready      ),      
               .std__pe26__lane24_strm0_cntl          ( std__pe26__lane24_strm0_cntl       ),      
               .std__pe26__lane24_strm0_data          ( std__pe26__lane24_strm0_data       ),      
               .std__pe26__lane24_strm0_data_valid    ( std__pe26__lane24_strm0_data_valid ),      
               .std__pe26__lane24_strm0_data_mask     ( std__pe26__lane24_strm0_data_mask  ),      

               .pe26__std__lane24_strm1_ready         ( pe26__std__lane24_strm1_ready      ),      
               .std__pe26__lane24_strm1_cntl          ( std__pe26__lane24_strm1_cntl       ),      
               .std__pe26__lane24_strm1_data          ( std__pe26__lane24_strm1_data       ),      
               .std__pe26__lane24_strm1_data_valid    ( std__pe26__lane24_strm1_data_valid ),      
               .std__pe26__lane24_strm1_data_mask     ( std__pe26__lane24_strm1_data_mask  ),      

               // PE 26, Lane 25                 
               .pe26__std__lane25_strm0_ready         ( pe26__std__lane25_strm0_ready      ),      
               .std__pe26__lane25_strm0_cntl          ( std__pe26__lane25_strm0_cntl       ),      
               .std__pe26__lane25_strm0_data          ( std__pe26__lane25_strm0_data       ),      
               .std__pe26__lane25_strm0_data_valid    ( std__pe26__lane25_strm0_data_valid ),      
               .std__pe26__lane25_strm0_data_mask     ( std__pe26__lane25_strm0_data_mask  ),      

               .pe26__std__lane25_strm1_ready         ( pe26__std__lane25_strm1_ready      ),      
               .std__pe26__lane25_strm1_cntl          ( std__pe26__lane25_strm1_cntl       ),      
               .std__pe26__lane25_strm1_data          ( std__pe26__lane25_strm1_data       ),      
               .std__pe26__lane25_strm1_data_valid    ( std__pe26__lane25_strm1_data_valid ),      
               .std__pe26__lane25_strm1_data_mask     ( std__pe26__lane25_strm1_data_mask  ),      

               // PE 26, Lane 26                 
               .pe26__std__lane26_strm0_ready         ( pe26__std__lane26_strm0_ready      ),      
               .std__pe26__lane26_strm0_cntl          ( std__pe26__lane26_strm0_cntl       ),      
               .std__pe26__lane26_strm0_data          ( std__pe26__lane26_strm0_data       ),      
               .std__pe26__lane26_strm0_data_valid    ( std__pe26__lane26_strm0_data_valid ),      
               .std__pe26__lane26_strm0_data_mask     ( std__pe26__lane26_strm0_data_mask  ),      

               .pe26__std__lane26_strm1_ready         ( pe26__std__lane26_strm1_ready      ),      
               .std__pe26__lane26_strm1_cntl          ( std__pe26__lane26_strm1_cntl       ),      
               .std__pe26__lane26_strm1_data          ( std__pe26__lane26_strm1_data       ),      
               .std__pe26__lane26_strm1_data_valid    ( std__pe26__lane26_strm1_data_valid ),      
               .std__pe26__lane26_strm1_data_mask     ( std__pe26__lane26_strm1_data_mask  ),      

               // PE 26, Lane 27                 
               .pe26__std__lane27_strm0_ready         ( pe26__std__lane27_strm0_ready      ),      
               .std__pe26__lane27_strm0_cntl          ( std__pe26__lane27_strm0_cntl       ),      
               .std__pe26__lane27_strm0_data          ( std__pe26__lane27_strm0_data       ),      
               .std__pe26__lane27_strm0_data_valid    ( std__pe26__lane27_strm0_data_valid ),      
               .std__pe26__lane27_strm0_data_mask     ( std__pe26__lane27_strm0_data_mask  ),      

               .pe26__std__lane27_strm1_ready         ( pe26__std__lane27_strm1_ready      ),      
               .std__pe26__lane27_strm1_cntl          ( std__pe26__lane27_strm1_cntl       ),      
               .std__pe26__lane27_strm1_data          ( std__pe26__lane27_strm1_data       ),      
               .std__pe26__lane27_strm1_data_valid    ( std__pe26__lane27_strm1_data_valid ),      
               .std__pe26__lane27_strm1_data_mask     ( std__pe26__lane27_strm1_data_mask  ),      

               // PE 26, Lane 28                 
               .pe26__std__lane28_strm0_ready         ( pe26__std__lane28_strm0_ready      ),      
               .std__pe26__lane28_strm0_cntl          ( std__pe26__lane28_strm0_cntl       ),      
               .std__pe26__lane28_strm0_data          ( std__pe26__lane28_strm0_data       ),      
               .std__pe26__lane28_strm0_data_valid    ( std__pe26__lane28_strm0_data_valid ),      
               .std__pe26__lane28_strm0_data_mask     ( std__pe26__lane28_strm0_data_mask  ),      

               .pe26__std__lane28_strm1_ready         ( pe26__std__lane28_strm1_ready      ),      
               .std__pe26__lane28_strm1_cntl          ( std__pe26__lane28_strm1_cntl       ),      
               .std__pe26__lane28_strm1_data          ( std__pe26__lane28_strm1_data       ),      
               .std__pe26__lane28_strm1_data_valid    ( std__pe26__lane28_strm1_data_valid ),      
               .std__pe26__lane28_strm1_data_mask     ( std__pe26__lane28_strm1_data_mask  ),      

               // PE 26, Lane 29                 
               .pe26__std__lane29_strm0_ready         ( pe26__std__lane29_strm0_ready      ),      
               .std__pe26__lane29_strm0_cntl          ( std__pe26__lane29_strm0_cntl       ),      
               .std__pe26__lane29_strm0_data          ( std__pe26__lane29_strm0_data       ),      
               .std__pe26__lane29_strm0_data_valid    ( std__pe26__lane29_strm0_data_valid ),      
               .std__pe26__lane29_strm0_data_mask     ( std__pe26__lane29_strm0_data_mask  ),      

               .pe26__std__lane29_strm1_ready         ( pe26__std__lane29_strm1_ready      ),      
               .std__pe26__lane29_strm1_cntl          ( std__pe26__lane29_strm1_cntl       ),      
               .std__pe26__lane29_strm1_data          ( std__pe26__lane29_strm1_data       ),      
               .std__pe26__lane29_strm1_data_valid    ( std__pe26__lane29_strm1_data_valid ),      
               .std__pe26__lane29_strm1_data_mask     ( std__pe26__lane29_strm1_data_mask  ),      

               // PE 26, Lane 30                 
               .pe26__std__lane30_strm0_ready         ( pe26__std__lane30_strm0_ready      ),      
               .std__pe26__lane30_strm0_cntl          ( std__pe26__lane30_strm0_cntl       ),      
               .std__pe26__lane30_strm0_data          ( std__pe26__lane30_strm0_data       ),      
               .std__pe26__lane30_strm0_data_valid    ( std__pe26__lane30_strm0_data_valid ),      
               .std__pe26__lane30_strm0_data_mask     ( std__pe26__lane30_strm0_data_mask  ),      

               .pe26__std__lane30_strm1_ready         ( pe26__std__lane30_strm1_ready      ),      
               .std__pe26__lane30_strm1_cntl          ( std__pe26__lane30_strm1_cntl       ),      
               .std__pe26__lane30_strm1_data          ( std__pe26__lane30_strm1_data       ),      
               .std__pe26__lane30_strm1_data_valid    ( std__pe26__lane30_strm1_data_valid ),      
               .std__pe26__lane30_strm1_data_mask     ( std__pe26__lane30_strm1_data_mask  ),      

               // PE 26, Lane 31                 
               .pe26__std__lane31_strm0_ready         ( pe26__std__lane31_strm0_ready      ),      
               .std__pe26__lane31_strm0_cntl          ( std__pe26__lane31_strm0_cntl       ),      
               .std__pe26__lane31_strm0_data          ( std__pe26__lane31_strm0_data       ),      
               .std__pe26__lane31_strm0_data_valid    ( std__pe26__lane31_strm0_data_valid ),      
               .std__pe26__lane31_strm0_data_mask     ( std__pe26__lane31_strm0_data_mask  ),      

               .pe26__std__lane31_strm1_ready         ( pe26__std__lane31_strm1_ready      ),      
               .std__pe26__lane31_strm1_cntl          ( std__pe26__lane31_strm1_cntl       ),      
               .std__pe26__lane31_strm1_data          ( std__pe26__lane31_strm1_data       ),      
               .std__pe26__lane31_strm1_data_valid    ( std__pe26__lane31_strm1_data_valid ),      
               .std__pe26__lane31_strm1_data_mask     ( std__pe26__lane31_strm1_data_mask  ),      

               // PE 27, Lane 0                 
               .pe27__std__lane0_strm0_ready         ( pe27__std__lane0_strm0_ready      ),      
               .std__pe27__lane0_strm0_cntl          ( std__pe27__lane0_strm0_cntl       ),      
               .std__pe27__lane0_strm0_data          ( std__pe27__lane0_strm0_data       ),      
               .std__pe27__lane0_strm0_data_valid    ( std__pe27__lane0_strm0_data_valid ),      
               .std__pe27__lane0_strm0_data_mask     ( std__pe27__lane0_strm0_data_mask  ),      

               .pe27__std__lane0_strm1_ready         ( pe27__std__lane0_strm1_ready      ),      
               .std__pe27__lane0_strm1_cntl          ( std__pe27__lane0_strm1_cntl       ),      
               .std__pe27__lane0_strm1_data          ( std__pe27__lane0_strm1_data       ),      
               .std__pe27__lane0_strm1_data_valid    ( std__pe27__lane0_strm1_data_valid ),      
               .std__pe27__lane0_strm1_data_mask     ( std__pe27__lane0_strm1_data_mask  ),      

               // PE 27, Lane 1                 
               .pe27__std__lane1_strm0_ready         ( pe27__std__lane1_strm0_ready      ),      
               .std__pe27__lane1_strm0_cntl          ( std__pe27__lane1_strm0_cntl       ),      
               .std__pe27__lane1_strm0_data          ( std__pe27__lane1_strm0_data       ),      
               .std__pe27__lane1_strm0_data_valid    ( std__pe27__lane1_strm0_data_valid ),      
               .std__pe27__lane1_strm0_data_mask     ( std__pe27__lane1_strm0_data_mask  ),      

               .pe27__std__lane1_strm1_ready         ( pe27__std__lane1_strm1_ready      ),      
               .std__pe27__lane1_strm1_cntl          ( std__pe27__lane1_strm1_cntl       ),      
               .std__pe27__lane1_strm1_data          ( std__pe27__lane1_strm1_data       ),      
               .std__pe27__lane1_strm1_data_valid    ( std__pe27__lane1_strm1_data_valid ),      
               .std__pe27__lane1_strm1_data_mask     ( std__pe27__lane1_strm1_data_mask  ),      

               // PE 27, Lane 2                 
               .pe27__std__lane2_strm0_ready         ( pe27__std__lane2_strm0_ready      ),      
               .std__pe27__lane2_strm0_cntl          ( std__pe27__lane2_strm0_cntl       ),      
               .std__pe27__lane2_strm0_data          ( std__pe27__lane2_strm0_data       ),      
               .std__pe27__lane2_strm0_data_valid    ( std__pe27__lane2_strm0_data_valid ),      
               .std__pe27__lane2_strm0_data_mask     ( std__pe27__lane2_strm0_data_mask  ),      

               .pe27__std__lane2_strm1_ready         ( pe27__std__lane2_strm1_ready      ),      
               .std__pe27__lane2_strm1_cntl          ( std__pe27__lane2_strm1_cntl       ),      
               .std__pe27__lane2_strm1_data          ( std__pe27__lane2_strm1_data       ),      
               .std__pe27__lane2_strm1_data_valid    ( std__pe27__lane2_strm1_data_valid ),      
               .std__pe27__lane2_strm1_data_mask     ( std__pe27__lane2_strm1_data_mask  ),      

               // PE 27, Lane 3                 
               .pe27__std__lane3_strm0_ready         ( pe27__std__lane3_strm0_ready      ),      
               .std__pe27__lane3_strm0_cntl          ( std__pe27__lane3_strm0_cntl       ),      
               .std__pe27__lane3_strm0_data          ( std__pe27__lane3_strm0_data       ),      
               .std__pe27__lane3_strm0_data_valid    ( std__pe27__lane3_strm0_data_valid ),      
               .std__pe27__lane3_strm0_data_mask     ( std__pe27__lane3_strm0_data_mask  ),      

               .pe27__std__lane3_strm1_ready         ( pe27__std__lane3_strm1_ready      ),      
               .std__pe27__lane3_strm1_cntl          ( std__pe27__lane3_strm1_cntl       ),      
               .std__pe27__lane3_strm1_data          ( std__pe27__lane3_strm1_data       ),      
               .std__pe27__lane3_strm1_data_valid    ( std__pe27__lane3_strm1_data_valid ),      
               .std__pe27__lane3_strm1_data_mask     ( std__pe27__lane3_strm1_data_mask  ),      

               // PE 27, Lane 4                 
               .pe27__std__lane4_strm0_ready         ( pe27__std__lane4_strm0_ready      ),      
               .std__pe27__lane4_strm0_cntl          ( std__pe27__lane4_strm0_cntl       ),      
               .std__pe27__lane4_strm0_data          ( std__pe27__lane4_strm0_data       ),      
               .std__pe27__lane4_strm0_data_valid    ( std__pe27__lane4_strm0_data_valid ),      
               .std__pe27__lane4_strm0_data_mask     ( std__pe27__lane4_strm0_data_mask  ),      

               .pe27__std__lane4_strm1_ready         ( pe27__std__lane4_strm1_ready      ),      
               .std__pe27__lane4_strm1_cntl          ( std__pe27__lane4_strm1_cntl       ),      
               .std__pe27__lane4_strm1_data          ( std__pe27__lane4_strm1_data       ),      
               .std__pe27__lane4_strm1_data_valid    ( std__pe27__lane4_strm1_data_valid ),      
               .std__pe27__lane4_strm1_data_mask     ( std__pe27__lane4_strm1_data_mask  ),      

               // PE 27, Lane 5                 
               .pe27__std__lane5_strm0_ready         ( pe27__std__lane5_strm0_ready      ),      
               .std__pe27__lane5_strm0_cntl          ( std__pe27__lane5_strm0_cntl       ),      
               .std__pe27__lane5_strm0_data          ( std__pe27__lane5_strm0_data       ),      
               .std__pe27__lane5_strm0_data_valid    ( std__pe27__lane5_strm0_data_valid ),      
               .std__pe27__lane5_strm0_data_mask     ( std__pe27__lane5_strm0_data_mask  ),      

               .pe27__std__lane5_strm1_ready         ( pe27__std__lane5_strm1_ready      ),      
               .std__pe27__lane5_strm1_cntl          ( std__pe27__lane5_strm1_cntl       ),      
               .std__pe27__lane5_strm1_data          ( std__pe27__lane5_strm1_data       ),      
               .std__pe27__lane5_strm1_data_valid    ( std__pe27__lane5_strm1_data_valid ),      
               .std__pe27__lane5_strm1_data_mask     ( std__pe27__lane5_strm1_data_mask  ),      

               // PE 27, Lane 6                 
               .pe27__std__lane6_strm0_ready         ( pe27__std__lane6_strm0_ready      ),      
               .std__pe27__lane6_strm0_cntl          ( std__pe27__lane6_strm0_cntl       ),      
               .std__pe27__lane6_strm0_data          ( std__pe27__lane6_strm0_data       ),      
               .std__pe27__lane6_strm0_data_valid    ( std__pe27__lane6_strm0_data_valid ),      
               .std__pe27__lane6_strm0_data_mask     ( std__pe27__lane6_strm0_data_mask  ),      

               .pe27__std__lane6_strm1_ready         ( pe27__std__lane6_strm1_ready      ),      
               .std__pe27__lane6_strm1_cntl          ( std__pe27__lane6_strm1_cntl       ),      
               .std__pe27__lane6_strm1_data          ( std__pe27__lane6_strm1_data       ),      
               .std__pe27__lane6_strm1_data_valid    ( std__pe27__lane6_strm1_data_valid ),      
               .std__pe27__lane6_strm1_data_mask     ( std__pe27__lane6_strm1_data_mask  ),      

               // PE 27, Lane 7                 
               .pe27__std__lane7_strm0_ready         ( pe27__std__lane7_strm0_ready      ),      
               .std__pe27__lane7_strm0_cntl          ( std__pe27__lane7_strm0_cntl       ),      
               .std__pe27__lane7_strm0_data          ( std__pe27__lane7_strm0_data       ),      
               .std__pe27__lane7_strm0_data_valid    ( std__pe27__lane7_strm0_data_valid ),      
               .std__pe27__lane7_strm0_data_mask     ( std__pe27__lane7_strm0_data_mask  ),      

               .pe27__std__lane7_strm1_ready         ( pe27__std__lane7_strm1_ready      ),      
               .std__pe27__lane7_strm1_cntl          ( std__pe27__lane7_strm1_cntl       ),      
               .std__pe27__lane7_strm1_data          ( std__pe27__lane7_strm1_data       ),      
               .std__pe27__lane7_strm1_data_valid    ( std__pe27__lane7_strm1_data_valid ),      
               .std__pe27__lane7_strm1_data_mask     ( std__pe27__lane7_strm1_data_mask  ),      

               // PE 27, Lane 8                 
               .pe27__std__lane8_strm0_ready         ( pe27__std__lane8_strm0_ready      ),      
               .std__pe27__lane8_strm0_cntl          ( std__pe27__lane8_strm0_cntl       ),      
               .std__pe27__lane8_strm0_data          ( std__pe27__lane8_strm0_data       ),      
               .std__pe27__lane8_strm0_data_valid    ( std__pe27__lane8_strm0_data_valid ),      
               .std__pe27__lane8_strm0_data_mask     ( std__pe27__lane8_strm0_data_mask  ),      

               .pe27__std__lane8_strm1_ready         ( pe27__std__lane8_strm1_ready      ),      
               .std__pe27__lane8_strm1_cntl          ( std__pe27__lane8_strm1_cntl       ),      
               .std__pe27__lane8_strm1_data          ( std__pe27__lane8_strm1_data       ),      
               .std__pe27__lane8_strm1_data_valid    ( std__pe27__lane8_strm1_data_valid ),      
               .std__pe27__lane8_strm1_data_mask     ( std__pe27__lane8_strm1_data_mask  ),      

               // PE 27, Lane 9                 
               .pe27__std__lane9_strm0_ready         ( pe27__std__lane9_strm0_ready      ),      
               .std__pe27__lane9_strm0_cntl          ( std__pe27__lane9_strm0_cntl       ),      
               .std__pe27__lane9_strm0_data          ( std__pe27__lane9_strm0_data       ),      
               .std__pe27__lane9_strm0_data_valid    ( std__pe27__lane9_strm0_data_valid ),      
               .std__pe27__lane9_strm0_data_mask     ( std__pe27__lane9_strm0_data_mask  ),      

               .pe27__std__lane9_strm1_ready         ( pe27__std__lane9_strm1_ready      ),      
               .std__pe27__lane9_strm1_cntl          ( std__pe27__lane9_strm1_cntl       ),      
               .std__pe27__lane9_strm1_data          ( std__pe27__lane9_strm1_data       ),      
               .std__pe27__lane9_strm1_data_valid    ( std__pe27__lane9_strm1_data_valid ),      
               .std__pe27__lane9_strm1_data_mask     ( std__pe27__lane9_strm1_data_mask  ),      

               // PE 27, Lane 10                 
               .pe27__std__lane10_strm0_ready         ( pe27__std__lane10_strm0_ready      ),      
               .std__pe27__lane10_strm0_cntl          ( std__pe27__lane10_strm0_cntl       ),      
               .std__pe27__lane10_strm0_data          ( std__pe27__lane10_strm0_data       ),      
               .std__pe27__lane10_strm0_data_valid    ( std__pe27__lane10_strm0_data_valid ),      
               .std__pe27__lane10_strm0_data_mask     ( std__pe27__lane10_strm0_data_mask  ),      

               .pe27__std__lane10_strm1_ready         ( pe27__std__lane10_strm1_ready      ),      
               .std__pe27__lane10_strm1_cntl          ( std__pe27__lane10_strm1_cntl       ),      
               .std__pe27__lane10_strm1_data          ( std__pe27__lane10_strm1_data       ),      
               .std__pe27__lane10_strm1_data_valid    ( std__pe27__lane10_strm1_data_valid ),      
               .std__pe27__lane10_strm1_data_mask     ( std__pe27__lane10_strm1_data_mask  ),      

               // PE 27, Lane 11                 
               .pe27__std__lane11_strm0_ready         ( pe27__std__lane11_strm0_ready      ),      
               .std__pe27__lane11_strm0_cntl          ( std__pe27__lane11_strm0_cntl       ),      
               .std__pe27__lane11_strm0_data          ( std__pe27__lane11_strm0_data       ),      
               .std__pe27__lane11_strm0_data_valid    ( std__pe27__lane11_strm0_data_valid ),      
               .std__pe27__lane11_strm0_data_mask     ( std__pe27__lane11_strm0_data_mask  ),      

               .pe27__std__lane11_strm1_ready         ( pe27__std__lane11_strm1_ready      ),      
               .std__pe27__lane11_strm1_cntl          ( std__pe27__lane11_strm1_cntl       ),      
               .std__pe27__lane11_strm1_data          ( std__pe27__lane11_strm1_data       ),      
               .std__pe27__lane11_strm1_data_valid    ( std__pe27__lane11_strm1_data_valid ),      
               .std__pe27__lane11_strm1_data_mask     ( std__pe27__lane11_strm1_data_mask  ),      

               // PE 27, Lane 12                 
               .pe27__std__lane12_strm0_ready         ( pe27__std__lane12_strm0_ready      ),      
               .std__pe27__lane12_strm0_cntl          ( std__pe27__lane12_strm0_cntl       ),      
               .std__pe27__lane12_strm0_data          ( std__pe27__lane12_strm0_data       ),      
               .std__pe27__lane12_strm0_data_valid    ( std__pe27__lane12_strm0_data_valid ),      
               .std__pe27__lane12_strm0_data_mask     ( std__pe27__lane12_strm0_data_mask  ),      

               .pe27__std__lane12_strm1_ready         ( pe27__std__lane12_strm1_ready      ),      
               .std__pe27__lane12_strm1_cntl          ( std__pe27__lane12_strm1_cntl       ),      
               .std__pe27__lane12_strm1_data          ( std__pe27__lane12_strm1_data       ),      
               .std__pe27__lane12_strm1_data_valid    ( std__pe27__lane12_strm1_data_valid ),      
               .std__pe27__lane12_strm1_data_mask     ( std__pe27__lane12_strm1_data_mask  ),      

               // PE 27, Lane 13                 
               .pe27__std__lane13_strm0_ready         ( pe27__std__lane13_strm0_ready      ),      
               .std__pe27__lane13_strm0_cntl          ( std__pe27__lane13_strm0_cntl       ),      
               .std__pe27__lane13_strm0_data          ( std__pe27__lane13_strm0_data       ),      
               .std__pe27__lane13_strm0_data_valid    ( std__pe27__lane13_strm0_data_valid ),      
               .std__pe27__lane13_strm0_data_mask     ( std__pe27__lane13_strm0_data_mask  ),      

               .pe27__std__lane13_strm1_ready         ( pe27__std__lane13_strm1_ready      ),      
               .std__pe27__lane13_strm1_cntl          ( std__pe27__lane13_strm1_cntl       ),      
               .std__pe27__lane13_strm1_data          ( std__pe27__lane13_strm1_data       ),      
               .std__pe27__lane13_strm1_data_valid    ( std__pe27__lane13_strm1_data_valid ),      
               .std__pe27__lane13_strm1_data_mask     ( std__pe27__lane13_strm1_data_mask  ),      

               // PE 27, Lane 14                 
               .pe27__std__lane14_strm0_ready         ( pe27__std__lane14_strm0_ready      ),      
               .std__pe27__lane14_strm0_cntl          ( std__pe27__lane14_strm0_cntl       ),      
               .std__pe27__lane14_strm0_data          ( std__pe27__lane14_strm0_data       ),      
               .std__pe27__lane14_strm0_data_valid    ( std__pe27__lane14_strm0_data_valid ),      
               .std__pe27__lane14_strm0_data_mask     ( std__pe27__lane14_strm0_data_mask  ),      

               .pe27__std__lane14_strm1_ready         ( pe27__std__lane14_strm1_ready      ),      
               .std__pe27__lane14_strm1_cntl          ( std__pe27__lane14_strm1_cntl       ),      
               .std__pe27__lane14_strm1_data          ( std__pe27__lane14_strm1_data       ),      
               .std__pe27__lane14_strm1_data_valid    ( std__pe27__lane14_strm1_data_valid ),      
               .std__pe27__lane14_strm1_data_mask     ( std__pe27__lane14_strm1_data_mask  ),      

               // PE 27, Lane 15                 
               .pe27__std__lane15_strm0_ready         ( pe27__std__lane15_strm0_ready      ),      
               .std__pe27__lane15_strm0_cntl          ( std__pe27__lane15_strm0_cntl       ),      
               .std__pe27__lane15_strm0_data          ( std__pe27__lane15_strm0_data       ),      
               .std__pe27__lane15_strm0_data_valid    ( std__pe27__lane15_strm0_data_valid ),      
               .std__pe27__lane15_strm0_data_mask     ( std__pe27__lane15_strm0_data_mask  ),      

               .pe27__std__lane15_strm1_ready         ( pe27__std__lane15_strm1_ready      ),      
               .std__pe27__lane15_strm1_cntl          ( std__pe27__lane15_strm1_cntl       ),      
               .std__pe27__lane15_strm1_data          ( std__pe27__lane15_strm1_data       ),      
               .std__pe27__lane15_strm1_data_valid    ( std__pe27__lane15_strm1_data_valid ),      
               .std__pe27__lane15_strm1_data_mask     ( std__pe27__lane15_strm1_data_mask  ),      

               // PE 27, Lane 16                 
               .pe27__std__lane16_strm0_ready         ( pe27__std__lane16_strm0_ready      ),      
               .std__pe27__lane16_strm0_cntl          ( std__pe27__lane16_strm0_cntl       ),      
               .std__pe27__lane16_strm0_data          ( std__pe27__lane16_strm0_data       ),      
               .std__pe27__lane16_strm0_data_valid    ( std__pe27__lane16_strm0_data_valid ),      
               .std__pe27__lane16_strm0_data_mask     ( std__pe27__lane16_strm0_data_mask  ),      

               .pe27__std__lane16_strm1_ready         ( pe27__std__lane16_strm1_ready      ),      
               .std__pe27__lane16_strm1_cntl          ( std__pe27__lane16_strm1_cntl       ),      
               .std__pe27__lane16_strm1_data          ( std__pe27__lane16_strm1_data       ),      
               .std__pe27__lane16_strm1_data_valid    ( std__pe27__lane16_strm1_data_valid ),      
               .std__pe27__lane16_strm1_data_mask     ( std__pe27__lane16_strm1_data_mask  ),      

               // PE 27, Lane 17                 
               .pe27__std__lane17_strm0_ready         ( pe27__std__lane17_strm0_ready      ),      
               .std__pe27__lane17_strm0_cntl          ( std__pe27__lane17_strm0_cntl       ),      
               .std__pe27__lane17_strm0_data          ( std__pe27__lane17_strm0_data       ),      
               .std__pe27__lane17_strm0_data_valid    ( std__pe27__lane17_strm0_data_valid ),      
               .std__pe27__lane17_strm0_data_mask     ( std__pe27__lane17_strm0_data_mask  ),      

               .pe27__std__lane17_strm1_ready         ( pe27__std__lane17_strm1_ready      ),      
               .std__pe27__lane17_strm1_cntl          ( std__pe27__lane17_strm1_cntl       ),      
               .std__pe27__lane17_strm1_data          ( std__pe27__lane17_strm1_data       ),      
               .std__pe27__lane17_strm1_data_valid    ( std__pe27__lane17_strm1_data_valid ),      
               .std__pe27__lane17_strm1_data_mask     ( std__pe27__lane17_strm1_data_mask  ),      

               // PE 27, Lane 18                 
               .pe27__std__lane18_strm0_ready         ( pe27__std__lane18_strm0_ready      ),      
               .std__pe27__lane18_strm0_cntl          ( std__pe27__lane18_strm0_cntl       ),      
               .std__pe27__lane18_strm0_data          ( std__pe27__lane18_strm0_data       ),      
               .std__pe27__lane18_strm0_data_valid    ( std__pe27__lane18_strm0_data_valid ),      
               .std__pe27__lane18_strm0_data_mask     ( std__pe27__lane18_strm0_data_mask  ),      

               .pe27__std__lane18_strm1_ready         ( pe27__std__lane18_strm1_ready      ),      
               .std__pe27__lane18_strm1_cntl          ( std__pe27__lane18_strm1_cntl       ),      
               .std__pe27__lane18_strm1_data          ( std__pe27__lane18_strm1_data       ),      
               .std__pe27__lane18_strm1_data_valid    ( std__pe27__lane18_strm1_data_valid ),      
               .std__pe27__lane18_strm1_data_mask     ( std__pe27__lane18_strm1_data_mask  ),      

               // PE 27, Lane 19                 
               .pe27__std__lane19_strm0_ready         ( pe27__std__lane19_strm0_ready      ),      
               .std__pe27__lane19_strm0_cntl          ( std__pe27__lane19_strm0_cntl       ),      
               .std__pe27__lane19_strm0_data          ( std__pe27__lane19_strm0_data       ),      
               .std__pe27__lane19_strm0_data_valid    ( std__pe27__lane19_strm0_data_valid ),      
               .std__pe27__lane19_strm0_data_mask     ( std__pe27__lane19_strm0_data_mask  ),      

               .pe27__std__lane19_strm1_ready         ( pe27__std__lane19_strm1_ready      ),      
               .std__pe27__lane19_strm1_cntl          ( std__pe27__lane19_strm1_cntl       ),      
               .std__pe27__lane19_strm1_data          ( std__pe27__lane19_strm1_data       ),      
               .std__pe27__lane19_strm1_data_valid    ( std__pe27__lane19_strm1_data_valid ),      
               .std__pe27__lane19_strm1_data_mask     ( std__pe27__lane19_strm1_data_mask  ),      

               // PE 27, Lane 20                 
               .pe27__std__lane20_strm0_ready         ( pe27__std__lane20_strm0_ready      ),      
               .std__pe27__lane20_strm0_cntl          ( std__pe27__lane20_strm0_cntl       ),      
               .std__pe27__lane20_strm0_data          ( std__pe27__lane20_strm0_data       ),      
               .std__pe27__lane20_strm0_data_valid    ( std__pe27__lane20_strm0_data_valid ),      
               .std__pe27__lane20_strm0_data_mask     ( std__pe27__lane20_strm0_data_mask  ),      

               .pe27__std__lane20_strm1_ready         ( pe27__std__lane20_strm1_ready      ),      
               .std__pe27__lane20_strm1_cntl          ( std__pe27__lane20_strm1_cntl       ),      
               .std__pe27__lane20_strm1_data          ( std__pe27__lane20_strm1_data       ),      
               .std__pe27__lane20_strm1_data_valid    ( std__pe27__lane20_strm1_data_valid ),      
               .std__pe27__lane20_strm1_data_mask     ( std__pe27__lane20_strm1_data_mask  ),      

               // PE 27, Lane 21                 
               .pe27__std__lane21_strm0_ready         ( pe27__std__lane21_strm0_ready      ),      
               .std__pe27__lane21_strm0_cntl          ( std__pe27__lane21_strm0_cntl       ),      
               .std__pe27__lane21_strm0_data          ( std__pe27__lane21_strm0_data       ),      
               .std__pe27__lane21_strm0_data_valid    ( std__pe27__lane21_strm0_data_valid ),      
               .std__pe27__lane21_strm0_data_mask     ( std__pe27__lane21_strm0_data_mask  ),      

               .pe27__std__lane21_strm1_ready         ( pe27__std__lane21_strm1_ready      ),      
               .std__pe27__lane21_strm1_cntl          ( std__pe27__lane21_strm1_cntl       ),      
               .std__pe27__lane21_strm1_data          ( std__pe27__lane21_strm1_data       ),      
               .std__pe27__lane21_strm1_data_valid    ( std__pe27__lane21_strm1_data_valid ),      
               .std__pe27__lane21_strm1_data_mask     ( std__pe27__lane21_strm1_data_mask  ),      

               // PE 27, Lane 22                 
               .pe27__std__lane22_strm0_ready         ( pe27__std__lane22_strm0_ready      ),      
               .std__pe27__lane22_strm0_cntl          ( std__pe27__lane22_strm0_cntl       ),      
               .std__pe27__lane22_strm0_data          ( std__pe27__lane22_strm0_data       ),      
               .std__pe27__lane22_strm0_data_valid    ( std__pe27__lane22_strm0_data_valid ),      
               .std__pe27__lane22_strm0_data_mask     ( std__pe27__lane22_strm0_data_mask  ),      

               .pe27__std__lane22_strm1_ready         ( pe27__std__lane22_strm1_ready      ),      
               .std__pe27__lane22_strm1_cntl          ( std__pe27__lane22_strm1_cntl       ),      
               .std__pe27__lane22_strm1_data          ( std__pe27__lane22_strm1_data       ),      
               .std__pe27__lane22_strm1_data_valid    ( std__pe27__lane22_strm1_data_valid ),      
               .std__pe27__lane22_strm1_data_mask     ( std__pe27__lane22_strm1_data_mask  ),      

               // PE 27, Lane 23                 
               .pe27__std__lane23_strm0_ready         ( pe27__std__lane23_strm0_ready      ),      
               .std__pe27__lane23_strm0_cntl          ( std__pe27__lane23_strm0_cntl       ),      
               .std__pe27__lane23_strm0_data          ( std__pe27__lane23_strm0_data       ),      
               .std__pe27__lane23_strm0_data_valid    ( std__pe27__lane23_strm0_data_valid ),      
               .std__pe27__lane23_strm0_data_mask     ( std__pe27__lane23_strm0_data_mask  ),      

               .pe27__std__lane23_strm1_ready         ( pe27__std__lane23_strm1_ready      ),      
               .std__pe27__lane23_strm1_cntl          ( std__pe27__lane23_strm1_cntl       ),      
               .std__pe27__lane23_strm1_data          ( std__pe27__lane23_strm1_data       ),      
               .std__pe27__lane23_strm1_data_valid    ( std__pe27__lane23_strm1_data_valid ),      
               .std__pe27__lane23_strm1_data_mask     ( std__pe27__lane23_strm1_data_mask  ),      

               // PE 27, Lane 24                 
               .pe27__std__lane24_strm0_ready         ( pe27__std__lane24_strm0_ready      ),      
               .std__pe27__lane24_strm0_cntl          ( std__pe27__lane24_strm0_cntl       ),      
               .std__pe27__lane24_strm0_data          ( std__pe27__lane24_strm0_data       ),      
               .std__pe27__lane24_strm0_data_valid    ( std__pe27__lane24_strm0_data_valid ),      
               .std__pe27__lane24_strm0_data_mask     ( std__pe27__lane24_strm0_data_mask  ),      

               .pe27__std__lane24_strm1_ready         ( pe27__std__lane24_strm1_ready      ),      
               .std__pe27__lane24_strm1_cntl          ( std__pe27__lane24_strm1_cntl       ),      
               .std__pe27__lane24_strm1_data          ( std__pe27__lane24_strm1_data       ),      
               .std__pe27__lane24_strm1_data_valid    ( std__pe27__lane24_strm1_data_valid ),      
               .std__pe27__lane24_strm1_data_mask     ( std__pe27__lane24_strm1_data_mask  ),      

               // PE 27, Lane 25                 
               .pe27__std__lane25_strm0_ready         ( pe27__std__lane25_strm0_ready      ),      
               .std__pe27__lane25_strm0_cntl          ( std__pe27__lane25_strm0_cntl       ),      
               .std__pe27__lane25_strm0_data          ( std__pe27__lane25_strm0_data       ),      
               .std__pe27__lane25_strm0_data_valid    ( std__pe27__lane25_strm0_data_valid ),      
               .std__pe27__lane25_strm0_data_mask     ( std__pe27__lane25_strm0_data_mask  ),      

               .pe27__std__lane25_strm1_ready         ( pe27__std__lane25_strm1_ready      ),      
               .std__pe27__lane25_strm1_cntl          ( std__pe27__lane25_strm1_cntl       ),      
               .std__pe27__lane25_strm1_data          ( std__pe27__lane25_strm1_data       ),      
               .std__pe27__lane25_strm1_data_valid    ( std__pe27__lane25_strm1_data_valid ),      
               .std__pe27__lane25_strm1_data_mask     ( std__pe27__lane25_strm1_data_mask  ),      

               // PE 27, Lane 26                 
               .pe27__std__lane26_strm0_ready         ( pe27__std__lane26_strm0_ready      ),      
               .std__pe27__lane26_strm0_cntl          ( std__pe27__lane26_strm0_cntl       ),      
               .std__pe27__lane26_strm0_data          ( std__pe27__lane26_strm0_data       ),      
               .std__pe27__lane26_strm0_data_valid    ( std__pe27__lane26_strm0_data_valid ),      
               .std__pe27__lane26_strm0_data_mask     ( std__pe27__lane26_strm0_data_mask  ),      

               .pe27__std__lane26_strm1_ready         ( pe27__std__lane26_strm1_ready      ),      
               .std__pe27__lane26_strm1_cntl          ( std__pe27__lane26_strm1_cntl       ),      
               .std__pe27__lane26_strm1_data          ( std__pe27__lane26_strm1_data       ),      
               .std__pe27__lane26_strm1_data_valid    ( std__pe27__lane26_strm1_data_valid ),      
               .std__pe27__lane26_strm1_data_mask     ( std__pe27__lane26_strm1_data_mask  ),      

               // PE 27, Lane 27                 
               .pe27__std__lane27_strm0_ready         ( pe27__std__lane27_strm0_ready      ),      
               .std__pe27__lane27_strm0_cntl          ( std__pe27__lane27_strm0_cntl       ),      
               .std__pe27__lane27_strm0_data          ( std__pe27__lane27_strm0_data       ),      
               .std__pe27__lane27_strm0_data_valid    ( std__pe27__lane27_strm0_data_valid ),      
               .std__pe27__lane27_strm0_data_mask     ( std__pe27__lane27_strm0_data_mask  ),      

               .pe27__std__lane27_strm1_ready         ( pe27__std__lane27_strm1_ready      ),      
               .std__pe27__lane27_strm1_cntl          ( std__pe27__lane27_strm1_cntl       ),      
               .std__pe27__lane27_strm1_data          ( std__pe27__lane27_strm1_data       ),      
               .std__pe27__lane27_strm1_data_valid    ( std__pe27__lane27_strm1_data_valid ),      
               .std__pe27__lane27_strm1_data_mask     ( std__pe27__lane27_strm1_data_mask  ),      

               // PE 27, Lane 28                 
               .pe27__std__lane28_strm0_ready         ( pe27__std__lane28_strm0_ready      ),      
               .std__pe27__lane28_strm0_cntl          ( std__pe27__lane28_strm0_cntl       ),      
               .std__pe27__lane28_strm0_data          ( std__pe27__lane28_strm0_data       ),      
               .std__pe27__lane28_strm0_data_valid    ( std__pe27__lane28_strm0_data_valid ),      
               .std__pe27__lane28_strm0_data_mask     ( std__pe27__lane28_strm0_data_mask  ),      

               .pe27__std__lane28_strm1_ready         ( pe27__std__lane28_strm1_ready      ),      
               .std__pe27__lane28_strm1_cntl          ( std__pe27__lane28_strm1_cntl       ),      
               .std__pe27__lane28_strm1_data          ( std__pe27__lane28_strm1_data       ),      
               .std__pe27__lane28_strm1_data_valid    ( std__pe27__lane28_strm1_data_valid ),      
               .std__pe27__lane28_strm1_data_mask     ( std__pe27__lane28_strm1_data_mask  ),      

               // PE 27, Lane 29                 
               .pe27__std__lane29_strm0_ready         ( pe27__std__lane29_strm0_ready      ),      
               .std__pe27__lane29_strm0_cntl          ( std__pe27__lane29_strm0_cntl       ),      
               .std__pe27__lane29_strm0_data          ( std__pe27__lane29_strm0_data       ),      
               .std__pe27__lane29_strm0_data_valid    ( std__pe27__lane29_strm0_data_valid ),      
               .std__pe27__lane29_strm0_data_mask     ( std__pe27__lane29_strm0_data_mask  ),      

               .pe27__std__lane29_strm1_ready         ( pe27__std__lane29_strm1_ready      ),      
               .std__pe27__lane29_strm1_cntl          ( std__pe27__lane29_strm1_cntl       ),      
               .std__pe27__lane29_strm1_data          ( std__pe27__lane29_strm1_data       ),      
               .std__pe27__lane29_strm1_data_valid    ( std__pe27__lane29_strm1_data_valid ),      
               .std__pe27__lane29_strm1_data_mask     ( std__pe27__lane29_strm1_data_mask  ),      

               // PE 27, Lane 30                 
               .pe27__std__lane30_strm0_ready         ( pe27__std__lane30_strm0_ready      ),      
               .std__pe27__lane30_strm0_cntl          ( std__pe27__lane30_strm0_cntl       ),      
               .std__pe27__lane30_strm0_data          ( std__pe27__lane30_strm0_data       ),      
               .std__pe27__lane30_strm0_data_valid    ( std__pe27__lane30_strm0_data_valid ),      
               .std__pe27__lane30_strm0_data_mask     ( std__pe27__lane30_strm0_data_mask  ),      

               .pe27__std__lane30_strm1_ready         ( pe27__std__lane30_strm1_ready      ),      
               .std__pe27__lane30_strm1_cntl          ( std__pe27__lane30_strm1_cntl       ),      
               .std__pe27__lane30_strm1_data          ( std__pe27__lane30_strm1_data       ),      
               .std__pe27__lane30_strm1_data_valid    ( std__pe27__lane30_strm1_data_valid ),      
               .std__pe27__lane30_strm1_data_mask     ( std__pe27__lane30_strm1_data_mask  ),      

               // PE 27, Lane 31                 
               .pe27__std__lane31_strm0_ready         ( pe27__std__lane31_strm0_ready      ),      
               .std__pe27__lane31_strm0_cntl          ( std__pe27__lane31_strm0_cntl       ),      
               .std__pe27__lane31_strm0_data          ( std__pe27__lane31_strm0_data       ),      
               .std__pe27__lane31_strm0_data_valid    ( std__pe27__lane31_strm0_data_valid ),      
               .std__pe27__lane31_strm0_data_mask     ( std__pe27__lane31_strm0_data_mask  ),      

               .pe27__std__lane31_strm1_ready         ( pe27__std__lane31_strm1_ready      ),      
               .std__pe27__lane31_strm1_cntl          ( std__pe27__lane31_strm1_cntl       ),      
               .std__pe27__lane31_strm1_data          ( std__pe27__lane31_strm1_data       ),      
               .std__pe27__lane31_strm1_data_valid    ( std__pe27__lane31_strm1_data_valid ),      
               .std__pe27__lane31_strm1_data_mask     ( std__pe27__lane31_strm1_data_mask  ),      

               // PE 28, Lane 0                 
               .pe28__std__lane0_strm0_ready         ( pe28__std__lane0_strm0_ready      ),      
               .std__pe28__lane0_strm0_cntl          ( std__pe28__lane0_strm0_cntl       ),      
               .std__pe28__lane0_strm0_data          ( std__pe28__lane0_strm0_data       ),      
               .std__pe28__lane0_strm0_data_valid    ( std__pe28__lane0_strm0_data_valid ),      
               .std__pe28__lane0_strm0_data_mask     ( std__pe28__lane0_strm0_data_mask  ),      

               .pe28__std__lane0_strm1_ready         ( pe28__std__lane0_strm1_ready      ),      
               .std__pe28__lane0_strm1_cntl          ( std__pe28__lane0_strm1_cntl       ),      
               .std__pe28__lane0_strm1_data          ( std__pe28__lane0_strm1_data       ),      
               .std__pe28__lane0_strm1_data_valid    ( std__pe28__lane0_strm1_data_valid ),      
               .std__pe28__lane0_strm1_data_mask     ( std__pe28__lane0_strm1_data_mask  ),      

               // PE 28, Lane 1                 
               .pe28__std__lane1_strm0_ready         ( pe28__std__lane1_strm0_ready      ),      
               .std__pe28__lane1_strm0_cntl          ( std__pe28__lane1_strm0_cntl       ),      
               .std__pe28__lane1_strm0_data          ( std__pe28__lane1_strm0_data       ),      
               .std__pe28__lane1_strm0_data_valid    ( std__pe28__lane1_strm0_data_valid ),      
               .std__pe28__lane1_strm0_data_mask     ( std__pe28__lane1_strm0_data_mask  ),      

               .pe28__std__lane1_strm1_ready         ( pe28__std__lane1_strm1_ready      ),      
               .std__pe28__lane1_strm1_cntl          ( std__pe28__lane1_strm1_cntl       ),      
               .std__pe28__lane1_strm1_data          ( std__pe28__lane1_strm1_data       ),      
               .std__pe28__lane1_strm1_data_valid    ( std__pe28__lane1_strm1_data_valid ),      
               .std__pe28__lane1_strm1_data_mask     ( std__pe28__lane1_strm1_data_mask  ),      

               // PE 28, Lane 2                 
               .pe28__std__lane2_strm0_ready         ( pe28__std__lane2_strm0_ready      ),      
               .std__pe28__lane2_strm0_cntl          ( std__pe28__lane2_strm0_cntl       ),      
               .std__pe28__lane2_strm0_data          ( std__pe28__lane2_strm0_data       ),      
               .std__pe28__lane2_strm0_data_valid    ( std__pe28__lane2_strm0_data_valid ),      
               .std__pe28__lane2_strm0_data_mask     ( std__pe28__lane2_strm0_data_mask  ),      

               .pe28__std__lane2_strm1_ready         ( pe28__std__lane2_strm1_ready      ),      
               .std__pe28__lane2_strm1_cntl          ( std__pe28__lane2_strm1_cntl       ),      
               .std__pe28__lane2_strm1_data          ( std__pe28__lane2_strm1_data       ),      
               .std__pe28__lane2_strm1_data_valid    ( std__pe28__lane2_strm1_data_valid ),      
               .std__pe28__lane2_strm1_data_mask     ( std__pe28__lane2_strm1_data_mask  ),      

               // PE 28, Lane 3                 
               .pe28__std__lane3_strm0_ready         ( pe28__std__lane3_strm0_ready      ),      
               .std__pe28__lane3_strm0_cntl          ( std__pe28__lane3_strm0_cntl       ),      
               .std__pe28__lane3_strm0_data          ( std__pe28__lane3_strm0_data       ),      
               .std__pe28__lane3_strm0_data_valid    ( std__pe28__lane3_strm0_data_valid ),      
               .std__pe28__lane3_strm0_data_mask     ( std__pe28__lane3_strm0_data_mask  ),      

               .pe28__std__lane3_strm1_ready         ( pe28__std__lane3_strm1_ready      ),      
               .std__pe28__lane3_strm1_cntl          ( std__pe28__lane3_strm1_cntl       ),      
               .std__pe28__lane3_strm1_data          ( std__pe28__lane3_strm1_data       ),      
               .std__pe28__lane3_strm1_data_valid    ( std__pe28__lane3_strm1_data_valid ),      
               .std__pe28__lane3_strm1_data_mask     ( std__pe28__lane3_strm1_data_mask  ),      

               // PE 28, Lane 4                 
               .pe28__std__lane4_strm0_ready         ( pe28__std__lane4_strm0_ready      ),      
               .std__pe28__lane4_strm0_cntl          ( std__pe28__lane4_strm0_cntl       ),      
               .std__pe28__lane4_strm0_data          ( std__pe28__lane4_strm0_data       ),      
               .std__pe28__lane4_strm0_data_valid    ( std__pe28__lane4_strm0_data_valid ),      
               .std__pe28__lane4_strm0_data_mask     ( std__pe28__lane4_strm0_data_mask  ),      

               .pe28__std__lane4_strm1_ready         ( pe28__std__lane4_strm1_ready      ),      
               .std__pe28__lane4_strm1_cntl          ( std__pe28__lane4_strm1_cntl       ),      
               .std__pe28__lane4_strm1_data          ( std__pe28__lane4_strm1_data       ),      
               .std__pe28__lane4_strm1_data_valid    ( std__pe28__lane4_strm1_data_valid ),      
               .std__pe28__lane4_strm1_data_mask     ( std__pe28__lane4_strm1_data_mask  ),      

               // PE 28, Lane 5                 
               .pe28__std__lane5_strm0_ready         ( pe28__std__lane5_strm0_ready      ),      
               .std__pe28__lane5_strm0_cntl          ( std__pe28__lane5_strm0_cntl       ),      
               .std__pe28__lane5_strm0_data          ( std__pe28__lane5_strm0_data       ),      
               .std__pe28__lane5_strm0_data_valid    ( std__pe28__lane5_strm0_data_valid ),      
               .std__pe28__lane5_strm0_data_mask     ( std__pe28__lane5_strm0_data_mask  ),      

               .pe28__std__lane5_strm1_ready         ( pe28__std__lane5_strm1_ready      ),      
               .std__pe28__lane5_strm1_cntl          ( std__pe28__lane5_strm1_cntl       ),      
               .std__pe28__lane5_strm1_data          ( std__pe28__lane5_strm1_data       ),      
               .std__pe28__lane5_strm1_data_valid    ( std__pe28__lane5_strm1_data_valid ),      
               .std__pe28__lane5_strm1_data_mask     ( std__pe28__lane5_strm1_data_mask  ),      

               // PE 28, Lane 6                 
               .pe28__std__lane6_strm0_ready         ( pe28__std__lane6_strm0_ready      ),      
               .std__pe28__lane6_strm0_cntl          ( std__pe28__lane6_strm0_cntl       ),      
               .std__pe28__lane6_strm0_data          ( std__pe28__lane6_strm0_data       ),      
               .std__pe28__lane6_strm0_data_valid    ( std__pe28__lane6_strm0_data_valid ),      
               .std__pe28__lane6_strm0_data_mask     ( std__pe28__lane6_strm0_data_mask  ),      

               .pe28__std__lane6_strm1_ready         ( pe28__std__lane6_strm1_ready      ),      
               .std__pe28__lane6_strm1_cntl          ( std__pe28__lane6_strm1_cntl       ),      
               .std__pe28__lane6_strm1_data          ( std__pe28__lane6_strm1_data       ),      
               .std__pe28__lane6_strm1_data_valid    ( std__pe28__lane6_strm1_data_valid ),      
               .std__pe28__lane6_strm1_data_mask     ( std__pe28__lane6_strm1_data_mask  ),      

               // PE 28, Lane 7                 
               .pe28__std__lane7_strm0_ready         ( pe28__std__lane7_strm0_ready      ),      
               .std__pe28__lane7_strm0_cntl          ( std__pe28__lane7_strm0_cntl       ),      
               .std__pe28__lane7_strm0_data          ( std__pe28__lane7_strm0_data       ),      
               .std__pe28__lane7_strm0_data_valid    ( std__pe28__lane7_strm0_data_valid ),      
               .std__pe28__lane7_strm0_data_mask     ( std__pe28__lane7_strm0_data_mask  ),      

               .pe28__std__lane7_strm1_ready         ( pe28__std__lane7_strm1_ready      ),      
               .std__pe28__lane7_strm1_cntl          ( std__pe28__lane7_strm1_cntl       ),      
               .std__pe28__lane7_strm1_data          ( std__pe28__lane7_strm1_data       ),      
               .std__pe28__lane7_strm1_data_valid    ( std__pe28__lane7_strm1_data_valid ),      
               .std__pe28__lane7_strm1_data_mask     ( std__pe28__lane7_strm1_data_mask  ),      

               // PE 28, Lane 8                 
               .pe28__std__lane8_strm0_ready         ( pe28__std__lane8_strm0_ready      ),      
               .std__pe28__lane8_strm0_cntl          ( std__pe28__lane8_strm0_cntl       ),      
               .std__pe28__lane8_strm0_data          ( std__pe28__lane8_strm0_data       ),      
               .std__pe28__lane8_strm0_data_valid    ( std__pe28__lane8_strm0_data_valid ),      
               .std__pe28__lane8_strm0_data_mask     ( std__pe28__lane8_strm0_data_mask  ),      

               .pe28__std__lane8_strm1_ready         ( pe28__std__lane8_strm1_ready      ),      
               .std__pe28__lane8_strm1_cntl          ( std__pe28__lane8_strm1_cntl       ),      
               .std__pe28__lane8_strm1_data          ( std__pe28__lane8_strm1_data       ),      
               .std__pe28__lane8_strm1_data_valid    ( std__pe28__lane8_strm1_data_valid ),      
               .std__pe28__lane8_strm1_data_mask     ( std__pe28__lane8_strm1_data_mask  ),      

               // PE 28, Lane 9                 
               .pe28__std__lane9_strm0_ready         ( pe28__std__lane9_strm0_ready      ),      
               .std__pe28__lane9_strm0_cntl          ( std__pe28__lane9_strm0_cntl       ),      
               .std__pe28__lane9_strm0_data          ( std__pe28__lane9_strm0_data       ),      
               .std__pe28__lane9_strm0_data_valid    ( std__pe28__lane9_strm0_data_valid ),      
               .std__pe28__lane9_strm0_data_mask     ( std__pe28__lane9_strm0_data_mask  ),      

               .pe28__std__lane9_strm1_ready         ( pe28__std__lane9_strm1_ready      ),      
               .std__pe28__lane9_strm1_cntl          ( std__pe28__lane9_strm1_cntl       ),      
               .std__pe28__lane9_strm1_data          ( std__pe28__lane9_strm1_data       ),      
               .std__pe28__lane9_strm1_data_valid    ( std__pe28__lane9_strm1_data_valid ),      
               .std__pe28__lane9_strm1_data_mask     ( std__pe28__lane9_strm1_data_mask  ),      

               // PE 28, Lane 10                 
               .pe28__std__lane10_strm0_ready         ( pe28__std__lane10_strm0_ready      ),      
               .std__pe28__lane10_strm0_cntl          ( std__pe28__lane10_strm0_cntl       ),      
               .std__pe28__lane10_strm0_data          ( std__pe28__lane10_strm0_data       ),      
               .std__pe28__lane10_strm0_data_valid    ( std__pe28__lane10_strm0_data_valid ),      
               .std__pe28__lane10_strm0_data_mask     ( std__pe28__lane10_strm0_data_mask  ),      

               .pe28__std__lane10_strm1_ready         ( pe28__std__lane10_strm1_ready      ),      
               .std__pe28__lane10_strm1_cntl          ( std__pe28__lane10_strm1_cntl       ),      
               .std__pe28__lane10_strm1_data          ( std__pe28__lane10_strm1_data       ),      
               .std__pe28__lane10_strm1_data_valid    ( std__pe28__lane10_strm1_data_valid ),      
               .std__pe28__lane10_strm1_data_mask     ( std__pe28__lane10_strm1_data_mask  ),      

               // PE 28, Lane 11                 
               .pe28__std__lane11_strm0_ready         ( pe28__std__lane11_strm0_ready      ),      
               .std__pe28__lane11_strm0_cntl          ( std__pe28__lane11_strm0_cntl       ),      
               .std__pe28__lane11_strm0_data          ( std__pe28__lane11_strm0_data       ),      
               .std__pe28__lane11_strm0_data_valid    ( std__pe28__lane11_strm0_data_valid ),      
               .std__pe28__lane11_strm0_data_mask     ( std__pe28__lane11_strm0_data_mask  ),      

               .pe28__std__lane11_strm1_ready         ( pe28__std__lane11_strm1_ready      ),      
               .std__pe28__lane11_strm1_cntl          ( std__pe28__lane11_strm1_cntl       ),      
               .std__pe28__lane11_strm1_data          ( std__pe28__lane11_strm1_data       ),      
               .std__pe28__lane11_strm1_data_valid    ( std__pe28__lane11_strm1_data_valid ),      
               .std__pe28__lane11_strm1_data_mask     ( std__pe28__lane11_strm1_data_mask  ),      

               // PE 28, Lane 12                 
               .pe28__std__lane12_strm0_ready         ( pe28__std__lane12_strm0_ready      ),      
               .std__pe28__lane12_strm0_cntl          ( std__pe28__lane12_strm0_cntl       ),      
               .std__pe28__lane12_strm0_data          ( std__pe28__lane12_strm0_data       ),      
               .std__pe28__lane12_strm0_data_valid    ( std__pe28__lane12_strm0_data_valid ),      
               .std__pe28__lane12_strm0_data_mask     ( std__pe28__lane12_strm0_data_mask  ),      

               .pe28__std__lane12_strm1_ready         ( pe28__std__lane12_strm1_ready      ),      
               .std__pe28__lane12_strm1_cntl          ( std__pe28__lane12_strm1_cntl       ),      
               .std__pe28__lane12_strm1_data          ( std__pe28__lane12_strm1_data       ),      
               .std__pe28__lane12_strm1_data_valid    ( std__pe28__lane12_strm1_data_valid ),      
               .std__pe28__lane12_strm1_data_mask     ( std__pe28__lane12_strm1_data_mask  ),      

               // PE 28, Lane 13                 
               .pe28__std__lane13_strm0_ready         ( pe28__std__lane13_strm0_ready      ),      
               .std__pe28__lane13_strm0_cntl          ( std__pe28__lane13_strm0_cntl       ),      
               .std__pe28__lane13_strm0_data          ( std__pe28__lane13_strm0_data       ),      
               .std__pe28__lane13_strm0_data_valid    ( std__pe28__lane13_strm0_data_valid ),      
               .std__pe28__lane13_strm0_data_mask     ( std__pe28__lane13_strm0_data_mask  ),      

               .pe28__std__lane13_strm1_ready         ( pe28__std__lane13_strm1_ready      ),      
               .std__pe28__lane13_strm1_cntl          ( std__pe28__lane13_strm1_cntl       ),      
               .std__pe28__lane13_strm1_data          ( std__pe28__lane13_strm1_data       ),      
               .std__pe28__lane13_strm1_data_valid    ( std__pe28__lane13_strm1_data_valid ),      
               .std__pe28__lane13_strm1_data_mask     ( std__pe28__lane13_strm1_data_mask  ),      

               // PE 28, Lane 14                 
               .pe28__std__lane14_strm0_ready         ( pe28__std__lane14_strm0_ready      ),      
               .std__pe28__lane14_strm0_cntl          ( std__pe28__lane14_strm0_cntl       ),      
               .std__pe28__lane14_strm0_data          ( std__pe28__lane14_strm0_data       ),      
               .std__pe28__lane14_strm0_data_valid    ( std__pe28__lane14_strm0_data_valid ),      
               .std__pe28__lane14_strm0_data_mask     ( std__pe28__lane14_strm0_data_mask  ),      

               .pe28__std__lane14_strm1_ready         ( pe28__std__lane14_strm1_ready      ),      
               .std__pe28__lane14_strm1_cntl          ( std__pe28__lane14_strm1_cntl       ),      
               .std__pe28__lane14_strm1_data          ( std__pe28__lane14_strm1_data       ),      
               .std__pe28__lane14_strm1_data_valid    ( std__pe28__lane14_strm1_data_valid ),      
               .std__pe28__lane14_strm1_data_mask     ( std__pe28__lane14_strm1_data_mask  ),      

               // PE 28, Lane 15                 
               .pe28__std__lane15_strm0_ready         ( pe28__std__lane15_strm0_ready      ),      
               .std__pe28__lane15_strm0_cntl          ( std__pe28__lane15_strm0_cntl       ),      
               .std__pe28__lane15_strm0_data          ( std__pe28__lane15_strm0_data       ),      
               .std__pe28__lane15_strm0_data_valid    ( std__pe28__lane15_strm0_data_valid ),      
               .std__pe28__lane15_strm0_data_mask     ( std__pe28__lane15_strm0_data_mask  ),      

               .pe28__std__lane15_strm1_ready         ( pe28__std__lane15_strm1_ready      ),      
               .std__pe28__lane15_strm1_cntl          ( std__pe28__lane15_strm1_cntl       ),      
               .std__pe28__lane15_strm1_data          ( std__pe28__lane15_strm1_data       ),      
               .std__pe28__lane15_strm1_data_valid    ( std__pe28__lane15_strm1_data_valid ),      
               .std__pe28__lane15_strm1_data_mask     ( std__pe28__lane15_strm1_data_mask  ),      

               // PE 28, Lane 16                 
               .pe28__std__lane16_strm0_ready         ( pe28__std__lane16_strm0_ready      ),      
               .std__pe28__lane16_strm0_cntl          ( std__pe28__lane16_strm0_cntl       ),      
               .std__pe28__lane16_strm0_data          ( std__pe28__lane16_strm0_data       ),      
               .std__pe28__lane16_strm0_data_valid    ( std__pe28__lane16_strm0_data_valid ),      
               .std__pe28__lane16_strm0_data_mask     ( std__pe28__lane16_strm0_data_mask  ),      

               .pe28__std__lane16_strm1_ready         ( pe28__std__lane16_strm1_ready      ),      
               .std__pe28__lane16_strm1_cntl          ( std__pe28__lane16_strm1_cntl       ),      
               .std__pe28__lane16_strm1_data          ( std__pe28__lane16_strm1_data       ),      
               .std__pe28__lane16_strm1_data_valid    ( std__pe28__lane16_strm1_data_valid ),      
               .std__pe28__lane16_strm1_data_mask     ( std__pe28__lane16_strm1_data_mask  ),      

               // PE 28, Lane 17                 
               .pe28__std__lane17_strm0_ready         ( pe28__std__lane17_strm0_ready      ),      
               .std__pe28__lane17_strm0_cntl          ( std__pe28__lane17_strm0_cntl       ),      
               .std__pe28__lane17_strm0_data          ( std__pe28__lane17_strm0_data       ),      
               .std__pe28__lane17_strm0_data_valid    ( std__pe28__lane17_strm0_data_valid ),      
               .std__pe28__lane17_strm0_data_mask     ( std__pe28__lane17_strm0_data_mask  ),      

               .pe28__std__lane17_strm1_ready         ( pe28__std__lane17_strm1_ready      ),      
               .std__pe28__lane17_strm1_cntl          ( std__pe28__lane17_strm1_cntl       ),      
               .std__pe28__lane17_strm1_data          ( std__pe28__lane17_strm1_data       ),      
               .std__pe28__lane17_strm1_data_valid    ( std__pe28__lane17_strm1_data_valid ),      
               .std__pe28__lane17_strm1_data_mask     ( std__pe28__lane17_strm1_data_mask  ),      

               // PE 28, Lane 18                 
               .pe28__std__lane18_strm0_ready         ( pe28__std__lane18_strm0_ready      ),      
               .std__pe28__lane18_strm0_cntl          ( std__pe28__lane18_strm0_cntl       ),      
               .std__pe28__lane18_strm0_data          ( std__pe28__lane18_strm0_data       ),      
               .std__pe28__lane18_strm0_data_valid    ( std__pe28__lane18_strm0_data_valid ),      
               .std__pe28__lane18_strm0_data_mask     ( std__pe28__lane18_strm0_data_mask  ),      

               .pe28__std__lane18_strm1_ready         ( pe28__std__lane18_strm1_ready      ),      
               .std__pe28__lane18_strm1_cntl          ( std__pe28__lane18_strm1_cntl       ),      
               .std__pe28__lane18_strm1_data          ( std__pe28__lane18_strm1_data       ),      
               .std__pe28__lane18_strm1_data_valid    ( std__pe28__lane18_strm1_data_valid ),      
               .std__pe28__lane18_strm1_data_mask     ( std__pe28__lane18_strm1_data_mask  ),      

               // PE 28, Lane 19                 
               .pe28__std__lane19_strm0_ready         ( pe28__std__lane19_strm0_ready      ),      
               .std__pe28__lane19_strm0_cntl          ( std__pe28__lane19_strm0_cntl       ),      
               .std__pe28__lane19_strm0_data          ( std__pe28__lane19_strm0_data       ),      
               .std__pe28__lane19_strm0_data_valid    ( std__pe28__lane19_strm0_data_valid ),      
               .std__pe28__lane19_strm0_data_mask     ( std__pe28__lane19_strm0_data_mask  ),      

               .pe28__std__lane19_strm1_ready         ( pe28__std__lane19_strm1_ready      ),      
               .std__pe28__lane19_strm1_cntl          ( std__pe28__lane19_strm1_cntl       ),      
               .std__pe28__lane19_strm1_data          ( std__pe28__lane19_strm1_data       ),      
               .std__pe28__lane19_strm1_data_valid    ( std__pe28__lane19_strm1_data_valid ),      
               .std__pe28__lane19_strm1_data_mask     ( std__pe28__lane19_strm1_data_mask  ),      

               // PE 28, Lane 20                 
               .pe28__std__lane20_strm0_ready         ( pe28__std__lane20_strm0_ready      ),      
               .std__pe28__lane20_strm0_cntl          ( std__pe28__lane20_strm0_cntl       ),      
               .std__pe28__lane20_strm0_data          ( std__pe28__lane20_strm0_data       ),      
               .std__pe28__lane20_strm0_data_valid    ( std__pe28__lane20_strm0_data_valid ),      
               .std__pe28__lane20_strm0_data_mask     ( std__pe28__lane20_strm0_data_mask  ),      

               .pe28__std__lane20_strm1_ready         ( pe28__std__lane20_strm1_ready      ),      
               .std__pe28__lane20_strm1_cntl          ( std__pe28__lane20_strm1_cntl       ),      
               .std__pe28__lane20_strm1_data          ( std__pe28__lane20_strm1_data       ),      
               .std__pe28__lane20_strm1_data_valid    ( std__pe28__lane20_strm1_data_valid ),      
               .std__pe28__lane20_strm1_data_mask     ( std__pe28__lane20_strm1_data_mask  ),      

               // PE 28, Lane 21                 
               .pe28__std__lane21_strm0_ready         ( pe28__std__lane21_strm0_ready      ),      
               .std__pe28__lane21_strm0_cntl          ( std__pe28__lane21_strm0_cntl       ),      
               .std__pe28__lane21_strm0_data          ( std__pe28__lane21_strm0_data       ),      
               .std__pe28__lane21_strm0_data_valid    ( std__pe28__lane21_strm0_data_valid ),      
               .std__pe28__lane21_strm0_data_mask     ( std__pe28__lane21_strm0_data_mask  ),      

               .pe28__std__lane21_strm1_ready         ( pe28__std__lane21_strm1_ready      ),      
               .std__pe28__lane21_strm1_cntl          ( std__pe28__lane21_strm1_cntl       ),      
               .std__pe28__lane21_strm1_data          ( std__pe28__lane21_strm1_data       ),      
               .std__pe28__lane21_strm1_data_valid    ( std__pe28__lane21_strm1_data_valid ),      
               .std__pe28__lane21_strm1_data_mask     ( std__pe28__lane21_strm1_data_mask  ),      

               // PE 28, Lane 22                 
               .pe28__std__lane22_strm0_ready         ( pe28__std__lane22_strm0_ready      ),      
               .std__pe28__lane22_strm0_cntl          ( std__pe28__lane22_strm0_cntl       ),      
               .std__pe28__lane22_strm0_data          ( std__pe28__lane22_strm0_data       ),      
               .std__pe28__lane22_strm0_data_valid    ( std__pe28__lane22_strm0_data_valid ),      
               .std__pe28__lane22_strm0_data_mask     ( std__pe28__lane22_strm0_data_mask  ),      

               .pe28__std__lane22_strm1_ready         ( pe28__std__lane22_strm1_ready      ),      
               .std__pe28__lane22_strm1_cntl          ( std__pe28__lane22_strm1_cntl       ),      
               .std__pe28__lane22_strm1_data          ( std__pe28__lane22_strm1_data       ),      
               .std__pe28__lane22_strm1_data_valid    ( std__pe28__lane22_strm1_data_valid ),      
               .std__pe28__lane22_strm1_data_mask     ( std__pe28__lane22_strm1_data_mask  ),      

               // PE 28, Lane 23                 
               .pe28__std__lane23_strm0_ready         ( pe28__std__lane23_strm0_ready      ),      
               .std__pe28__lane23_strm0_cntl          ( std__pe28__lane23_strm0_cntl       ),      
               .std__pe28__lane23_strm0_data          ( std__pe28__lane23_strm0_data       ),      
               .std__pe28__lane23_strm0_data_valid    ( std__pe28__lane23_strm0_data_valid ),      
               .std__pe28__lane23_strm0_data_mask     ( std__pe28__lane23_strm0_data_mask  ),      

               .pe28__std__lane23_strm1_ready         ( pe28__std__lane23_strm1_ready      ),      
               .std__pe28__lane23_strm1_cntl          ( std__pe28__lane23_strm1_cntl       ),      
               .std__pe28__lane23_strm1_data          ( std__pe28__lane23_strm1_data       ),      
               .std__pe28__lane23_strm1_data_valid    ( std__pe28__lane23_strm1_data_valid ),      
               .std__pe28__lane23_strm1_data_mask     ( std__pe28__lane23_strm1_data_mask  ),      

               // PE 28, Lane 24                 
               .pe28__std__lane24_strm0_ready         ( pe28__std__lane24_strm0_ready      ),      
               .std__pe28__lane24_strm0_cntl          ( std__pe28__lane24_strm0_cntl       ),      
               .std__pe28__lane24_strm0_data          ( std__pe28__lane24_strm0_data       ),      
               .std__pe28__lane24_strm0_data_valid    ( std__pe28__lane24_strm0_data_valid ),      
               .std__pe28__lane24_strm0_data_mask     ( std__pe28__lane24_strm0_data_mask  ),      

               .pe28__std__lane24_strm1_ready         ( pe28__std__lane24_strm1_ready      ),      
               .std__pe28__lane24_strm1_cntl          ( std__pe28__lane24_strm1_cntl       ),      
               .std__pe28__lane24_strm1_data          ( std__pe28__lane24_strm1_data       ),      
               .std__pe28__lane24_strm1_data_valid    ( std__pe28__lane24_strm1_data_valid ),      
               .std__pe28__lane24_strm1_data_mask     ( std__pe28__lane24_strm1_data_mask  ),      

               // PE 28, Lane 25                 
               .pe28__std__lane25_strm0_ready         ( pe28__std__lane25_strm0_ready      ),      
               .std__pe28__lane25_strm0_cntl          ( std__pe28__lane25_strm0_cntl       ),      
               .std__pe28__lane25_strm0_data          ( std__pe28__lane25_strm0_data       ),      
               .std__pe28__lane25_strm0_data_valid    ( std__pe28__lane25_strm0_data_valid ),      
               .std__pe28__lane25_strm0_data_mask     ( std__pe28__lane25_strm0_data_mask  ),      

               .pe28__std__lane25_strm1_ready         ( pe28__std__lane25_strm1_ready      ),      
               .std__pe28__lane25_strm1_cntl          ( std__pe28__lane25_strm1_cntl       ),      
               .std__pe28__lane25_strm1_data          ( std__pe28__lane25_strm1_data       ),      
               .std__pe28__lane25_strm1_data_valid    ( std__pe28__lane25_strm1_data_valid ),      
               .std__pe28__lane25_strm1_data_mask     ( std__pe28__lane25_strm1_data_mask  ),      

               // PE 28, Lane 26                 
               .pe28__std__lane26_strm0_ready         ( pe28__std__lane26_strm0_ready      ),      
               .std__pe28__lane26_strm0_cntl          ( std__pe28__lane26_strm0_cntl       ),      
               .std__pe28__lane26_strm0_data          ( std__pe28__lane26_strm0_data       ),      
               .std__pe28__lane26_strm0_data_valid    ( std__pe28__lane26_strm0_data_valid ),      
               .std__pe28__lane26_strm0_data_mask     ( std__pe28__lane26_strm0_data_mask  ),      

               .pe28__std__lane26_strm1_ready         ( pe28__std__lane26_strm1_ready      ),      
               .std__pe28__lane26_strm1_cntl          ( std__pe28__lane26_strm1_cntl       ),      
               .std__pe28__lane26_strm1_data          ( std__pe28__lane26_strm1_data       ),      
               .std__pe28__lane26_strm1_data_valid    ( std__pe28__lane26_strm1_data_valid ),      
               .std__pe28__lane26_strm1_data_mask     ( std__pe28__lane26_strm1_data_mask  ),      

               // PE 28, Lane 27                 
               .pe28__std__lane27_strm0_ready         ( pe28__std__lane27_strm0_ready      ),      
               .std__pe28__lane27_strm0_cntl          ( std__pe28__lane27_strm0_cntl       ),      
               .std__pe28__lane27_strm0_data          ( std__pe28__lane27_strm0_data       ),      
               .std__pe28__lane27_strm0_data_valid    ( std__pe28__lane27_strm0_data_valid ),      
               .std__pe28__lane27_strm0_data_mask     ( std__pe28__lane27_strm0_data_mask  ),      

               .pe28__std__lane27_strm1_ready         ( pe28__std__lane27_strm1_ready      ),      
               .std__pe28__lane27_strm1_cntl          ( std__pe28__lane27_strm1_cntl       ),      
               .std__pe28__lane27_strm1_data          ( std__pe28__lane27_strm1_data       ),      
               .std__pe28__lane27_strm1_data_valid    ( std__pe28__lane27_strm1_data_valid ),      
               .std__pe28__lane27_strm1_data_mask     ( std__pe28__lane27_strm1_data_mask  ),      

               // PE 28, Lane 28                 
               .pe28__std__lane28_strm0_ready         ( pe28__std__lane28_strm0_ready      ),      
               .std__pe28__lane28_strm0_cntl          ( std__pe28__lane28_strm0_cntl       ),      
               .std__pe28__lane28_strm0_data          ( std__pe28__lane28_strm0_data       ),      
               .std__pe28__lane28_strm0_data_valid    ( std__pe28__lane28_strm0_data_valid ),      
               .std__pe28__lane28_strm0_data_mask     ( std__pe28__lane28_strm0_data_mask  ),      

               .pe28__std__lane28_strm1_ready         ( pe28__std__lane28_strm1_ready      ),      
               .std__pe28__lane28_strm1_cntl          ( std__pe28__lane28_strm1_cntl       ),      
               .std__pe28__lane28_strm1_data          ( std__pe28__lane28_strm1_data       ),      
               .std__pe28__lane28_strm1_data_valid    ( std__pe28__lane28_strm1_data_valid ),      
               .std__pe28__lane28_strm1_data_mask     ( std__pe28__lane28_strm1_data_mask  ),      

               // PE 28, Lane 29                 
               .pe28__std__lane29_strm0_ready         ( pe28__std__lane29_strm0_ready      ),      
               .std__pe28__lane29_strm0_cntl          ( std__pe28__lane29_strm0_cntl       ),      
               .std__pe28__lane29_strm0_data          ( std__pe28__lane29_strm0_data       ),      
               .std__pe28__lane29_strm0_data_valid    ( std__pe28__lane29_strm0_data_valid ),      
               .std__pe28__lane29_strm0_data_mask     ( std__pe28__lane29_strm0_data_mask  ),      

               .pe28__std__lane29_strm1_ready         ( pe28__std__lane29_strm1_ready      ),      
               .std__pe28__lane29_strm1_cntl          ( std__pe28__lane29_strm1_cntl       ),      
               .std__pe28__lane29_strm1_data          ( std__pe28__lane29_strm1_data       ),      
               .std__pe28__lane29_strm1_data_valid    ( std__pe28__lane29_strm1_data_valid ),      
               .std__pe28__lane29_strm1_data_mask     ( std__pe28__lane29_strm1_data_mask  ),      

               // PE 28, Lane 30                 
               .pe28__std__lane30_strm0_ready         ( pe28__std__lane30_strm0_ready      ),      
               .std__pe28__lane30_strm0_cntl          ( std__pe28__lane30_strm0_cntl       ),      
               .std__pe28__lane30_strm0_data          ( std__pe28__lane30_strm0_data       ),      
               .std__pe28__lane30_strm0_data_valid    ( std__pe28__lane30_strm0_data_valid ),      
               .std__pe28__lane30_strm0_data_mask     ( std__pe28__lane30_strm0_data_mask  ),      

               .pe28__std__lane30_strm1_ready         ( pe28__std__lane30_strm1_ready      ),      
               .std__pe28__lane30_strm1_cntl          ( std__pe28__lane30_strm1_cntl       ),      
               .std__pe28__lane30_strm1_data          ( std__pe28__lane30_strm1_data       ),      
               .std__pe28__lane30_strm1_data_valid    ( std__pe28__lane30_strm1_data_valid ),      
               .std__pe28__lane30_strm1_data_mask     ( std__pe28__lane30_strm1_data_mask  ),      

               // PE 28, Lane 31                 
               .pe28__std__lane31_strm0_ready         ( pe28__std__lane31_strm0_ready      ),      
               .std__pe28__lane31_strm0_cntl          ( std__pe28__lane31_strm0_cntl       ),      
               .std__pe28__lane31_strm0_data          ( std__pe28__lane31_strm0_data       ),      
               .std__pe28__lane31_strm0_data_valid    ( std__pe28__lane31_strm0_data_valid ),      
               .std__pe28__lane31_strm0_data_mask     ( std__pe28__lane31_strm0_data_mask  ),      

               .pe28__std__lane31_strm1_ready         ( pe28__std__lane31_strm1_ready      ),      
               .std__pe28__lane31_strm1_cntl          ( std__pe28__lane31_strm1_cntl       ),      
               .std__pe28__lane31_strm1_data          ( std__pe28__lane31_strm1_data       ),      
               .std__pe28__lane31_strm1_data_valid    ( std__pe28__lane31_strm1_data_valid ),      
               .std__pe28__lane31_strm1_data_mask     ( std__pe28__lane31_strm1_data_mask  ),      

               // PE 29, Lane 0                 
               .pe29__std__lane0_strm0_ready         ( pe29__std__lane0_strm0_ready      ),      
               .std__pe29__lane0_strm0_cntl          ( std__pe29__lane0_strm0_cntl       ),      
               .std__pe29__lane0_strm0_data          ( std__pe29__lane0_strm0_data       ),      
               .std__pe29__lane0_strm0_data_valid    ( std__pe29__lane0_strm0_data_valid ),      
               .std__pe29__lane0_strm0_data_mask     ( std__pe29__lane0_strm0_data_mask  ),      

               .pe29__std__lane0_strm1_ready         ( pe29__std__lane0_strm1_ready      ),      
               .std__pe29__lane0_strm1_cntl          ( std__pe29__lane0_strm1_cntl       ),      
               .std__pe29__lane0_strm1_data          ( std__pe29__lane0_strm1_data       ),      
               .std__pe29__lane0_strm1_data_valid    ( std__pe29__lane0_strm1_data_valid ),      
               .std__pe29__lane0_strm1_data_mask     ( std__pe29__lane0_strm1_data_mask  ),      

               // PE 29, Lane 1                 
               .pe29__std__lane1_strm0_ready         ( pe29__std__lane1_strm0_ready      ),      
               .std__pe29__lane1_strm0_cntl          ( std__pe29__lane1_strm0_cntl       ),      
               .std__pe29__lane1_strm0_data          ( std__pe29__lane1_strm0_data       ),      
               .std__pe29__lane1_strm0_data_valid    ( std__pe29__lane1_strm0_data_valid ),      
               .std__pe29__lane1_strm0_data_mask     ( std__pe29__lane1_strm0_data_mask  ),      

               .pe29__std__lane1_strm1_ready         ( pe29__std__lane1_strm1_ready      ),      
               .std__pe29__lane1_strm1_cntl          ( std__pe29__lane1_strm1_cntl       ),      
               .std__pe29__lane1_strm1_data          ( std__pe29__lane1_strm1_data       ),      
               .std__pe29__lane1_strm1_data_valid    ( std__pe29__lane1_strm1_data_valid ),      
               .std__pe29__lane1_strm1_data_mask     ( std__pe29__lane1_strm1_data_mask  ),      

               // PE 29, Lane 2                 
               .pe29__std__lane2_strm0_ready         ( pe29__std__lane2_strm0_ready      ),      
               .std__pe29__lane2_strm0_cntl          ( std__pe29__lane2_strm0_cntl       ),      
               .std__pe29__lane2_strm0_data          ( std__pe29__lane2_strm0_data       ),      
               .std__pe29__lane2_strm0_data_valid    ( std__pe29__lane2_strm0_data_valid ),      
               .std__pe29__lane2_strm0_data_mask     ( std__pe29__lane2_strm0_data_mask  ),      

               .pe29__std__lane2_strm1_ready         ( pe29__std__lane2_strm1_ready      ),      
               .std__pe29__lane2_strm1_cntl          ( std__pe29__lane2_strm1_cntl       ),      
               .std__pe29__lane2_strm1_data          ( std__pe29__lane2_strm1_data       ),      
               .std__pe29__lane2_strm1_data_valid    ( std__pe29__lane2_strm1_data_valid ),      
               .std__pe29__lane2_strm1_data_mask     ( std__pe29__lane2_strm1_data_mask  ),      

               // PE 29, Lane 3                 
               .pe29__std__lane3_strm0_ready         ( pe29__std__lane3_strm0_ready      ),      
               .std__pe29__lane3_strm0_cntl          ( std__pe29__lane3_strm0_cntl       ),      
               .std__pe29__lane3_strm0_data          ( std__pe29__lane3_strm0_data       ),      
               .std__pe29__lane3_strm0_data_valid    ( std__pe29__lane3_strm0_data_valid ),      
               .std__pe29__lane3_strm0_data_mask     ( std__pe29__lane3_strm0_data_mask  ),      

               .pe29__std__lane3_strm1_ready         ( pe29__std__lane3_strm1_ready      ),      
               .std__pe29__lane3_strm1_cntl          ( std__pe29__lane3_strm1_cntl       ),      
               .std__pe29__lane3_strm1_data          ( std__pe29__lane3_strm1_data       ),      
               .std__pe29__lane3_strm1_data_valid    ( std__pe29__lane3_strm1_data_valid ),      
               .std__pe29__lane3_strm1_data_mask     ( std__pe29__lane3_strm1_data_mask  ),      

               // PE 29, Lane 4                 
               .pe29__std__lane4_strm0_ready         ( pe29__std__lane4_strm0_ready      ),      
               .std__pe29__lane4_strm0_cntl          ( std__pe29__lane4_strm0_cntl       ),      
               .std__pe29__lane4_strm0_data          ( std__pe29__lane4_strm0_data       ),      
               .std__pe29__lane4_strm0_data_valid    ( std__pe29__lane4_strm0_data_valid ),      
               .std__pe29__lane4_strm0_data_mask     ( std__pe29__lane4_strm0_data_mask  ),      

               .pe29__std__lane4_strm1_ready         ( pe29__std__lane4_strm1_ready      ),      
               .std__pe29__lane4_strm1_cntl          ( std__pe29__lane4_strm1_cntl       ),      
               .std__pe29__lane4_strm1_data          ( std__pe29__lane4_strm1_data       ),      
               .std__pe29__lane4_strm1_data_valid    ( std__pe29__lane4_strm1_data_valid ),      
               .std__pe29__lane4_strm1_data_mask     ( std__pe29__lane4_strm1_data_mask  ),      

               // PE 29, Lane 5                 
               .pe29__std__lane5_strm0_ready         ( pe29__std__lane5_strm0_ready      ),      
               .std__pe29__lane5_strm0_cntl          ( std__pe29__lane5_strm0_cntl       ),      
               .std__pe29__lane5_strm0_data          ( std__pe29__lane5_strm0_data       ),      
               .std__pe29__lane5_strm0_data_valid    ( std__pe29__lane5_strm0_data_valid ),      
               .std__pe29__lane5_strm0_data_mask     ( std__pe29__lane5_strm0_data_mask  ),      

               .pe29__std__lane5_strm1_ready         ( pe29__std__lane5_strm1_ready      ),      
               .std__pe29__lane5_strm1_cntl          ( std__pe29__lane5_strm1_cntl       ),      
               .std__pe29__lane5_strm1_data          ( std__pe29__lane5_strm1_data       ),      
               .std__pe29__lane5_strm1_data_valid    ( std__pe29__lane5_strm1_data_valid ),      
               .std__pe29__lane5_strm1_data_mask     ( std__pe29__lane5_strm1_data_mask  ),      

               // PE 29, Lane 6                 
               .pe29__std__lane6_strm0_ready         ( pe29__std__lane6_strm0_ready      ),      
               .std__pe29__lane6_strm0_cntl          ( std__pe29__lane6_strm0_cntl       ),      
               .std__pe29__lane6_strm0_data          ( std__pe29__lane6_strm0_data       ),      
               .std__pe29__lane6_strm0_data_valid    ( std__pe29__lane6_strm0_data_valid ),      
               .std__pe29__lane6_strm0_data_mask     ( std__pe29__lane6_strm0_data_mask  ),      

               .pe29__std__lane6_strm1_ready         ( pe29__std__lane6_strm1_ready      ),      
               .std__pe29__lane6_strm1_cntl          ( std__pe29__lane6_strm1_cntl       ),      
               .std__pe29__lane6_strm1_data          ( std__pe29__lane6_strm1_data       ),      
               .std__pe29__lane6_strm1_data_valid    ( std__pe29__lane6_strm1_data_valid ),      
               .std__pe29__lane6_strm1_data_mask     ( std__pe29__lane6_strm1_data_mask  ),      

               // PE 29, Lane 7                 
               .pe29__std__lane7_strm0_ready         ( pe29__std__lane7_strm0_ready      ),      
               .std__pe29__lane7_strm0_cntl          ( std__pe29__lane7_strm0_cntl       ),      
               .std__pe29__lane7_strm0_data          ( std__pe29__lane7_strm0_data       ),      
               .std__pe29__lane7_strm0_data_valid    ( std__pe29__lane7_strm0_data_valid ),      
               .std__pe29__lane7_strm0_data_mask     ( std__pe29__lane7_strm0_data_mask  ),      

               .pe29__std__lane7_strm1_ready         ( pe29__std__lane7_strm1_ready      ),      
               .std__pe29__lane7_strm1_cntl          ( std__pe29__lane7_strm1_cntl       ),      
               .std__pe29__lane7_strm1_data          ( std__pe29__lane7_strm1_data       ),      
               .std__pe29__lane7_strm1_data_valid    ( std__pe29__lane7_strm1_data_valid ),      
               .std__pe29__lane7_strm1_data_mask     ( std__pe29__lane7_strm1_data_mask  ),      

               // PE 29, Lane 8                 
               .pe29__std__lane8_strm0_ready         ( pe29__std__lane8_strm0_ready      ),      
               .std__pe29__lane8_strm0_cntl          ( std__pe29__lane8_strm0_cntl       ),      
               .std__pe29__lane8_strm0_data          ( std__pe29__lane8_strm0_data       ),      
               .std__pe29__lane8_strm0_data_valid    ( std__pe29__lane8_strm0_data_valid ),      
               .std__pe29__lane8_strm0_data_mask     ( std__pe29__lane8_strm0_data_mask  ),      

               .pe29__std__lane8_strm1_ready         ( pe29__std__lane8_strm1_ready      ),      
               .std__pe29__lane8_strm1_cntl          ( std__pe29__lane8_strm1_cntl       ),      
               .std__pe29__lane8_strm1_data          ( std__pe29__lane8_strm1_data       ),      
               .std__pe29__lane8_strm1_data_valid    ( std__pe29__lane8_strm1_data_valid ),      
               .std__pe29__lane8_strm1_data_mask     ( std__pe29__lane8_strm1_data_mask  ),      

               // PE 29, Lane 9                 
               .pe29__std__lane9_strm0_ready         ( pe29__std__lane9_strm0_ready      ),      
               .std__pe29__lane9_strm0_cntl          ( std__pe29__lane9_strm0_cntl       ),      
               .std__pe29__lane9_strm0_data          ( std__pe29__lane9_strm0_data       ),      
               .std__pe29__lane9_strm0_data_valid    ( std__pe29__lane9_strm0_data_valid ),      
               .std__pe29__lane9_strm0_data_mask     ( std__pe29__lane9_strm0_data_mask  ),      

               .pe29__std__lane9_strm1_ready         ( pe29__std__lane9_strm1_ready      ),      
               .std__pe29__lane9_strm1_cntl          ( std__pe29__lane9_strm1_cntl       ),      
               .std__pe29__lane9_strm1_data          ( std__pe29__lane9_strm1_data       ),      
               .std__pe29__lane9_strm1_data_valid    ( std__pe29__lane9_strm1_data_valid ),      
               .std__pe29__lane9_strm1_data_mask     ( std__pe29__lane9_strm1_data_mask  ),      

               // PE 29, Lane 10                 
               .pe29__std__lane10_strm0_ready         ( pe29__std__lane10_strm0_ready      ),      
               .std__pe29__lane10_strm0_cntl          ( std__pe29__lane10_strm0_cntl       ),      
               .std__pe29__lane10_strm0_data          ( std__pe29__lane10_strm0_data       ),      
               .std__pe29__lane10_strm0_data_valid    ( std__pe29__lane10_strm0_data_valid ),      
               .std__pe29__lane10_strm0_data_mask     ( std__pe29__lane10_strm0_data_mask  ),      

               .pe29__std__lane10_strm1_ready         ( pe29__std__lane10_strm1_ready      ),      
               .std__pe29__lane10_strm1_cntl          ( std__pe29__lane10_strm1_cntl       ),      
               .std__pe29__lane10_strm1_data          ( std__pe29__lane10_strm1_data       ),      
               .std__pe29__lane10_strm1_data_valid    ( std__pe29__lane10_strm1_data_valid ),      
               .std__pe29__lane10_strm1_data_mask     ( std__pe29__lane10_strm1_data_mask  ),      

               // PE 29, Lane 11                 
               .pe29__std__lane11_strm0_ready         ( pe29__std__lane11_strm0_ready      ),      
               .std__pe29__lane11_strm0_cntl          ( std__pe29__lane11_strm0_cntl       ),      
               .std__pe29__lane11_strm0_data          ( std__pe29__lane11_strm0_data       ),      
               .std__pe29__lane11_strm0_data_valid    ( std__pe29__lane11_strm0_data_valid ),      
               .std__pe29__lane11_strm0_data_mask     ( std__pe29__lane11_strm0_data_mask  ),      

               .pe29__std__lane11_strm1_ready         ( pe29__std__lane11_strm1_ready      ),      
               .std__pe29__lane11_strm1_cntl          ( std__pe29__lane11_strm1_cntl       ),      
               .std__pe29__lane11_strm1_data          ( std__pe29__lane11_strm1_data       ),      
               .std__pe29__lane11_strm1_data_valid    ( std__pe29__lane11_strm1_data_valid ),      
               .std__pe29__lane11_strm1_data_mask     ( std__pe29__lane11_strm1_data_mask  ),      

               // PE 29, Lane 12                 
               .pe29__std__lane12_strm0_ready         ( pe29__std__lane12_strm0_ready      ),      
               .std__pe29__lane12_strm0_cntl          ( std__pe29__lane12_strm0_cntl       ),      
               .std__pe29__lane12_strm0_data          ( std__pe29__lane12_strm0_data       ),      
               .std__pe29__lane12_strm0_data_valid    ( std__pe29__lane12_strm0_data_valid ),      
               .std__pe29__lane12_strm0_data_mask     ( std__pe29__lane12_strm0_data_mask  ),      

               .pe29__std__lane12_strm1_ready         ( pe29__std__lane12_strm1_ready      ),      
               .std__pe29__lane12_strm1_cntl          ( std__pe29__lane12_strm1_cntl       ),      
               .std__pe29__lane12_strm1_data          ( std__pe29__lane12_strm1_data       ),      
               .std__pe29__lane12_strm1_data_valid    ( std__pe29__lane12_strm1_data_valid ),      
               .std__pe29__lane12_strm1_data_mask     ( std__pe29__lane12_strm1_data_mask  ),      

               // PE 29, Lane 13                 
               .pe29__std__lane13_strm0_ready         ( pe29__std__lane13_strm0_ready      ),      
               .std__pe29__lane13_strm0_cntl          ( std__pe29__lane13_strm0_cntl       ),      
               .std__pe29__lane13_strm0_data          ( std__pe29__lane13_strm0_data       ),      
               .std__pe29__lane13_strm0_data_valid    ( std__pe29__lane13_strm0_data_valid ),      
               .std__pe29__lane13_strm0_data_mask     ( std__pe29__lane13_strm0_data_mask  ),      

               .pe29__std__lane13_strm1_ready         ( pe29__std__lane13_strm1_ready      ),      
               .std__pe29__lane13_strm1_cntl          ( std__pe29__lane13_strm1_cntl       ),      
               .std__pe29__lane13_strm1_data          ( std__pe29__lane13_strm1_data       ),      
               .std__pe29__lane13_strm1_data_valid    ( std__pe29__lane13_strm1_data_valid ),      
               .std__pe29__lane13_strm1_data_mask     ( std__pe29__lane13_strm1_data_mask  ),      

               // PE 29, Lane 14                 
               .pe29__std__lane14_strm0_ready         ( pe29__std__lane14_strm0_ready      ),      
               .std__pe29__lane14_strm0_cntl          ( std__pe29__lane14_strm0_cntl       ),      
               .std__pe29__lane14_strm0_data          ( std__pe29__lane14_strm0_data       ),      
               .std__pe29__lane14_strm0_data_valid    ( std__pe29__lane14_strm0_data_valid ),      
               .std__pe29__lane14_strm0_data_mask     ( std__pe29__lane14_strm0_data_mask  ),      

               .pe29__std__lane14_strm1_ready         ( pe29__std__lane14_strm1_ready      ),      
               .std__pe29__lane14_strm1_cntl          ( std__pe29__lane14_strm1_cntl       ),      
               .std__pe29__lane14_strm1_data          ( std__pe29__lane14_strm1_data       ),      
               .std__pe29__lane14_strm1_data_valid    ( std__pe29__lane14_strm1_data_valid ),      
               .std__pe29__lane14_strm1_data_mask     ( std__pe29__lane14_strm1_data_mask  ),      

               // PE 29, Lane 15                 
               .pe29__std__lane15_strm0_ready         ( pe29__std__lane15_strm0_ready      ),      
               .std__pe29__lane15_strm0_cntl          ( std__pe29__lane15_strm0_cntl       ),      
               .std__pe29__lane15_strm0_data          ( std__pe29__lane15_strm0_data       ),      
               .std__pe29__lane15_strm0_data_valid    ( std__pe29__lane15_strm0_data_valid ),      
               .std__pe29__lane15_strm0_data_mask     ( std__pe29__lane15_strm0_data_mask  ),      

               .pe29__std__lane15_strm1_ready         ( pe29__std__lane15_strm1_ready      ),      
               .std__pe29__lane15_strm1_cntl          ( std__pe29__lane15_strm1_cntl       ),      
               .std__pe29__lane15_strm1_data          ( std__pe29__lane15_strm1_data       ),      
               .std__pe29__lane15_strm1_data_valid    ( std__pe29__lane15_strm1_data_valid ),      
               .std__pe29__lane15_strm1_data_mask     ( std__pe29__lane15_strm1_data_mask  ),      

               // PE 29, Lane 16                 
               .pe29__std__lane16_strm0_ready         ( pe29__std__lane16_strm0_ready      ),      
               .std__pe29__lane16_strm0_cntl          ( std__pe29__lane16_strm0_cntl       ),      
               .std__pe29__lane16_strm0_data          ( std__pe29__lane16_strm0_data       ),      
               .std__pe29__lane16_strm0_data_valid    ( std__pe29__lane16_strm0_data_valid ),      
               .std__pe29__lane16_strm0_data_mask     ( std__pe29__lane16_strm0_data_mask  ),      

               .pe29__std__lane16_strm1_ready         ( pe29__std__lane16_strm1_ready      ),      
               .std__pe29__lane16_strm1_cntl          ( std__pe29__lane16_strm1_cntl       ),      
               .std__pe29__lane16_strm1_data          ( std__pe29__lane16_strm1_data       ),      
               .std__pe29__lane16_strm1_data_valid    ( std__pe29__lane16_strm1_data_valid ),      
               .std__pe29__lane16_strm1_data_mask     ( std__pe29__lane16_strm1_data_mask  ),      

               // PE 29, Lane 17                 
               .pe29__std__lane17_strm0_ready         ( pe29__std__lane17_strm0_ready      ),      
               .std__pe29__lane17_strm0_cntl          ( std__pe29__lane17_strm0_cntl       ),      
               .std__pe29__lane17_strm0_data          ( std__pe29__lane17_strm0_data       ),      
               .std__pe29__lane17_strm0_data_valid    ( std__pe29__lane17_strm0_data_valid ),      
               .std__pe29__lane17_strm0_data_mask     ( std__pe29__lane17_strm0_data_mask  ),      

               .pe29__std__lane17_strm1_ready         ( pe29__std__lane17_strm1_ready      ),      
               .std__pe29__lane17_strm1_cntl          ( std__pe29__lane17_strm1_cntl       ),      
               .std__pe29__lane17_strm1_data          ( std__pe29__lane17_strm1_data       ),      
               .std__pe29__lane17_strm1_data_valid    ( std__pe29__lane17_strm1_data_valid ),      
               .std__pe29__lane17_strm1_data_mask     ( std__pe29__lane17_strm1_data_mask  ),      

               // PE 29, Lane 18                 
               .pe29__std__lane18_strm0_ready         ( pe29__std__lane18_strm0_ready      ),      
               .std__pe29__lane18_strm0_cntl          ( std__pe29__lane18_strm0_cntl       ),      
               .std__pe29__lane18_strm0_data          ( std__pe29__lane18_strm0_data       ),      
               .std__pe29__lane18_strm0_data_valid    ( std__pe29__lane18_strm0_data_valid ),      
               .std__pe29__lane18_strm0_data_mask     ( std__pe29__lane18_strm0_data_mask  ),      

               .pe29__std__lane18_strm1_ready         ( pe29__std__lane18_strm1_ready      ),      
               .std__pe29__lane18_strm1_cntl          ( std__pe29__lane18_strm1_cntl       ),      
               .std__pe29__lane18_strm1_data          ( std__pe29__lane18_strm1_data       ),      
               .std__pe29__lane18_strm1_data_valid    ( std__pe29__lane18_strm1_data_valid ),      
               .std__pe29__lane18_strm1_data_mask     ( std__pe29__lane18_strm1_data_mask  ),      

               // PE 29, Lane 19                 
               .pe29__std__lane19_strm0_ready         ( pe29__std__lane19_strm0_ready      ),      
               .std__pe29__lane19_strm0_cntl          ( std__pe29__lane19_strm0_cntl       ),      
               .std__pe29__lane19_strm0_data          ( std__pe29__lane19_strm0_data       ),      
               .std__pe29__lane19_strm0_data_valid    ( std__pe29__lane19_strm0_data_valid ),      
               .std__pe29__lane19_strm0_data_mask     ( std__pe29__lane19_strm0_data_mask  ),      

               .pe29__std__lane19_strm1_ready         ( pe29__std__lane19_strm1_ready      ),      
               .std__pe29__lane19_strm1_cntl          ( std__pe29__lane19_strm1_cntl       ),      
               .std__pe29__lane19_strm1_data          ( std__pe29__lane19_strm1_data       ),      
               .std__pe29__lane19_strm1_data_valid    ( std__pe29__lane19_strm1_data_valid ),      
               .std__pe29__lane19_strm1_data_mask     ( std__pe29__lane19_strm1_data_mask  ),      

               // PE 29, Lane 20                 
               .pe29__std__lane20_strm0_ready         ( pe29__std__lane20_strm0_ready      ),      
               .std__pe29__lane20_strm0_cntl          ( std__pe29__lane20_strm0_cntl       ),      
               .std__pe29__lane20_strm0_data          ( std__pe29__lane20_strm0_data       ),      
               .std__pe29__lane20_strm0_data_valid    ( std__pe29__lane20_strm0_data_valid ),      
               .std__pe29__lane20_strm0_data_mask     ( std__pe29__lane20_strm0_data_mask  ),      

               .pe29__std__lane20_strm1_ready         ( pe29__std__lane20_strm1_ready      ),      
               .std__pe29__lane20_strm1_cntl          ( std__pe29__lane20_strm1_cntl       ),      
               .std__pe29__lane20_strm1_data          ( std__pe29__lane20_strm1_data       ),      
               .std__pe29__lane20_strm1_data_valid    ( std__pe29__lane20_strm1_data_valid ),      
               .std__pe29__lane20_strm1_data_mask     ( std__pe29__lane20_strm1_data_mask  ),      

               // PE 29, Lane 21                 
               .pe29__std__lane21_strm0_ready         ( pe29__std__lane21_strm0_ready      ),      
               .std__pe29__lane21_strm0_cntl          ( std__pe29__lane21_strm0_cntl       ),      
               .std__pe29__lane21_strm0_data          ( std__pe29__lane21_strm0_data       ),      
               .std__pe29__lane21_strm0_data_valid    ( std__pe29__lane21_strm0_data_valid ),      
               .std__pe29__lane21_strm0_data_mask     ( std__pe29__lane21_strm0_data_mask  ),      

               .pe29__std__lane21_strm1_ready         ( pe29__std__lane21_strm1_ready      ),      
               .std__pe29__lane21_strm1_cntl          ( std__pe29__lane21_strm1_cntl       ),      
               .std__pe29__lane21_strm1_data          ( std__pe29__lane21_strm1_data       ),      
               .std__pe29__lane21_strm1_data_valid    ( std__pe29__lane21_strm1_data_valid ),      
               .std__pe29__lane21_strm1_data_mask     ( std__pe29__lane21_strm1_data_mask  ),      

               // PE 29, Lane 22                 
               .pe29__std__lane22_strm0_ready         ( pe29__std__lane22_strm0_ready      ),      
               .std__pe29__lane22_strm0_cntl          ( std__pe29__lane22_strm0_cntl       ),      
               .std__pe29__lane22_strm0_data          ( std__pe29__lane22_strm0_data       ),      
               .std__pe29__lane22_strm0_data_valid    ( std__pe29__lane22_strm0_data_valid ),      
               .std__pe29__lane22_strm0_data_mask     ( std__pe29__lane22_strm0_data_mask  ),      

               .pe29__std__lane22_strm1_ready         ( pe29__std__lane22_strm1_ready      ),      
               .std__pe29__lane22_strm1_cntl          ( std__pe29__lane22_strm1_cntl       ),      
               .std__pe29__lane22_strm1_data          ( std__pe29__lane22_strm1_data       ),      
               .std__pe29__lane22_strm1_data_valid    ( std__pe29__lane22_strm1_data_valid ),      
               .std__pe29__lane22_strm1_data_mask     ( std__pe29__lane22_strm1_data_mask  ),      

               // PE 29, Lane 23                 
               .pe29__std__lane23_strm0_ready         ( pe29__std__lane23_strm0_ready      ),      
               .std__pe29__lane23_strm0_cntl          ( std__pe29__lane23_strm0_cntl       ),      
               .std__pe29__lane23_strm0_data          ( std__pe29__lane23_strm0_data       ),      
               .std__pe29__lane23_strm0_data_valid    ( std__pe29__lane23_strm0_data_valid ),      
               .std__pe29__lane23_strm0_data_mask     ( std__pe29__lane23_strm0_data_mask  ),      

               .pe29__std__lane23_strm1_ready         ( pe29__std__lane23_strm1_ready      ),      
               .std__pe29__lane23_strm1_cntl          ( std__pe29__lane23_strm1_cntl       ),      
               .std__pe29__lane23_strm1_data          ( std__pe29__lane23_strm1_data       ),      
               .std__pe29__lane23_strm1_data_valid    ( std__pe29__lane23_strm1_data_valid ),      
               .std__pe29__lane23_strm1_data_mask     ( std__pe29__lane23_strm1_data_mask  ),      

               // PE 29, Lane 24                 
               .pe29__std__lane24_strm0_ready         ( pe29__std__lane24_strm0_ready      ),      
               .std__pe29__lane24_strm0_cntl          ( std__pe29__lane24_strm0_cntl       ),      
               .std__pe29__lane24_strm0_data          ( std__pe29__lane24_strm0_data       ),      
               .std__pe29__lane24_strm0_data_valid    ( std__pe29__lane24_strm0_data_valid ),      
               .std__pe29__lane24_strm0_data_mask     ( std__pe29__lane24_strm0_data_mask  ),      

               .pe29__std__lane24_strm1_ready         ( pe29__std__lane24_strm1_ready      ),      
               .std__pe29__lane24_strm1_cntl          ( std__pe29__lane24_strm1_cntl       ),      
               .std__pe29__lane24_strm1_data          ( std__pe29__lane24_strm1_data       ),      
               .std__pe29__lane24_strm1_data_valid    ( std__pe29__lane24_strm1_data_valid ),      
               .std__pe29__lane24_strm1_data_mask     ( std__pe29__lane24_strm1_data_mask  ),      

               // PE 29, Lane 25                 
               .pe29__std__lane25_strm0_ready         ( pe29__std__lane25_strm0_ready      ),      
               .std__pe29__lane25_strm0_cntl          ( std__pe29__lane25_strm0_cntl       ),      
               .std__pe29__lane25_strm0_data          ( std__pe29__lane25_strm0_data       ),      
               .std__pe29__lane25_strm0_data_valid    ( std__pe29__lane25_strm0_data_valid ),      
               .std__pe29__lane25_strm0_data_mask     ( std__pe29__lane25_strm0_data_mask  ),      

               .pe29__std__lane25_strm1_ready         ( pe29__std__lane25_strm1_ready      ),      
               .std__pe29__lane25_strm1_cntl          ( std__pe29__lane25_strm1_cntl       ),      
               .std__pe29__lane25_strm1_data          ( std__pe29__lane25_strm1_data       ),      
               .std__pe29__lane25_strm1_data_valid    ( std__pe29__lane25_strm1_data_valid ),      
               .std__pe29__lane25_strm1_data_mask     ( std__pe29__lane25_strm1_data_mask  ),      

               // PE 29, Lane 26                 
               .pe29__std__lane26_strm0_ready         ( pe29__std__lane26_strm0_ready      ),      
               .std__pe29__lane26_strm0_cntl          ( std__pe29__lane26_strm0_cntl       ),      
               .std__pe29__lane26_strm0_data          ( std__pe29__lane26_strm0_data       ),      
               .std__pe29__lane26_strm0_data_valid    ( std__pe29__lane26_strm0_data_valid ),      
               .std__pe29__lane26_strm0_data_mask     ( std__pe29__lane26_strm0_data_mask  ),      

               .pe29__std__lane26_strm1_ready         ( pe29__std__lane26_strm1_ready      ),      
               .std__pe29__lane26_strm1_cntl          ( std__pe29__lane26_strm1_cntl       ),      
               .std__pe29__lane26_strm1_data          ( std__pe29__lane26_strm1_data       ),      
               .std__pe29__lane26_strm1_data_valid    ( std__pe29__lane26_strm1_data_valid ),      
               .std__pe29__lane26_strm1_data_mask     ( std__pe29__lane26_strm1_data_mask  ),      

               // PE 29, Lane 27                 
               .pe29__std__lane27_strm0_ready         ( pe29__std__lane27_strm0_ready      ),      
               .std__pe29__lane27_strm0_cntl          ( std__pe29__lane27_strm0_cntl       ),      
               .std__pe29__lane27_strm0_data          ( std__pe29__lane27_strm0_data       ),      
               .std__pe29__lane27_strm0_data_valid    ( std__pe29__lane27_strm0_data_valid ),      
               .std__pe29__lane27_strm0_data_mask     ( std__pe29__lane27_strm0_data_mask  ),      

               .pe29__std__lane27_strm1_ready         ( pe29__std__lane27_strm1_ready      ),      
               .std__pe29__lane27_strm1_cntl          ( std__pe29__lane27_strm1_cntl       ),      
               .std__pe29__lane27_strm1_data          ( std__pe29__lane27_strm1_data       ),      
               .std__pe29__lane27_strm1_data_valid    ( std__pe29__lane27_strm1_data_valid ),      
               .std__pe29__lane27_strm1_data_mask     ( std__pe29__lane27_strm1_data_mask  ),      

               // PE 29, Lane 28                 
               .pe29__std__lane28_strm0_ready         ( pe29__std__lane28_strm0_ready      ),      
               .std__pe29__lane28_strm0_cntl          ( std__pe29__lane28_strm0_cntl       ),      
               .std__pe29__lane28_strm0_data          ( std__pe29__lane28_strm0_data       ),      
               .std__pe29__lane28_strm0_data_valid    ( std__pe29__lane28_strm0_data_valid ),      
               .std__pe29__lane28_strm0_data_mask     ( std__pe29__lane28_strm0_data_mask  ),      

               .pe29__std__lane28_strm1_ready         ( pe29__std__lane28_strm1_ready      ),      
               .std__pe29__lane28_strm1_cntl          ( std__pe29__lane28_strm1_cntl       ),      
               .std__pe29__lane28_strm1_data          ( std__pe29__lane28_strm1_data       ),      
               .std__pe29__lane28_strm1_data_valid    ( std__pe29__lane28_strm1_data_valid ),      
               .std__pe29__lane28_strm1_data_mask     ( std__pe29__lane28_strm1_data_mask  ),      

               // PE 29, Lane 29                 
               .pe29__std__lane29_strm0_ready         ( pe29__std__lane29_strm0_ready      ),      
               .std__pe29__lane29_strm0_cntl          ( std__pe29__lane29_strm0_cntl       ),      
               .std__pe29__lane29_strm0_data          ( std__pe29__lane29_strm0_data       ),      
               .std__pe29__lane29_strm0_data_valid    ( std__pe29__lane29_strm0_data_valid ),      
               .std__pe29__lane29_strm0_data_mask     ( std__pe29__lane29_strm0_data_mask  ),      

               .pe29__std__lane29_strm1_ready         ( pe29__std__lane29_strm1_ready      ),      
               .std__pe29__lane29_strm1_cntl          ( std__pe29__lane29_strm1_cntl       ),      
               .std__pe29__lane29_strm1_data          ( std__pe29__lane29_strm1_data       ),      
               .std__pe29__lane29_strm1_data_valid    ( std__pe29__lane29_strm1_data_valid ),      
               .std__pe29__lane29_strm1_data_mask     ( std__pe29__lane29_strm1_data_mask  ),      

               // PE 29, Lane 30                 
               .pe29__std__lane30_strm0_ready         ( pe29__std__lane30_strm0_ready      ),      
               .std__pe29__lane30_strm0_cntl          ( std__pe29__lane30_strm0_cntl       ),      
               .std__pe29__lane30_strm0_data          ( std__pe29__lane30_strm0_data       ),      
               .std__pe29__lane30_strm0_data_valid    ( std__pe29__lane30_strm0_data_valid ),      
               .std__pe29__lane30_strm0_data_mask     ( std__pe29__lane30_strm0_data_mask  ),      

               .pe29__std__lane30_strm1_ready         ( pe29__std__lane30_strm1_ready      ),      
               .std__pe29__lane30_strm1_cntl          ( std__pe29__lane30_strm1_cntl       ),      
               .std__pe29__lane30_strm1_data          ( std__pe29__lane30_strm1_data       ),      
               .std__pe29__lane30_strm1_data_valid    ( std__pe29__lane30_strm1_data_valid ),      
               .std__pe29__lane30_strm1_data_mask     ( std__pe29__lane30_strm1_data_mask  ),      

               // PE 29, Lane 31                 
               .pe29__std__lane31_strm0_ready         ( pe29__std__lane31_strm0_ready      ),      
               .std__pe29__lane31_strm0_cntl          ( std__pe29__lane31_strm0_cntl       ),      
               .std__pe29__lane31_strm0_data          ( std__pe29__lane31_strm0_data       ),      
               .std__pe29__lane31_strm0_data_valid    ( std__pe29__lane31_strm0_data_valid ),      
               .std__pe29__lane31_strm0_data_mask     ( std__pe29__lane31_strm0_data_mask  ),      

               .pe29__std__lane31_strm1_ready         ( pe29__std__lane31_strm1_ready      ),      
               .std__pe29__lane31_strm1_cntl          ( std__pe29__lane31_strm1_cntl       ),      
               .std__pe29__lane31_strm1_data          ( std__pe29__lane31_strm1_data       ),      
               .std__pe29__lane31_strm1_data_valid    ( std__pe29__lane31_strm1_data_valid ),      
               .std__pe29__lane31_strm1_data_mask     ( std__pe29__lane31_strm1_data_mask  ),      

               // PE 30, Lane 0                 
               .pe30__std__lane0_strm0_ready         ( pe30__std__lane0_strm0_ready      ),      
               .std__pe30__lane0_strm0_cntl          ( std__pe30__lane0_strm0_cntl       ),      
               .std__pe30__lane0_strm0_data          ( std__pe30__lane0_strm0_data       ),      
               .std__pe30__lane0_strm0_data_valid    ( std__pe30__lane0_strm0_data_valid ),      
               .std__pe30__lane0_strm0_data_mask     ( std__pe30__lane0_strm0_data_mask  ),      

               .pe30__std__lane0_strm1_ready         ( pe30__std__lane0_strm1_ready      ),      
               .std__pe30__lane0_strm1_cntl          ( std__pe30__lane0_strm1_cntl       ),      
               .std__pe30__lane0_strm1_data          ( std__pe30__lane0_strm1_data       ),      
               .std__pe30__lane0_strm1_data_valid    ( std__pe30__lane0_strm1_data_valid ),      
               .std__pe30__lane0_strm1_data_mask     ( std__pe30__lane0_strm1_data_mask  ),      

               // PE 30, Lane 1                 
               .pe30__std__lane1_strm0_ready         ( pe30__std__lane1_strm0_ready      ),      
               .std__pe30__lane1_strm0_cntl          ( std__pe30__lane1_strm0_cntl       ),      
               .std__pe30__lane1_strm0_data          ( std__pe30__lane1_strm0_data       ),      
               .std__pe30__lane1_strm0_data_valid    ( std__pe30__lane1_strm0_data_valid ),      
               .std__pe30__lane1_strm0_data_mask     ( std__pe30__lane1_strm0_data_mask  ),      

               .pe30__std__lane1_strm1_ready         ( pe30__std__lane1_strm1_ready      ),      
               .std__pe30__lane1_strm1_cntl          ( std__pe30__lane1_strm1_cntl       ),      
               .std__pe30__lane1_strm1_data          ( std__pe30__lane1_strm1_data       ),      
               .std__pe30__lane1_strm1_data_valid    ( std__pe30__lane1_strm1_data_valid ),      
               .std__pe30__lane1_strm1_data_mask     ( std__pe30__lane1_strm1_data_mask  ),      

               // PE 30, Lane 2                 
               .pe30__std__lane2_strm0_ready         ( pe30__std__lane2_strm0_ready      ),      
               .std__pe30__lane2_strm0_cntl          ( std__pe30__lane2_strm0_cntl       ),      
               .std__pe30__lane2_strm0_data          ( std__pe30__lane2_strm0_data       ),      
               .std__pe30__lane2_strm0_data_valid    ( std__pe30__lane2_strm0_data_valid ),      
               .std__pe30__lane2_strm0_data_mask     ( std__pe30__lane2_strm0_data_mask  ),      

               .pe30__std__lane2_strm1_ready         ( pe30__std__lane2_strm1_ready      ),      
               .std__pe30__lane2_strm1_cntl          ( std__pe30__lane2_strm1_cntl       ),      
               .std__pe30__lane2_strm1_data          ( std__pe30__lane2_strm1_data       ),      
               .std__pe30__lane2_strm1_data_valid    ( std__pe30__lane2_strm1_data_valid ),      
               .std__pe30__lane2_strm1_data_mask     ( std__pe30__lane2_strm1_data_mask  ),      

               // PE 30, Lane 3                 
               .pe30__std__lane3_strm0_ready         ( pe30__std__lane3_strm0_ready      ),      
               .std__pe30__lane3_strm0_cntl          ( std__pe30__lane3_strm0_cntl       ),      
               .std__pe30__lane3_strm0_data          ( std__pe30__lane3_strm0_data       ),      
               .std__pe30__lane3_strm0_data_valid    ( std__pe30__lane3_strm0_data_valid ),      
               .std__pe30__lane3_strm0_data_mask     ( std__pe30__lane3_strm0_data_mask  ),      

               .pe30__std__lane3_strm1_ready         ( pe30__std__lane3_strm1_ready      ),      
               .std__pe30__lane3_strm1_cntl          ( std__pe30__lane3_strm1_cntl       ),      
               .std__pe30__lane3_strm1_data          ( std__pe30__lane3_strm1_data       ),      
               .std__pe30__lane3_strm1_data_valid    ( std__pe30__lane3_strm1_data_valid ),      
               .std__pe30__lane3_strm1_data_mask     ( std__pe30__lane3_strm1_data_mask  ),      

               // PE 30, Lane 4                 
               .pe30__std__lane4_strm0_ready         ( pe30__std__lane4_strm0_ready      ),      
               .std__pe30__lane4_strm0_cntl          ( std__pe30__lane4_strm0_cntl       ),      
               .std__pe30__lane4_strm0_data          ( std__pe30__lane4_strm0_data       ),      
               .std__pe30__lane4_strm0_data_valid    ( std__pe30__lane4_strm0_data_valid ),      
               .std__pe30__lane4_strm0_data_mask     ( std__pe30__lane4_strm0_data_mask  ),      

               .pe30__std__lane4_strm1_ready         ( pe30__std__lane4_strm1_ready      ),      
               .std__pe30__lane4_strm1_cntl          ( std__pe30__lane4_strm1_cntl       ),      
               .std__pe30__lane4_strm1_data          ( std__pe30__lane4_strm1_data       ),      
               .std__pe30__lane4_strm1_data_valid    ( std__pe30__lane4_strm1_data_valid ),      
               .std__pe30__lane4_strm1_data_mask     ( std__pe30__lane4_strm1_data_mask  ),      

               // PE 30, Lane 5                 
               .pe30__std__lane5_strm0_ready         ( pe30__std__lane5_strm0_ready      ),      
               .std__pe30__lane5_strm0_cntl          ( std__pe30__lane5_strm0_cntl       ),      
               .std__pe30__lane5_strm0_data          ( std__pe30__lane5_strm0_data       ),      
               .std__pe30__lane5_strm0_data_valid    ( std__pe30__lane5_strm0_data_valid ),      
               .std__pe30__lane5_strm0_data_mask     ( std__pe30__lane5_strm0_data_mask  ),      

               .pe30__std__lane5_strm1_ready         ( pe30__std__lane5_strm1_ready      ),      
               .std__pe30__lane5_strm1_cntl          ( std__pe30__lane5_strm1_cntl       ),      
               .std__pe30__lane5_strm1_data          ( std__pe30__lane5_strm1_data       ),      
               .std__pe30__lane5_strm1_data_valid    ( std__pe30__lane5_strm1_data_valid ),      
               .std__pe30__lane5_strm1_data_mask     ( std__pe30__lane5_strm1_data_mask  ),      

               // PE 30, Lane 6                 
               .pe30__std__lane6_strm0_ready         ( pe30__std__lane6_strm0_ready      ),      
               .std__pe30__lane6_strm0_cntl          ( std__pe30__lane6_strm0_cntl       ),      
               .std__pe30__lane6_strm0_data          ( std__pe30__lane6_strm0_data       ),      
               .std__pe30__lane6_strm0_data_valid    ( std__pe30__lane6_strm0_data_valid ),      
               .std__pe30__lane6_strm0_data_mask     ( std__pe30__lane6_strm0_data_mask  ),      

               .pe30__std__lane6_strm1_ready         ( pe30__std__lane6_strm1_ready      ),      
               .std__pe30__lane6_strm1_cntl          ( std__pe30__lane6_strm1_cntl       ),      
               .std__pe30__lane6_strm1_data          ( std__pe30__lane6_strm1_data       ),      
               .std__pe30__lane6_strm1_data_valid    ( std__pe30__lane6_strm1_data_valid ),      
               .std__pe30__lane6_strm1_data_mask     ( std__pe30__lane6_strm1_data_mask  ),      

               // PE 30, Lane 7                 
               .pe30__std__lane7_strm0_ready         ( pe30__std__lane7_strm0_ready      ),      
               .std__pe30__lane7_strm0_cntl          ( std__pe30__lane7_strm0_cntl       ),      
               .std__pe30__lane7_strm0_data          ( std__pe30__lane7_strm0_data       ),      
               .std__pe30__lane7_strm0_data_valid    ( std__pe30__lane7_strm0_data_valid ),      
               .std__pe30__lane7_strm0_data_mask     ( std__pe30__lane7_strm0_data_mask  ),      

               .pe30__std__lane7_strm1_ready         ( pe30__std__lane7_strm1_ready      ),      
               .std__pe30__lane7_strm1_cntl          ( std__pe30__lane7_strm1_cntl       ),      
               .std__pe30__lane7_strm1_data          ( std__pe30__lane7_strm1_data       ),      
               .std__pe30__lane7_strm1_data_valid    ( std__pe30__lane7_strm1_data_valid ),      
               .std__pe30__lane7_strm1_data_mask     ( std__pe30__lane7_strm1_data_mask  ),      

               // PE 30, Lane 8                 
               .pe30__std__lane8_strm0_ready         ( pe30__std__lane8_strm0_ready      ),      
               .std__pe30__lane8_strm0_cntl          ( std__pe30__lane8_strm0_cntl       ),      
               .std__pe30__lane8_strm0_data          ( std__pe30__lane8_strm0_data       ),      
               .std__pe30__lane8_strm0_data_valid    ( std__pe30__lane8_strm0_data_valid ),      
               .std__pe30__lane8_strm0_data_mask     ( std__pe30__lane8_strm0_data_mask  ),      

               .pe30__std__lane8_strm1_ready         ( pe30__std__lane8_strm1_ready      ),      
               .std__pe30__lane8_strm1_cntl          ( std__pe30__lane8_strm1_cntl       ),      
               .std__pe30__lane8_strm1_data          ( std__pe30__lane8_strm1_data       ),      
               .std__pe30__lane8_strm1_data_valid    ( std__pe30__lane8_strm1_data_valid ),      
               .std__pe30__lane8_strm1_data_mask     ( std__pe30__lane8_strm1_data_mask  ),      

               // PE 30, Lane 9                 
               .pe30__std__lane9_strm0_ready         ( pe30__std__lane9_strm0_ready      ),      
               .std__pe30__lane9_strm0_cntl          ( std__pe30__lane9_strm0_cntl       ),      
               .std__pe30__lane9_strm0_data          ( std__pe30__lane9_strm0_data       ),      
               .std__pe30__lane9_strm0_data_valid    ( std__pe30__lane9_strm0_data_valid ),      
               .std__pe30__lane9_strm0_data_mask     ( std__pe30__lane9_strm0_data_mask  ),      

               .pe30__std__lane9_strm1_ready         ( pe30__std__lane9_strm1_ready      ),      
               .std__pe30__lane9_strm1_cntl          ( std__pe30__lane9_strm1_cntl       ),      
               .std__pe30__lane9_strm1_data          ( std__pe30__lane9_strm1_data       ),      
               .std__pe30__lane9_strm1_data_valid    ( std__pe30__lane9_strm1_data_valid ),      
               .std__pe30__lane9_strm1_data_mask     ( std__pe30__lane9_strm1_data_mask  ),      

               // PE 30, Lane 10                 
               .pe30__std__lane10_strm0_ready         ( pe30__std__lane10_strm0_ready      ),      
               .std__pe30__lane10_strm0_cntl          ( std__pe30__lane10_strm0_cntl       ),      
               .std__pe30__lane10_strm0_data          ( std__pe30__lane10_strm0_data       ),      
               .std__pe30__lane10_strm0_data_valid    ( std__pe30__lane10_strm0_data_valid ),      
               .std__pe30__lane10_strm0_data_mask     ( std__pe30__lane10_strm0_data_mask  ),      

               .pe30__std__lane10_strm1_ready         ( pe30__std__lane10_strm1_ready      ),      
               .std__pe30__lane10_strm1_cntl          ( std__pe30__lane10_strm1_cntl       ),      
               .std__pe30__lane10_strm1_data          ( std__pe30__lane10_strm1_data       ),      
               .std__pe30__lane10_strm1_data_valid    ( std__pe30__lane10_strm1_data_valid ),      
               .std__pe30__lane10_strm1_data_mask     ( std__pe30__lane10_strm1_data_mask  ),      

               // PE 30, Lane 11                 
               .pe30__std__lane11_strm0_ready         ( pe30__std__lane11_strm0_ready      ),      
               .std__pe30__lane11_strm0_cntl          ( std__pe30__lane11_strm0_cntl       ),      
               .std__pe30__lane11_strm0_data          ( std__pe30__lane11_strm0_data       ),      
               .std__pe30__lane11_strm0_data_valid    ( std__pe30__lane11_strm0_data_valid ),      
               .std__pe30__lane11_strm0_data_mask     ( std__pe30__lane11_strm0_data_mask  ),      

               .pe30__std__lane11_strm1_ready         ( pe30__std__lane11_strm1_ready      ),      
               .std__pe30__lane11_strm1_cntl          ( std__pe30__lane11_strm1_cntl       ),      
               .std__pe30__lane11_strm1_data          ( std__pe30__lane11_strm1_data       ),      
               .std__pe30__lane11_strm1_data_valid    ( std__pe30__lane11_strm1_data_valid ),      
               .std__pe30__lane11_strm1_data_mask     ( std__pe30__lane11_strm1_data_mask  ),      

               // PE 30, Lane 12                 
               .pe30__std__lane12_strm0_ready         ( pe30__std__lane12_strm0_ready      ),      
               .std__pe30__lane12_strm0_cntl          ( std__pe30__lane12_strm0_cntl       ),      
               .std__pe30__lane12_strm0_data          ( std__pe30__lane12_strm0_data       ),      
               .std__pe30__lane12_strm0_data_valid    ( std__pe30__lane12_strm0_data_valid ),      
               .std__pe30__lane12_strm0_data_mask     ( std__pe30__lane12_strm0_data_mask  ),      

               .pe30__std__lane12_strm1_ready         ( pe30__std__lane12_strm1_ready      ),      
               .std__pe30__lane12_strm1_cntl          ( std__pe30__lane12_strm1_cntl       ),      
               .std__pe30__lane12_strm1_data          ( std__pe30__lane12_strm1_data       ),      
               .std__pe30__lane12_strm1_data_valid    ( std__pe30__lane12_strm1_data_valid ),      
               .std__pe30__lane12_strm1_data_mask     ( std__pe30__lane12_strm1_data_mask  ),      

               // PE 30, Lane 13                 
               .pe30__std__lane13_strm0_ready         ( pe30__std__lane13_strm0_ready      ),      
               .std__pe30__lane13_strm0_cntl          ( std__pe30__lane13_strm0_cntl       ),      
               .std__pe30__lane13_strm0_data          ( std__pe30__lane13_strm0_data       ),      
               .std__pe30__lane13_strm0_data_valid    ( std__pe30__lane13_strm0_data_valid ),      
               .std__pe30__lane13_strm0_data_mask     ( std__pe30__lane13_strm0_data_mask  ),      

               .pe30__std__lane13_strm1_ready         ( pe30__std__lane13_strm1_ready      ),      
               .std__pe30__lane13_strm1_cntl          ( std__pe30__lane13_strm1_cntl       ),      
               .std__pe30__lane13_strm1_data          ( std__pe30__lane13_strm1_data       ),      
               .std__pe30__lane13_strm1_data_valid    ( std__pe30__lane13_strm1_data_valid ),      
               .std__pe30__lane13_strm1_data_mask     ( std__pe30__lane13_strm1_data_mask  ),      

               // PE 30, Lane 14                 
               .pe30__std__lane14_strm0_ready         ( pe30__std__lane14_strm0_ready      ),      
               .std__pe30__lane14_strm0_cntl          ( std__pe30__lane14_strm0_cntl       ),      
               .std__pe30__lane14_strm0_data          ( std__pe30__lane14_strm0_data       ),      
               .std__pe30__lane14_strm0_data_valid    ( std__pe30__lane14_strm0_data_valid ),      
               .std__pe30__lane14_strm0_data_mask     ( std__pe30__lane14_strm0_data_mask  ),      

               .pe30__std__lane14_strm1_ready         ( pe30__std__lane14_strm1_ready      ),      
               .std__pe30__lane14_strm1_cntl          ( std__pe30__lane14_strm1_cntl       ),      
               .std__pe30__lane14_strm1_data          ( std__pe30__lane14_strm1_data       ),      
               .std__pe30__lane14_strm1_data_valid    ( std__pe30__lane14_strm1_data_valid ),      
               .std__pe30__lane14_strm1_data_mask     ( std__pe30__lane14_strm1_data_mask  ),      

               // PE 30, Lane 15                 
               .pe30__std__lane15_strm0_ready         ( pe30__std__lane15_strm0_ready      ),      
               .std__pe30__lane15_strm0_cntl          ( std__pe30__lane15_strm0_cntl       ),      
               .std__pe30__lane15_strm0_data          ( std__pe30__lane15_strm0_data       ),      
               .std__pe30__lane15_strm0_data_valid    ( std__pe30__lane15_strm0_data_valid ),      
               .std__pe30__lane15_strm0_data_mask     ( std__pe30__lane15_strm0_data_mask  ),      

               .pe30__std__lane15_strm1_ready         ( pe30__std__lane15_strm1_ready      ),      
               .std__pe30__lane15_strm1_cntl          ( std__pe30__lane15_strm1_cntl       ),      
               .std__pe30__lane15_strm1_data          ( std__pe30__lane15_strm1_data       ),      
               .std__pe30__lane15_strm1_data_valid    ( std__pe30__lane15_strm1_data_valid ),      
               .std__pe30__lane15_strm1_data_mask     ( std__pe30__lane15_strm1_data_mask  ),      

               // PE 30, Lane 16                 
               .pe30__std__lane16_strm0_ready         ( pe30__std__lane16_strm0_ready      ),      
               .std__pe30__lane16_strm0_cntl          ( std__pe30__lane16_strm0_cntl       ),      
               .std__pe30__lane16_strm0_data          ( std__pe30__lane16_strm0_data       ),      
               .std__pe30__lane16_strm0_data_valid    ( std__pe30__lane16_strm0_data_valid ),      
               .std__pe30__lane16_strm0_data_mask     ( std__pe30__lane16_strm0_data_mask  ),      

               .pe30__std__lane16_strm1_ready         ( pe30__std__lane16_strm1_ready      ),      
               .std__pe30__lane16_strm1_cntl          ( std__pe30__lane16_strm1_cntl       ),      
               .std__pe30__lane16_strm1_data          ( std__pe30__lane16_strm1_data       ),      
               .std__pe30__lane16_strm1_data_valid    ( std__pe30__lane16_strm1_data_valid ),      
               .std__pe30__lane16_strm1_data_mask     ( std__pe30__lane16_strm1_data_mask  ),      

               // PE 30, Lane 17                 
               .pe30__std__lane17_strm0_ready         ( pe30__std__lane17_strm0_ready      ),      
               .std__pe30__lane17_strm0_cntl          ( std__pe30__lane17_strm0_cntl       ),      
               .std__pe30__lane17_strm0_data          ( std__pe30__lane17_strm0_data       ),      
               .std__pe30__lane17_strm0_data_valid    ( std__pe30__lane17_strm0_data_valid ),      
               .std__pe30__lane17_strm0_data_mask     ( std__pe30__lane17_strm0_data_mask  ),      

               .pe30__std__lane17_strm1_ready         ( pe30__std__lane17_strm1_ready      ),      
               .std__pe30__lane17_strm1_cntl          ( std__pe30__lane17_strm1_cntl       ),      
               .std__pe30__lane17_strm1_data          ( std__pe30__lane17_strm1_data       ),      
               .std__pe30__lane17_strm1_data_valid    ( std__pe30__lane17_strm1_data_valid ),      
               .std__pe30__lane17_strm1_data_mask     ( std__pe30__lane17_strm1_data_mask  ),      

               // PE 30, Lane 18                 
               .pe30__std__lane18_strm0_ready         ( pe30__std__lane18_strm0_ready      ),      
               .std__pe30__lane18_strm0_cntl          ( std__pe30__lane18_strm0_cntl       ),      
               .std__pe30__lane18_strm0_data          ( std__pe30__lane18_strm0_data       ),      
               .std__pe30__lane18_strm0_data_valid    ( std__pe30__lane18_strm0_data_valid ),      
               .std__pe30__lane18_strm0_data_mask     ( std__pe30__lane18_strm0_data_mask  ),      

               .pe30__std__lane18_strm1_ready         ( pe30__std__lane18_strm1_ready      ),      
               .std__pe30__lane18_strm1_cntl          ( std__pe30__lane18_strm1_cntl       ),      
               .std__pe30__lane18_strm1_data          ( std__pe30__lane18_strm1_data       ),      
               .std__pe30__lane18_strm1_data_valid    ( std__pe30__lane18_strm1_data_valid ),      
               .std__pe30__lane18_strm1_data_mask     ( std__pe30__lane18_strm1_data_mask  ),      

               // PE 30, Lane 19                 
               .pe30__std__lane19_strm0_ready         ( pe30__std__lane19_strm0_ready      ),      
               .std__pe30__lane19_strm0_cntl          ( std__pe30__lane19_strm0_cntl       ),      
               .std__pe30__lane19_strm0_data          ( std__pe30__lane19_strm0_data       ),      
               .std__pe30__lane19_strm0_data_valid    ( std__pe30__lane19_strm0_data_valid ),      
               .std__pe30__lane19_strm0_data_mask     ( std__pe30__lane19_strm0_data_mask  ),      

               .pe30__std__lane19_strm1_ready         ( pe30__std__lane19_strm1_ready      ),      
               .std__pe30__lane19_strm1_cntl          ( std__pe30__lane19_strm1_cntl       ),      
               .std__pe30__lane19_strm1_data          ( std__pe30__lane19_strm1_data       ),      
               .std__pe30__lane19_strm1_data_valid    ( std__pe30__lane19_strm1_data_valid ),      
               .std__pe30__lane19_strm1_data_mask     ( std__pe30__lane19_strm1_data_mask  ),      

               // PE 30, Lane 20                 
               .pe30__std__lane20_strm0_ready         ( pe30__std__lane20_strm0_ready      ),      
               .std__pe30__lane20_strm0_cntl          ( std__pe30__lane20_strm0_cntl       ),      
               .std__pe30__lane20_strm0_data          ( std__pe30__lane20_strm0_data       ),      
               .std__pe30__lane20_strm0_data_valid    ( std__pe30__lane20_strm0_data_valid ),      
               .std__pe30__lane20_strm0_data_mask     ( std__pe30__lane20_strm0_data_mask  ),      

               .pe30__std__lane20_strm1_ready         ( pe30__std__lane20_strm1_ready      ),      
               .std__pe30__lane20_strm1_cntl          ( std__pe30__lane20_strm1_cntl       ),      
               .std__pe30__lane20_strm1_data          ( std__pe30__lane20_strm1_data       ),      
               .std__pe30__lane20_strm1_data_valid    ( std__pe30__lane20_strm1_data_valid ),      
               .std__pe30__lane20_strm1_data_mask     ( std__pe30__lane20_strm1_data_mask  ),      

               // PE 30, Lane 21                 
               .pe30__std__lane21_strm0_ready         ( pe30__std__lane21_strm0_ready      ),      
               .std__pe30__lane21_strm0_cntl          ( std__pe30__lane21_strm0_cntl       ),      
               .std__pe30__lane21_strm0_data          ( std__pe30__lane21_strm0_data       ),      
               .std__pe30__lane21_strm0_data_valid    ( std__pe30__lane21_strm0_data_valid ),      
               .std__pe30__lane21_strm0_data_mask     ( std__pe30__lane21_strm0_data_mask  ),      

               .pe30__std__lane21_strm1_ready         ( pe30__std__lane21_strm1_ready      ),      
               .std__pe30__lane21_strm1_cntl          ( std__pe30__lane21_strm1_cntl       ),      
               .std__pe30__lane21_strm1_data          ( std__pe30__lane21_strm1_data       ),      
               .std__pe30__lane21_strm1_data_valid    ( std__pe30__lane21_strm1_data_valid ),      
               .std__pe30__lane21_strm1_data_mask     ( std__pe30__lane21_strm1_data_mask  ),      

               // PE 30, Lane 22                 
               .pe30__std__lane22_strm0_ready         ( pe30__std__lane22_strm0_ready      ),      
               .std__pe30__lane22_strm0_cntl          ( std__pe30__lane22_strm0_cntl       ),      
               .std__pe30__lane22_strm0_data          ( std__pe30__lane22_strm0_data       ),      
               .std__pe30__lane22_strm0_data_valid    ( std__pe30__lane22_strm0_data_valid ),      
               .std__pe30__lane22_strm0_data_mask     ( std__pe30__lane22_strm0_data_mask  ),      

               .pe30__std__lane22_strm1_ready         ( pe30__std__lane22_strm1_ready      ),      
               .std__pe30__lane22_strm1_cntl          ( std__pe30__lane22_strm1_cntl       ),      
               .std__pe30__lane22_strm1_data          ( std__pe30__lane22_strm1_data       ),      
               .std__pe30__lane22_strm1_data_valid    ( std__pe30__lane22_strm1_data_valid ),      
               .std__pe30__lane22_strm1_data_mask     ( std__pe30__lane22_strm1_data_mask  ),      

               // PE 30, Lane 23                 
               .pe30__std__lane23_strm0_ready         ( pe30__std__lane23_strm0_ready      ),      
               .std__pe30__lane23_strm0_cntl          ( std__pe30__lane23_strm0_cntl       ),      
               .std__pe30__lane23_strm0_data          ( std__pe30__lane23_strm0_data       ),      
               .std__pe30__lane23_strm0_data_valid    ( std__pe30__lane23_strm0_data_valid ),      
               .std__pe30__lane23_strm0_data_mask     ( std__pe30__lane23_strm0_data_mask  ),      

               .pe30__std__lane23_strm1_ready         ( pe30__std__lane23_strm1_ready      ),      
               .std__pe30__lane23_strm1_cntl          ( std__pe30__lane23_strm1_cntl       ),      
               .std__pe30__lane23_strm1_data          ( std__pe30__lane23_strm1_data       ),      
               .std__pe30__lane23_strm1_data_valid    ( std__pe30__lane23_strm1_data_valid ),      
               .std__pe30__lane23_strm1_data_mask     ( std__pe30__lane23_strm1_data_mask  ),      

               // PE 30, Lane 24                 
               .pe30__std__lane24_strm0_ready         ( pe30__std__lane24_strm0_ready      ),      
               .std__pe30__lane24_strm0_cntl          ( std__pe30__lane24_strm0_cntl       ),      
               .std__pe30__lane24_strm0_data          ( std__pe30__lane24_strm0_data       ),      
               .std__pe30__lane24_strm0_data_valid    ( std__pe30__lane24_strm0_data_valid ),      
               .std__pe30__lane24_strm0_data_mask     ( std__pe30__lane24_strm0_data_mask  ),      

               .pe30__std__lane24_strm1_ready         ( pe30__std__lane24_strm1_ready      ),      
               .std__pe30__lane24_strm1_cntl          ( std__pe30__lane24_strm1_cntl       ),      
               .std__pe30__lane24_strm1_data          ( std__pe30__lane24_strm1_data       ),      
               .std__pe30__lane24_strm1_data_valid    ( std__pe30__lane24_strm1_data_valid ),      
               .std__pe30__lane24_strm1_data_mask     ( std__pe30__lane24_strm1_data_mask  ),      

               // PE 30, Lane 25                 
               .pe30__std__lane25_strm0_ready         ( pe30__std__lane25_strm0_ready      ),      
               .std__pe30__lane25_strm0_cntl          ( std__pe30__lane25_strm0_cntl       ),      
               .std__pe30__lane25_strm0_data          ( std__pe30__lane25_strm0_data       ),      
               .std__pe30__lane25_strm0_data_valid    ( std__pe30__lane25_strm0_data_valid ),      
               .std__pe30__lane25_strm0_data_mask     ( std__pe30__lane25_strm0_data_mask  ),      

               .pe30__std__lane25_strm1_ready         ( pe30__std__lane25_strm1_ready      ),      
               .std__pe30__lane25_strm1_cntl          ( std__pe30__lane25_strm1_cntl       ),      
               .std__pe30__lane25_strm1_data          ( std__pe30__lane25_strm1_data       ),      
               .std__pe30__lane25_strm1_data_valid    ( std__pe30__lane25_strm1_data_valid ),      
               .std__pe30__lane25_strm1_data_mask     ( std__pe30__lane25_strm1_data_mask  ),      

               // PE 30, Lane 26                 
               .pe30__std__lane26_strm0_ready         ( pe30__std__lane26_strm0_ready      ),      
               .std__pe30__lane26_strm0_cntl          ( std__pe30__lane26_strm0_cntl       ),      
               .std__pe30__lane26_strm0_data          ( std__pe30__lane26_strm0_data       ),      
               .std__pe30__lane26_strm0_data_valid    ( std__pe30__lane26_strm0_data_valid ),      
               .std__pe30__lane26_strm0_data_mask     ( std__pe30__lane26_strm0_data_mask  ),      

               .pe30__std__lane26_strm1_ready         ( pe30__std__lane26_strm1_ready      ),      
               .std__pe30__lane26_strm1_cntl          ( std__pe30__lane26_strm1_cntl       ),      
               .std__pe30__lane26_strm1_data          ( std__pe30__lane26_strm1_data       ),      
               .std__pe30__lane26_strm1_data_valid    ( std__pe30__lane26_strm1_data_valid ),      
               .std__pe30__lane26_strm1_data_mask     ( std__pe30__lane26_strm1_data_mask  ),      

               // PE 30, Lane 27                 
               .pe30__std__lane27_strm0_ready         ( pe30__std__lane27_strm0_ready      ),      
               .std__pe30__lane27_strm0_cntl          ( std__pe30__lane27_strm0_cntl       ),      
               .std__pe30__lane27_strm0_data          ( std__pe30__lane27_strm0_data       ),      
               .std__pe30__lane27_strm0_data_valid    ( std__pe30__lane27_strm0_data_valid ),      
               .std__pe30__lane27_strm0_data_mask     ( std__pe30__lane27_strm0_data_mask  ),      

               .pe30__std__lane27_strm1_ready         ( pe30__std__lane27_strm1_ready      ),      
               .std__pe30__lane27_strm1_cntl          ( std__pe30__lane27_strm1_cntl       ),      
               .std__pe30__lane27_strm1_data          ( std__pe30__lane27_strm1_data       ),      
               .std__pe30__lane27_strm1_data_valid    ( std__pe30__lane27_strm1_data_valid ),      
               .std__pe30__lane27_strm1_data_mask     ( std__pe30__lane27_strm1_data_mask  ),      

               // PE 30, Lane 28                 
               .pe30__std__lane28_strm0_ready         ( pe30__std__lane28_strm0_ready      ),      
               .std__pe30__lane28_strm0_cntl          ( std__pe30__lane28_strm0_cntl       ),      
               .std__pe30__lane28_strm0_data          ( std__pe30__lane28_strm0_data       ),      
               .std__pe30__lane28_strm0_data_valid    ( std__pe30__lane28_strm0_data_valid ),      
               .std__pe30__lane28_strm0_data_mask     ( std__pe30__lane28_strm0_data_mask  ),      

               .pe30__std__lane28_strm1_ready         ( pe30__std__lane28_strm1_ready      ),      
               .std__pe30__lane28_strm1_cntl          ( std__pe30__lane28_strm1_cntl       ),      
               .std__pe30__lane28_strm1_data          ( std__pe30__lane28_strm1_data       ),      
               .std__pe30__lane28_strm1_data_valid    ( std__pe30__lane28_strm1_data_valid ),      
               .std__pe30__lane28_strm1_data_mask     ( std__pe30__lane28_strm1_data_mask  ),      

               // PE 30, Lane 29                 
               .pe30__std__lane29_strm0_ready         ( pe30__std__lane29_strm0_ready      ),      
               .std__pe30__lane29_strm0_cntl          ( std__pe30__lane29_strm0_cntl       ),      
               .std__pe30__lane29_strm0_data          ( std__pe30__lane29_strm0_data       ),      
               .std__pe30__lane29_strm0_data_valid    ( std__pe30__lane29_strm0_data_valid ),      
               .std__pe30__lane29_strm0_data_mask     ( std__pe30__lane29_strm0_data_mask  ),      

               .pe30__std__lane29_strm1_ready         ( pe30__std__lane29_strm1_ready      ),      
               .std__pe30__lane29_strm1_cntl          ( std__pe30__lane29_strm1_cntl       ),      
               .std__pe30__lane29_strm1_data          ( std__pe30__lane29_strm1_data       ),      
               .std__pe30__lane29_strm1_data_valid    ( std__pe30__lane29_strm1_data_valid ),      
               .std__pe30__lane29_strm1_data_mask     ( std__pe30__lane29_strm1_data_mask  ),      

               // PE 30, Lane 30                 
               .pe30__std__lane30_strm0_ready         ( pe30__std__lane30_strm0_ready      ),      
               .std__pe30__lane30_strm0_cntl          ( std__pe30__lane30_strm0_cntl       ),      
               .std__pe30__lane30_strm0_data          ( std__pe30__lane30_strm0_data       ),      
               .std__pe30__lane30_strm0_data_valid    ( std__pe30__lane30_strm0_data_valid ),      
               .std__pe30__lane30_strm0_data_mask     ( std__pe30__lane30_strm0_data_mask  ),      

               .pe30__std__lane30_strm1_ready         ( pe30__std__lane30_strm1_ready      ),      
               .std__pe30__lane30_strm1_cntl          ( std__pe30__lane30_strm1_cntl       ),      
               .std__pe30__lane30_strm1_data          ( std__pe30__lane30_strm1_data       ),      
               .std__pe30__lane30_strm1_data_valid    ( std__pe30__lane30_strm1_data_valid ),      
               .std__pe30__lane30_strm1_data_mask     ( std__pe30__lane30_strm1_data_mask  ),      

               // PE 30, Lane 31                 
               .pe30__std__lane31_strm0_ready         ( pe30__std__lane31_strm0_ready      ),      
               .std__pe30__lane31_strm0_cntl          ( std__pe30__lane31_strm0_cntl       ),      
               .std__pe30__lane31_strm0_data          ( std__pe30__lane31_strm0_data       ),      
               .std__pe30__lane31_strm0_data_valid    ( std__pe30__lane31_strm0_data_valid ),      
               .std__pe30__lane31_strm0_data_mask     ( std__pe30__lane31_strm0_data_mask  ),      

               .pe30__std__lane31_strm1_ready         ( pe30__std__lane31_strm1_ready      ),      
               .std__pe30__lane31_strm1_cntl          ( std__pe30__lane31_strm1_cntl       ),      
               .std__pe30__lane31_strm1_data          ( std__pe30__lane31_strm1_data       ),      
               .std__pe30__lane31_strm1_data_valid    ( std__pe30__lane31_strm1_data_valid ),      
               .std__pe30__lane31_strm1_data_mask     ( std__pe30__lane31_strm1_data_mask  ),      

               // PE 31, Lane 0                 
               .pe31__std__lane0_strm0_ready         ( pe31__std__lane0_strm0_ready      ),      
               .std__pe31__lane0_strm0_cntl          ( std__pe31__lane0_strm0_cntl       ),      
               .std__pe31__lane0_strm0_data          ( std__pe31__lane0_strm0_data       ),      
               .std__pe31__lane0_strm0_data_valid    ( std__pe31__lane0_strm0_data_valid ),      
               .std__pe31__lane0_strm0_data_mask     ( std__pe31__lane0_strm0_data_mask  ),      

               .pe31__std__lane0_strm1_ready         ( pe31__std__lane0_strm1_ready      ),      
               .std__pe31__lane0_strm1_cntl          ( std__pe31__lane0_strm1_cntl       ),      
               .std__pe31__lane0_strm1_data          ( std__pe31__lane0_strm1_data       ),      
               .std__pe31__lane0_strm1_data_valid    ( std__pe31__lane0_strm1_data_valid ),      
               .std__pe31__lane0_strm1_data_mask     ( std__pe31__lane0_strm1_data_mask  ),      

               // PE 31, Lane 1                 
               .pe31__std__lane1_strm0_ready         ( pe31__std__lane1_strm0_ready      ),      
               .std__pe31__lane1_strm0_cntl          ( std__pe31__lane1_strm0_cntl       ),      
               .std__pe31__lane1_strm0_data          ( std__pe31__lane1_strm0_data       ),      
               .std__pe31__lane1_strm0_data_valid    ( std__pe31__lane1_strm0_data_valid ),      
               .std__pe31__lane1_strm0_data_mask     ( std__pe31__lane1_strm0_data_mask  ),      

               .pe31__std__lane1_strm1_ready         ( pe31__std__lane1_strm1_ready      ),      
               .std__pe31__lane1_strm1_cntl          ( std__pe31__lane1_strm1_cntl       ),      
               .std__pe31__lane1_strm1_data          ( std__pe31__lane1_strm1_data       ),      
               .std__pe31__lane1_strm1_data_valid    ( std__pe31__lane1_strm1_data_valid ),      
               .std__pe31__lane1_strm1_data_mask     ( std__pe31__lane1_strm1_data_mask  ),      

               // PE 31, Lane 2                 
               .pe31__std__lane2_strm0_ready         ( pe31__std__lane2_strm0_ready      ),      
               .std__pe31__lane2_strm0_cntl          ( std__pe31__lane2_strm0_cntl       ),      
               .std__pe31__lane2_strm0_data          ( std__pe31__lane2_strm0_data       ),      
               .std__pe31__lane2_strm0_data_valid    ( std__pe31__lane2_strm0_data_valid ),      
               .std__pe31__lane2_strm0_data_mask     ( std__pe31__lane2_strm0_data_mask  ),      

               .pe31__std__lane2_strm1_ready         ( pe31__std__lane2_strm1_ready      ),      
               .std__pe31__lane2_strm1_cntl          ( std__pe31__lane2_strm1_cntl       ),      
               .std__pe31__lane2_strm1_data          ( std__pe31__lane2_strm1_data       ),      
               .std__pe31__lane2_strm1_data_valid    ( std__pe31__lane2_strm1_data_valid ),      
               .std__pe31__lane2_strm1_data_mask     ( std__pe31__lane2_strm1_data_mask  ),      

               // PE 31, Lane 3                 
               .pe31__std__lane3_strm0_ready         ( pe31__std__lane3_strm0_ready      ),      
               .std__pe31__lane3_strm0_cntl          ( std__pe31__lane3_strm0_cntl       ),      
               .std__pe31__lane3_strm0_data          ( std__pe31__lane3_strm0_data       ),      
               .std__pe31__lane3_strm0_data_valid    ( std__pe31__lane3_strm0_data_valid ),      
               .std__pe31__lane3_strm0_data_mask     ( std__pe31__lane3_strm0_data_mask  ),      

               .pe31__std__lane3_strm1_ready         ( pe31__std__lane3_strm1_ready      ),      
               .std__pe31__lane3_strm1_cntl          ( std__pe31__lane3_strm1_cntl       ),      
               .std__pe31__lane3_strm1_data          ( std__pe31__lane3_strm1_data       ),      
               .std__pe31__lane3_strm1_data_valid    ( std__pe31__lane3_strm1_data_valid ),      
               .std__pe31__lane3_strm1_data_mask     ( std__pe31__lane3_strm1_data_mask  ),      

               // PE 31, Lane 4                 
               .pe31__std__lane4_strm0_ready         ( pe31__std__lane4_strm0_ready      ),      
               .std__pe31__lane4_strm0_cntl          ( std__pe31__lane4_strm0_cntl       ),      
               .std__pe31__lane4_strm0_data          ( std__pe31__lane4_strm0_data       ),      
               .std__pe31__lane4_strm0_data_valid    ( std__pe31__lane4_strm0_data_valid ),      
               .std__pe31__lane4_strm0_data_mask     ( std__pe31__lane4_strm0_data_mask  ),      

               .pe31__std__lane4_strm1_ready         ( pe31__std__lane4_strm1_ready      ),      
               .std__pe31__lane4_strm1_cntl          ( std__pe31__lane4_strm1_cntl       ),      
               .std__pe31__lane4_strm1_data          ( std__pe31__lane4_strm1_data       ),      
               .std__pe31__lane4_strm1_data_valid    ( std__pe31__lane4_strm1_data_valid ),      
               .std__pe31__lane4_strm1_data_mask     ( std__pe31__lane4_strm1_data_mask  ),      

               // PE 31, Lane 5                 
               .pe31__std__lane5_strm0_ready         ( pe31__std__lane5_strm0_ready      ),      
               .std__pe31__lane5_strm0_cntl          ( std__pe31__lane5_strm0_cntl       ),      
               .std__pe31__lane5_strm0_data          ( std__pe31__lane5_strm0_data       ),      
               .std__pe31__lane5_strm0_data_valid    ( std__pe31__lane5_strm0_data_valid ),      
               .std__pe31__lane5_strm0_data_mask     ( std__pe31__lane5_strm0_data_mask  ),      

               .pe31__std__lane5_strm1_ready         ( pe31__std__lane5_strm1_ready      ),      
               .std__pe31__lane5_strm1_cntl          ( std__pe31__lane5_strm1_cntl       ),      
               .std__pe31__lane5_strm1_data          ( std__pe31__lane5_strm1_data       ),      
               .std__pe31__lane5_strm1_data_valid    ( std__pe31__lane5_strm1_data_valid ),      
               .std__pe31__lane5_strm1_data_mask     ( std__pe31__lane5_strm1_data_mask  ),      

               // PE 31, Lane 6                 
               .pe31__std__lane6_strm0_ready         ( pe31__std__lane6_strm0_ready      ),      
               .std__pe31__lane6_strm0_cntl          ( std__pe31__lane6_strm0_cntl       ),      
               .std__pe31__lane6_strm0_data          ( std__pe31__lane6_strm0_data       ),      
               .std__pe31__lane6_strm0_data_valid    ( std__pe31__lane6_strm0_data_valid ),      
               .std__pe31__lane6_strm0_data_mask     ( std__pe31__lane6_strm0_data_mask  ),      

               .pe31__std__lane6_strm1_ready         ( pe31__std__lane6_strm1_ready      ),      
               .std__pe31__lane6_strm1_cntl          ( std__pe31__lane6_strm1_cntl       ),      
               .std__pe31__lane6_strm1_data          ( std__pe31__lane6_strm1_data       ),      
               .std__pe31__lane6_strm1_data_valid    ( std__pe31__lane6_strm1_data_valid ),      
               .std__pe31__lane6_strm1_data_mask     ( std__pe31__lane6_strm1_data_mask  ),      

               // PE 31, Lane 7                 
               .pe31__std__lane7_strm0_ready         ( pe31__std__lane7_strm0_ready      ),      
               .std__pe31__lane7_strm0_cntl          ( std__pe31__lane7_strm0_cntl       ),      
               .std__pe31__lane7_strm0_data          ( std__pe31__lane7_strm0_data       ),      
               .std__pe31__lane7_strm0_data_valid    ( std__pe31__lane7_strm0_data_valid ),      
               .std__pe31__lane7_strm0_data_mask     ( std__pe31__lane7_strm0_data_mask  ),      

               .pe31__std__lane7_strm1_ready         ( pe31__std__lane7_strm1_ready      ),      
               .std__pe31__lane7_strm1_cntl          ( std__pe31__lane7_strm1_cntl       ),      
               .std__pe31__lane7_strm1_data          ( std__pe31__lane7_strm1_data       ),      
               .std__pe31__lane7_strm1_data_valid    ( std__pe31__lane7_strm1_data_valid ),      
               .std__pe31__lane7_strm1_data_mask     ( std__pe31__lane7_strm1_data_mask  ),      

               // PE 31, Lane 8                 
               .pe31__std__lane8_strm0_ready         ( pe31__std__lane8_strm0_ready      ),      
               .std__pe31__lane8_strm0_cntl          ( std__pe31__lane8_strm0_cntl       ),      
               .std__pe31__lane8_strm0_data          ( std__pe31__lane8_strm0_data       ),      
               .std__pe31__lane8_strm0_data_valid    ( std__pe31__lane8_strm0_data_valid ),      
               .std__pe31__lane8_strm0_data_mask     ( std__pe31__lane8_strm0_data_mask  ),      

               .pe31__std__lane8_strm1_ready         ( pe31__std__lane8_strm1_ready      ),      
               .std__pe31__lane8_strm1_cntl          ( std__pe31__lane8_strm1_cntl       ),      
               .std__pe31__lane8_strm1_data          ( std__pe31__lane8_strm1_data       ),      
               .std__pe31__lane8_strm1_data_valid    ( std__pe31__lane8_strm1_data_valid ),      
               .std__pe31__lane8_strm1_data_mask     ( std__pe31__lane8_strm1_data_mask  ),      

               // PE 31, Lane 9                 
               .pe31__std__lane9_strm0_ready         ( pe31__std__lane9_strm0_ready      ),      
               .std__pe31__lane9_strm0_cntl          ( std__pe31__lane9_strm0_cntl       ),      
               .std__pe31__lane9_strm0_data          ( std__pe31__lane9_strm0_data       ),      
               .std__pe31__lane9_strm0_data_valid    ( std__pe31__lane9_strm0_data_valid ),      
               .std__pe31__lane9_strm0_data_mask     ( std__pe31__lane9_strm0_data_mask  ),      

               .pe31__std__lane9_strm1_ready         ( pe31__std__lane9_strm1_ready      ),      
               .std__pe31__lane9_strm1_cntl          ( std__pe31__lane9_strm1_cntl       ),      
               .std__pe31__lane9_strm1_data          ( std__pe31__lane9_strm1_data       ),      
               .std__pe31__lane9_strm1_data_valid    ( std__pe31__lane9_strm1_data_valid ),      
               .std__pe31__lane9_strm1_data_mask     ( std__pe31__lane9_strm1_data_mask  ),      

               // PE 31, Lane 10                 
               .pe31__std__lane10_strm0_ready         ( pe31__std__lane10_strm0_ready      ),      
               .std__pe31__lane10_strm0_cntl          ( std__pe31__lane10_strm0_cntl       ),      
               .std__pe31__lane10_strm0_data          ( std__pe31__lane10_strm0_data       ),      
               .std__pe31__lane10_strm0_data_valid    ( std__pe31__lane10_strm0_data_valid ),      
               .std__pe31__lane10_strm0_data_mask     ( std__pe31__lane10_strm0_data_mask  ),      

               .pe31__std__lane10_strm1_ready         ( pe31__std__lane10_strm1_ready      ),      
               .std__pe31__lane10_strm1_cntl          ( std__pe31__lane10_strm1_cntl       ),      
               .std__pe31__lane10_strm1_data          ( std__pe31__lane10_strm1_data       ),      
               .std__pe31__lane10_strm1_data_valid    ( std__pe31__lane10_strm1_data_valid ),      
               .std__pe31__lane10_strm1_data_mask     ( std__pe31__lane10_strm1_data_mask  ),      

               // PE 31, Lane 11                 
               .pe31__std__lane11_strm0_ready         ( pe31__std__lane11_strm0_ready      ),      
               .std__pe31__lane11_strm0_cntl          ( std__pe31__lane11_strm0_cntl       ),      
               .std__pe31__lane11_strm0_data          ( std__pe31__lane11_strm0_data       ),      
               .std__pe31__lane11_strm0_data_valid    ( std__pe31__lane11_strm0_data_valid ),      
               .std__pe31__lane11_strm0_data_mask     ( std__pe31__lane11_strm0_data_mask  ),      

               .pe31__std__lane11_strm1_ready         ( pe31__std__lane11_strm1_ready      ),      
               .std__pe31__lane11_strm1_cntl          ( std__pe31__lane11_strm1_cntl       ),      
               .std__pe31__lane11_strm1_data          ( std__pe31__lane11_strm1_data       ),      
               .std__pe31__lane11_strm1_data_valid    ( std__pe31__lane11_strm1_data_valid ),      
               .std__pe31__lane11_strm1_data_mask     ( std__pe31__lane11_strm1_data_mask  ),      

               // PE 31, Lane 12                 
               .pe31__std__lane12_strm0_ready         ( pe31__std__lane12_strm0_ready      ),      
               .std__pe31__lane12_strm0_cntl          ( std__pe31__lane12_strm0_cntl       ),      
               .std__pe31__lane12_strm0_data          ( std__pe31__lane12_strm0_data       ),      
               .std__pe31__lane12_strm0_data_valid    ( std__pe31__lane12_strm0_data_valid ),      
               .std__pe31__lane12_strm0_data_mask     ( std__pe31__lane12_strm0_data_mask  ),      

               .pe31__std__lane12_strm1_ready         ( pe31__std__lane12_strm1_ready      ),      
               .std__pe31__lane12_strm1_cntl          ( std__pe31__lane12_strm1_cntl       ),      
               .std__pe31__lane12_strm1_data          ( std__pe31__lane12_strm1_data       ),      
               .std__pe31__lane12_strm1_data_valid    ( std__pe31__lane12_strm1_data_valid ),      
               .std__pe31__lane12_strm1_data_mask     ( std__pe31__lane12_strm1_data_mask  ),      

               // PE 31, Lane 13                 
               .pe31__std__lane13_strm0_ready         ( pe31__std__lane13_strm0_ready      ),      
               .std__pe31__lane13_strm0_cntl          ( std__pe31__lane13_strm0_cntl       ),      
               .std__pe31__lane13_strm0_data          ( std__pe31__lane13_strm0_data       ),      
               .std__pe31__lane13_strm0_data_valid    ( std__pe31__lane13_strm0_data_valid ),      
               .std__pe31__lane13_strm0_data_mask     ( std__pe31__lane13_strm0_data_mask  ),      

               .pe31__std__lane13_strm1_ready         ( pe31__std__lane13_strm1_ready      ),      
               .std__pe31__lane13_strm1_cntl          ( std__pe31__lane13_strm1_cntl       ),      
               .std__pe31__lane13_strm1_data          ( std__pe31__lane13_strm1_data       ),      
               .std__pe31__lane13_strm1_data_valid    ( std__pe31__lane13_strm1_data_valid ),      
               .std__pe31__lane13_strm1_data_mask     ( std__pe31__lane13_strm1_data_mask  ),      

               // PE 31, Lane 14                 
               .pe31__std__lane14_strm0_ready         ( pe31__std__lane14_strm0_ready      ),      
               .std__pe31__lane14_strm0_cntl          ( std__pe31__lane14_strm0_cntl       ),      
               .std__pe31__lane14_strm0_data          ( std__pe31__lane14_strm0_data       ),      
               .std__pe31__lane14_strm0_data_valid    ( std__pe31__lane14_strm0_data_valid ),      
               .std__pe31__lane14_strm0_data_mask     ( std__pe31__lane14_strm0_data_mask  ),      

               .pe31__std__lane14_strm1_ready         ( pe31__std__lane14_strm1_ready      ),      
               .std__pe31__lane14_strm1_cntl          ( std__pe31__lane14_strm1_cntl       ),      
               .std__pe31__lane14_strm1_data          ( std__pe31__lane14_strm1_data       ),      
               .std__pe31__lane14_strm1_data_valid    ( std__pe31__lane14_strm1_data_valid ),      
               .std__pe31__lane14_strm1_data_mask     ( std__pe31__lane14_strm1_data_mask  ),      

               // PE 31, Lane 15                 
               .pe31__std__lane15_strm0_ready         ( pe31__std__lane15_strm0_ready      ),      
               .std__pe31__lane15_strm0_cntl          ( std__pe31__lane15_strm0_cntl       ),      
               .std__pe31__lane15_strm0_data          ( std__pe31__lane15_strm0_data       ),      
               .std__pe31__lane15_strm0_data_valid    ( std__pe31__lane15_strm0_data_valid ),      
               .std__pe31__lane15_strm0_data_mask     ( std__pe31__lane15_strm0_data_mask  ),      

               .pe31__std__lane15_strm1_ready         ( pe31__std__lane15_strm1_ready      ),      
               .std__pe31__lane15_strm1_cntl          ( std__pe31__lane15_strm1_cntl       ),      
               .std__pe31__lane15_strm1_data          ( std__pe31__lane15_strm1_data       ),      
               .std__pe31__lane15_strm1_data_valid    ( std__pe31__lane15_strm1_data_valid ),      
               .std__pe31__lane15_strm1_data_mask     ( std__pe31__lane15_strm1_data_mask  ),      

               // PE 31, Lane 16                 
               .pe31__std__lane16_strm0_ready         ( pe31__std__lane16_strm0_ready      ),      
               .std__pe31__lane16_strm0_cntl          ( std__pe31__lane16_strm0_cntl       ),      
               .std__pe31__lane16_strm0_data          ( std__pe31__lane16_strm0_data       ),      
               .std__pe31__lane16_strm0_data_valid    ( std__pe31__lane16_strm0_data_valid ),      
               .std__pe31__lane16_strm0_data_mask     ( std__pe31__lane16_strm0_data_mask  ),      

               .pe31__std__lane16_strm1_ready         ( pe31__std__lane16_strm1_ready      ),      
               .std__pe31__lane16_strm1_cntl          ( std__pe31__lane16_strm1_cntl       ),      
               .std__pe31__lane16_strm1_data          ( std__pe31__lane16_strm1_data       ),      
               .std__pe31__lane16_strm1_data_valid    ( std__pe31__lane16_strm1_data_valid ),      
               .std__pe31__lane16_strm1_data_mask     ( std__pe31__lane16_strm1_data_mask  ),      

               // PE 31, Lane 17                 
               .pe31__std__lane17_strm0_ready         ( pe31__std__lane17_strm0_ready      ),      
               .std__pe31__lane17_strm0_cntl          ( std__pe31__lane17_strm0_cntl       ),      
               .std__pe31__lane17_strm0_data          ( std__pe31__lane17_strm0_data       ),      
               .std__pe31__lane17_strm0_data_valid    ( std__pe31__lane17_strm0_data_valid ),      
               .std__pe31__lane17_strm0_data_mask     ( std__pe31__lane17_strm0_data_mask  ),      

               .pe31__std__lane17_strm1_ready         ( pe31__std__lane17_strm1_ready      ),      
               .std__pe31__lane17_strm1_cntl          ( std__pe31__lane17_strm1_cntl       ),      
               .std__pe31__lane17_strm1_data          ( std__pe31__lane17_strm1_data       ),      
               .std__pe31__lane17_strm1_data_valid    ( std__pe31__lane17_strm1_data_valid ),      
               .std__pe31__lane17_strm1_data_mask     ( std__pe31__lane17_strm1_data_mask  ),      

               // PE 31, Lane 18                 
               .pe31__std__lane18_strm0_ready         ( pe31__std__lane18_strm0_ready      ),      
               .std__pe31__lane18_strm0_cntl          ( std__pe31__lane18_strm0_cntl       ),      
               .std__pe31__lane18_strm0_data          ( std__pe31__lane18_strm0_data       ),      
               .std__pe31__lane18_strm0_data_valid    ( std__pe31__lane18_strm0_data_valid ),      
               .std__pe31__lane18_strm0_data_mask     ( std__pe31__lane18_strm0_data_mask  ),      

               .pe31__std__lane18_strm1_ready         ( pe31__std__lane18_strm1_ready      ),      
               .std__pe31__lane18_strm1_cntl          ( std__pe31__lane18_strm1_cntl       ),      
               .std__pe31__lane18_strm1_data          ( std__pe31__lane18_strm1_data       ),      
               .std__pe31__lane18_strm1_data_valid    ( std__pe31__lane18_strm1_data_valid ),      
               .std__pe31__lane18_strm1_data_mask     ( std__pe31__lane18_strm1_data_mask  ),      

               // PE 31, Lane 19                 
               .pe31__std__lane19_strm0_ready         ( pe31__std__lane19_strm0_ready      ),      
               .std__pe31__lane19_strm0_cntl          ( std__pe31__lane19_strm0_cntl       ),      
               .std__pe31__lane19_strm0_data          ( std__pe31__lane19_strm0_data       ),      
               .std__pe31__lane19_strm0_data_valid    ( std__pe31__lane19_strm0_data_valid ),      
               .std__pe31__lane19_strm0_data_mask     ( std__pe31__lane19_strm0_data_mask  ),      

               .pe31__std__lane19_strm1_ready         ( pe31__std__lane19_strm1_ready      ),      
               .std__pe31__lane19_strm1_cntl          ( std__pe31__lane19_strm1_cntl       ),      
               .std__pe31__lane19_strm1_data          ( std__pe31__lane19_strm1_data       ),      
               .std__pe31__lane19_strm1_data_valid    ( std__pe31__lane19_strm1_data_valid ),      
               .std__pe31__lane19_strm1_data_mask     ( std__pe31__lane19_strm1_data_mask  ),      

               // PE 31, Lane 20                 
               .pe31__std__lane20_strm0_ready         ( pe31__std__lane20_strm0_ready      ),      
               .std__pe31__lane20_strm0_cntl          ( std__pe31__lane20_strm0_cntl       ),      
               .std__pe31__lane20_strm0_data          ( std__pe31__lane20_strm0_data       ),      
               .std__pe31__lane20_strm0_data_valid    ( std__pe31__lane20_strm0_data_valid ),      
               .std__pe31__lane20_strm0_data_mask     ( std__pe31__lane20_strm0_data_mask  ),      

               .pe31__std__lane20_strm1_ready         ( pe31__std__lane20_strm1_ready      ),      
               .std__pe31__lane20_strm1_cntl          ( std__pe31__lane20_strm1_cntl       ),      
               .std__pe31__lane20_strm1_data          ( std__pe31__lane20_strm1_data       ),      
               .std__pe31__lane20_strm1_data_valid    ( std__pe31__lane20_strm1_data_valid ),      
               .std__pe31__lane20_strm1_data_mask     ( std__pe31__lane20_strm1_data_mask  ),      

               // PE 31, Lane 21                 
               .pe31__std__lane21_strm0_ready         ( pe31__std__lane21_strm0_ready      ),      
               .std__pe31__lane21_strm0_cntl          ( std__pe31__lane21_strm0_cntl       ),      
               .std__pe31__lane21_strm0_data          ( std__pe31__lane21_strm0_data       ),      
               .std__pe31__lane21_strm0_data_valid    ( std__pe31__lane21_strm0_data_valid ),      
               .std__pe31__lane21_strm0_data_mask     ( std__pe31__lane21_strm0_data_mask  ),      

               .pe31__std__lane21_strm1_ready         ( pe31__std__lane21_strm1_ready      ),      
               .std__pe31__lane21_strm1_cntl          ( std__pe31__lane21_strm1_cntl       ),      
               .std__pe31__lane21_strm1_data          ( std__pe31__lane21_strm1_data       ),      
               .std__pe31__lane21_strm1_data_valid    ( std__pe31__lane21_strm1_data_valid ),      
               .std__pe31__lane21_strm1_data_mask     ( std__pe31__lane21_strm1_data_mask  ),      

               // PE 31, Lane 22                 
               .pe31__std__lane22_strm0_ready         ( pe31__std__lane22_strm0_ready      ),      
               .std__pe31__lane22_strm0_cntl          ( std__pe31__lane22_strm0_cntl       ),      
               .std__pe31__lane22_strm0_data          ( std__pe31__lane22_strm0_data       ),      
               .std__pe31__lane22_strm0_data_valid    ( std__pe31__lane22_strm0_data_valid ),      
               .std__pe31__lane22_strm0_data_mask     ( std__pe31__lane22_strm0_data_mask  ),      

               .pe31__std__lane22_strm1_ready         ( pe31__std__lane22_strm1_ready      ),      
               .std__pe31__lane22_strm1_cntl          ( std__pe31__lane22_strm1_cntl       ),      
               .std__pe31__lane22_strm1_data          ( std__pe31__lane22_strm1_data       ),      
               .std__pe31__lane22_strm1_data_valid    ( std__pe31__lane22_strm1_data_valid ),      
               .std__pe31__lane22_strm1_data_mask     ( std__pe31__lane22_strm1_data_mask  ),      

               // PE 31, Lane 23                 
               .pe31__std__lane23_strm0_ready         ( pe31__std__lane23_strm0_ready      ),      
               .std__pe31__lane23_strm0_cntl          ( std__pe31__lane23_strm0_cntl       ),      
               .std__pe31__lane23_strm0_data          ( std__pe31__lane23_strm0_data       ),      
               .std__pe31__lane23_strm0_data_valid    ( std__pe31__lane23_strm0_data_valid ),      
               .std__pe31__lane23_strm0_data_mask     ( std__pe31__lane23_strm0_data_mask  ),      

               .pe31__std__lane23_strm1_ready         ( pe31__std__lane23_strm1_ready      ),      
               .std__pe31__lane23_strm1_cntl          ( std__pe31__lane23_strm1_cntl       ),      
               .std__pe31__lane23_strm1_data          ( std__pe31__lane23_strm1_data       ),      
               .std__pe31__lane23_strm1_data_valid    ( std__pe31__lane23_strm1_data_valid ),      
               .std__pe31__lane23_strm1_data_mask     ( std__pe31__lane23_strm1_data_mask  ),      

               // PE 31, Lane 24                 
               .pe31__std__lane24_strm0_ready         ( pe31__std__lane24_strm0_ready      ),      
               .std__pe31__lane24_strm0_cntl          ( std__pe31__lane24_strm0_cntl       ),      
               .std__pe31__lane24_strm0_data          ( std__pe31__lane24_strm0_data       ),      
               .std__pe31__lane24_strm0_data_valid    ( std__pe31__lane24_strm0_data_valid ),      
               .std__pe31__lane24_strm0_data_mask     ( std__pe31__lane24_strm0_data_mask  ),      

               .pe31__std__lane24_strm1_ready         ( pe31__std__lane24_strm1_ready      ),      
               .std__pe31__lane24_strm1_cntl          ( std__pe31__lane24_strm1_cntl       ),      
               .std__pe31__lane24_strm1_data          ( std__pe31__lane24_strm1_data       ),      
               .std__pe31__lane24_strm1_data_valid    ( std__pe31__lane24_strm1_data_valid ),      
               .std__pe31__lane24_strm1_data_mask     ( std__pe31__lane24_strm1_data_mask  ),      

               // PE 31, Lane 25                 
               .pe31__std__lane25_strm0_ready         ( pe31__std__lane25_strm0_ready      ),      
               .std__pe31__lane25_strm0_cntl          ( std__pe31__lane25_strm0_cntl       ),      
               .std__pe31__lane25_strm0_data          ( std__pe31__lane25_strm0_data       ),      
               .std__pe31__lane25_strm0_data_valid    ( std__pe31__lane25_strm0_data_valid ),      
               .std__pe31__lane25_strm0_data_mask     ( std__pe31__lane25_strm0_data_mask  ),      

               .pe31__std__lane25_strm1_ready         ( pe31__std__lane25_strm1_ready      ),      
               .std__pe31__lane25_strm1_cntl          ( std__pe31__lane25_strm1_cntl       ),      
               .std__pe31__lane25_strm1_data          ( std__pe31__lane25_strm1_data       ),      
               .std__pe31__lane25_strm1_data_valid    ( std__pe31__lane25_strm1_data_valid ),      
               .std__pe31__lane25_strm1_data_mask     ( std__pe31__lane25_strm1_data_mask  ),      

               // PE 31, Lane 26                 
               .pe31__std__lane26_strm0_ready         ( pe31__std__lane26_strm0_ready      ),      
               .std__pe31__lane26_strm0_cntl          ( std__pe31__lane26_strm0_cntl       ),      
               .std__pe31__lane26_strm0_data          ( std__pe31__lane26_strm0_data       ),      
               .std__pe31__lane26_strm0_data_valid    ( std__pe31__lane26_strm0_data_valid ),      
               .std__pe31__lane26_strm0_data_mask     ( std__pe31__lane26_strm0_data_mask  ),      

               .pe31__std__lane26_strm1_ready         ( pe31__std__lane26_strm1_ready      ),      
               .std__pe31__lane26_strm1_cntl          ( std__pe31__lane26_strm1_cntl       ),      
               .std__pe31__lane26_strm1_data          ( std__pe31__lane26_strm1_data       ),      
               .std__pe31__lane26_strm1_data_valid    ( std__pe31__lane26_strm1_data_valid ),      
               .std__pe31__lane26_strm1_data_mask     ( std__pe31__lane26_strm1_data_mask  ),      

               // PE 31, Lane 27                 
               .pe31__std__lane27_strm0_ready         ( pe31__std__lane27_strm0_ready      ),      
               .std__pe31__lane27_strm0_cntl          ( std__pe31__lane27_strm0_cntl       ),      
               .std__pe31__lane27_strm0_data          ( std__pe31__lane27_strm0_data       ),      
               .std__pe31__lane27_strm0_data_valid    ( std__pe31__lane27_strm0_data_valid ),      
               .std__pe31__lane27_strm0_data_mask     ( std__pe31__lane27_strm0_data_mask  ),      

               .pe31__std__lane27_strm1_ready         ( pe31__std__lane27_strm1_ready      ),      
               .std__pe31__lane27_strm1_cntl          ( std__pe31__lane27_strm1_cntl       ),      
               .std__pe31__lane27_strm1_data          ( std__pe31__lane27_strm1_data       ),      
               .std__pe31__lane27_strm1_data_valid    ( std__pe31__lane27_strm1_data_valid ),      
               .std__pe31__lane27_strm1_data_mask     ( std__pe31__lane27_strm1_data_mask  ),      

               // PE 31, Lane 28                 
               .pe31__std__lane28_strm0_ready         ( pe31__std__lane28_strm0_ready      ),      
               .std__pe31__lane28_strm0_cntl          ( std__pe31__lane28_strm0_cntl       ),      
               .std__pe31__lane28_strm0_data          ( std__pe31__lane28_strm0_data       ),      
               .std__pe31__lane28_strm0_data_valid    ( std__pe31__lane28_strm0_data_valid ),      
               .std__pe31__lane28_strm0_data_mask     ( std__pe31__lane28_strm0_data_mask  ),      

               .pe31__std__lane28_strm1_ready         ( pe31__std__lane28_strm1_ready      ),      
               .std__pe31__lane28_strm1_cntl          ( std__pe31__lane28_strm1_cntl       ),      
               .std__pe31__lane28_strm1_data          ( std__pe31__lane28_strm1_data       ),      
               .std__pe31__lane28_strm1_data_valid    ( std__pe31__lane28_strm1_data_valid ),      
               .std__pe31__lane28_strm1_data_mask     ( std__pe31__lane28_strm1_data_mask  ),      

               // PE 31, Lane 29                 
               .pe31__std__lane29_strm0_ready         ( pe31__std__lane29_strm0_ready      ),      
               .std__pe31__lane29_strm0_cntl          ( std__pe31__lane29_strm0_cntl       ),      
               .std__pe31__lane29_strm0_data          ( std__pe31__lane29_strm0_data       ),      
               .std__pe31__lane29_strm0_data_valid    ( std__pe31__lane29_strm0_data_valid ),      
               .std__pe31__lane29_strm0_data_mask     ( std__pe31__lane29_strm0_data_mask  ),      

               .pe31__std__lane29_strm1_ready         ( pe31__std__lane29_strm1_ready      ),      
               .std__pe31__lane29_strm1_cntl          ( std__pe31__lane29_strm1_cntl       ),      
               .std__pe31__lane29_strm1_data          ( std__pe31__lane29_strm1_data       ),      
               .std__pe31__lane29_strm1_data_valid    ( std__pe31__lane29_strm1_data_valid ),      
               .std__pe31__lane29_strm1_data_mask     ( std__pe31__lane29_strm1_data_mask  ),      

               // PE 31, Lane 30                 
               .pe31__std__lane30_strm0_ready         ( pe31__std__lane30_strm0_ready      ),      
               .std__pe31__lane30_strm0_cntl          ( std__pe31__lane30_strm0_cntl       ),      
               .std__pe31__lane30_strm0_data          ( std__pe31__lane30_strm0_data       ),      
               .std__pe31__lane30_strm0_data_valid    ( std__pe31__lane30_strm0_data_valid ),      
               .std__pe31__lane30_strm0_data_mask     ( std__pe31__lane30_strm0_data_mask  ),      

               .pe31__std__lane30_strm1_ready         ( pe31__std__lane30_strm1_ready      ),      
               .std__pe31__lane30_strm1_cntl          ( std__pe31__lane30_strm1_cntl       ),      
               .std__pe31__lane30_strm1_data          ( std__pe31__lane30_strm1_data       ),      
               .std__pe31__lane30_strm1_data_valid    ( std__pe31__lane30_strm1_data_valid ),      
               .std__pe31__lane30_strm1_data_mask     ( std__pe31__lane30_strm1_data_mask  ),      

               // PE 31, Lane 31                 
               .pe31__std__lane31_strm0_ready         ( pe31__std__lane31_strm0_ready      ),      
               .std__pe31__lane31_strm0_cntl          ( std__pe31__lane31_strm0_cntl       ),      
               .std__pe31__lane31_strm0_data          ( std__pe31__lane31_strm0_data       ),      
               .std__pe31__lane31_strm0_data_valid    ( std__pe31__lane31_strm0_data_valid ),      
               .std__pe31__lane31_strm0_data_mask     ( std__pe31__lane31_strm0_data_mask  ),      

               .pe31__std__lane31_strm1_ready         ( pe31__std__lane31_strm1_ready      ),      
               .std__pe31__lane31_strm1_cntl          ( std__pe31__lane31_strm1_cntl       ),      
               .std__pe31__lane31_strm1_data          ( std__pe31__lane31_strm1_data       ),      
               .std__pe31__lane31_strm1_data_valid    ( std__pe31__lane31_strm1_data_valid ),      
               .std__pe31__lane31_strm1_data_mask     ( std__pe31__lane31_strm1_data_mask  ),      

               // PE 32, Lane 0                 
               .pe32__std__lane0_strm0_ready         ( pe32__std__lane0_strm0_ready      ),      
               .std__pe32__lane0_strm0_cntl          ( std__pe32__lane0_strm0_cntl       ),      
               .std__pe32__lane0_strm0_data          ( std__pe32__lane0_strm0_data       ),      
               .std__pe32__lane0_strm0_data_valid    ( std__pe32__lane0_strm0_data_valid ),      
               .std__pe32__lane0_strm0_data_mask     ( std__pe32__lane0_strm0_data_mask  ),      

               .pe32__std__lane0_strm1_ready         ( pe32__std__lane0_strm1_ready      ),      
               .std__pe32__lane0_strm1_cntl          ( std__pe32__lane0_strm1_cntl       ),      
               .std__pe32__lane0_strm1_data          ( std__pe32__lane0_strm1_data       ),      
               .std__pe32__lane0_strm1_data_valid    ( std__pe32__lane0_strm1_data_valid ),      
               .std__pe32__lane0_strm1_data_mask     ( std__pe32__lane0_strm1_data_mask  ),      

               // PE 32, Lane 1                 
               .pe32__std__lane1_strm0_ready         ( pe32__std__lane1_strm0_ready      ),      
               .std__pe32__lane1_strm0_cntl          ( std__pe32__lane1_strm0_cntl       ),      
               .std__pe32__lane1_strm0_data          ( std__pe32__lane1_strm0_data       ),      
               .std__pe32__lane1_strm0_data_valid    ( std__pe32__lane1_strm0_data_valid ),      
               .std__pe32__lane1_strm0_data_mask     ( std__pe32__lane1_strm0_data_mask  ),      

               .pe32__std__lane1_strm1_ready         ( pe32__std__lane1_strm1_ready      ),      
               .std__pe32__lane1_strm1_cntl          ( std__pe32__lane1_strm1_cntl       ),      
               .std__pe32__lane1_strm1_data          ( std__pe32__lane1_strm1_data       ),      
               .std__pe32__lane1_strm1_data_valid    ( std__pe32__lane1_strm1_data_valid ),      
               .std__pe32__lane1_strm1_data_mask     ( std__pe32__lane1_strm1_data_mask  ),      

               // PE 32, Lane 2                 
               .pe32__std__lane2_strm0_ready         ( pe32__std__lane2_strm0_ready      ),      
               .std__pe32__lane2_strm0_cntl          ( std__pe32__lane2_strm0_cntl       ),      
               .std__pe32__lane2_strm0_data          ( std__pe32__lane2_strm0_data       ),      
               .std__pe32__lane2_strm0_data_valid    ( std__pe32__lane2_strm0_data_valid ),      
               .std__pe32__lane2_strm0_data_mask     ( std__pe32__lane2_strm0_data_mask  ),      

               .pe32__std__lane2_strm1_ready         ( pe32__std__lane2_strm1_ready      ),      
               .std__pe32__lane2_strm1_cntl          ( std__pe32__lane2_strm1_cntl       ),      
               .std__pe32__lane2_strm1_data          ( std__pe32__lane2_strm1_data       ),      
               .std__pe32__lane2_strm1_data_valid    ( std__pe32__lane2_strm1_data_valid ),      
               .std__pe32__lane2_strm1_data_mask     ( std__pe32__lane2_strm1_data_mask  ),      

               // PE 32, Lane 3                 
               .pe32__std__lane3_strm0_ready         ( pe32__std__lane3_strm0_ready      ),      
               .std__pe32__lane3_strm0_cntl          ( std__pe32__lane3_strm0_cntl       ),      
               .std__pe32__lane3_strm0_data          ( std__pe32__lane3_strm0_data       ),      
               .std__pe32__lane3_strm0_data_valid    ( std__pe32__lane3_strm0_data_valid ),      
               .std__pe32__lane3_strm0_data_mask     ( std__pe32__lane3_strm0_data_mask  ),      

               .pe32__std__lane3_strm1_ready         ( pe32__std__lane3_strm1_ready      ),      
               .std__pe32__lane3_strm1_cntl          ( std__pe32__lane3_strm1_cntl       ),      
               .std__pe32__lane3_strm1_data          ( std__pe32__lane3_strm1_data       ),      
               .std__pe32__lane3_strm1_data_valid    ( std__pe32__lane3_strm1_data_valid ),      
               .std__pe32__lane3_strm1_data_mask     ( std__pe32__lane3_strm1_data_mask  ),      

               // PE 32, Lane 4                 
               .pe32__std__lane4_strm0_ready         ( pe32__std__lane4_strm0_ready      ),      
               .std__pe32__lane4_strm0_cntl          ( std__pe32__lane4_strm0_cntl       ),      
               .std__pe32__lane4_strm0_data          ( std__pe32__lane4_strm0_data       ),      
               .std__pe32__lane4_strm0_data_valid    ( std__pe32__lane4_strm0_data_valid ),      
               .std__pe32__lane4_strm0_data_mask     ( std__pe32__lane4_strm0_data_mask  ),      

               .pe32__std__lane4_strm1_ready         ( pe32__std__lane4_strm1_ready      ),      
               .std__pe32__lane4_strm1_cntl          ( std__pe32__lane4_strm1_cntl       ),      
               .std__pe32__lane4_strm1_data          ( std__pe32__lane4_strm1_data       ),      
               .std__pe32__lane4_strm1_data_valid    ( std__pe32__lane4_strm1_data_valid ),      
               .std__pe32__lane4_strm1_data_mask     ( std__pe32__lane4_strm1_data_mask  ),      

               // PE 32, Lane 5                 
               .pe32__std__lane5_strm0_ready         ( pe32__std__lane5_strm0_ready      ),      
               .std__pe32__lane5_strm0_cntl          ( std__pe32__lane5_strm0_cntl       ),      
               .std__pe32__lane5_strm0_data          ( std__pe32__lane5_strm0_data       ),      
               .std__pe32__lane5_strm0_data_valid    ( std__pe32__lane5_strm0_data_valid ),      
               .std__pe32__lane5_strm0_data_mask     ( std__pe32__lane5_strm0_data_mask  ),      

               .pe32__std__lane5_strm1_ready         ( pe32__std__lane5_strm1_ready      ),      
               .std__pe32__lane5_strm1_cntl          ( std__pe32__lane5_strm1_cntl       ),      
               .std__pe32__lane5_strm1_data          ( std__pe32__lane5_strm1_data       ),      
               .std__pe32__lane5_strm1_data_valid    ( std__pe32__lane5_strm1_data_valid ),      
               .std__pe32__lane5_strm1_data_mask     ( std__pe32__lane5_strm1_data_mask  ),      

               // PE 32, Lane 6                 
               .pe32__std__lane6_strm0_ready         ( pe32__std__lane6_strm0_ready      ),      
               .std__pe32__lane6_strm0_cntl          ( std__pe32__lane6_strm0_cntl       ),      
               .std__pe32__lane6_strm0_data          ( std__pe32__lane6_strm0_data       ),      
               .std__pe32__lane6_strm0_data_valid    ( std__pe32__lane6_strm0_data_valid ),      
               .std__pe32__lane6_strm0_data_mask     ( std__pe32__lane6_strm0_data_mask  ),      

               .pe32__std__lane6_strm1_ready         ( pe32__std__lane6_strm1_ready      ),      
               .std__pe32__lane6_strm1_cntl          ( std__pe32__lane6_strm1_cntl       ),      
               .std__pe32__lane6_strm1_data          ( std__pe32__lane6_strm1_data       ),      
               .std__pe32__lane6_strm1_data_valid    ( std__pe32__lane6_strm1_data_valid ),      
               .std__pe32__lane6_strm1_data_mask     ( std__pe32__lane6_strm1_data_mask  ),      

               // PE 32, Lane 7                 
               .pe32__std__lane7_strm0_ready         ( pe32__std__lane7_strm0_ready      ),      
               .std__pe32__lane7_strm0_cntl          ( std__pe32__lane7_strm0_cntl       ),      
               .std__pe32__lane7_strm0_data          ( std__pe32__lane7_strm0_data       ),      
               .std__pe32__lane7_strm0_data_valid    ( std__pe32__lane7_strm0_data_valid ),      
               .std__pe32__lane7_strm0_data_mask     ( std__pe32__lane7_strm0_data_mask  ),      

               .pe32__std__lane7_strm1_ready         ( pe32__std__lane7_strm1_ready      ),      
               .std__pe32__lane7_strm1_cntl          ( std__pe32__lane7_strm1_cntl       ),      
               .std__pe32__lane7_strm1_data          ( std__pe32__lane7_strm1_data       ),      
               .std__pe32__lane7_strm1_data_valid    ( std__pe32__lane7_strm1_data_valid ),      
               .std__pe32__lane7_strm1_data_mask     ( std__pe32__lane7_strm1_data_mask  ),      

               // PE 32, Lane 8                 
               .pe32__std__lane8_strm0_ready         ( pe32__std__lane8_strm0_ready      ),      
               .std__pe32__lane8_strm0_cntl          ( std__pe32__lane8_strm0_cntl       ),      
               .std__pe32__lane8_strm0_data          ( std__pe32__lane8_strm0_data       ),      
               .std__pe32__lane8_strm0_data_valid    ( std__pe32__lane8_strm0_data_valid ),      
               .std__pe32__lane8_strm0_data_mask     ( std__pe32__lane8_strm0_data_mask  ),      

               .pe32__std__lane8_strm1_ready         ( pe32__std__lane8_strm1_ready      ),      
               .std__pe32__lane8_strm1_cntl          ( std__pe32__lane8_strm1_cntl       ),      
               .std__pe32__lane8_strm1_data          ( std__pe32__lane8_strm1_data       ),      
               .std__pe32__lane8_strm1_data_valid    ( std__pe32__lane8_strm1_data_valid ),      
               .std__pe32__lane8_strm1_data_mask     ( std__pe32__lane8_strm1_data_mask  ),      

               // PE 32, Lane 9                 
               .pe32__std__lane9_strm0_ready         ( pe32__std__lane9_strm0_ready      ),      
               .std__pe32__lane9_strm0_cntl          ( std__pe32__lane9_strm0_cntl       ),      
               .std__pe32__lane9_strm0_data          ( std__pe32__lane9_strm0_data       ),      
               .std__pe32__lane9_strm0_data_valid    ( std__pe32__lane9_strm0_data_valid ),      
               .std__pe32__lane9_strm0_data_mask     ( std__pe32__lane9_strm0_data_mask  ),      

               .pe32__std__lane9_strm1_ready         ( pe32__std__lane9_strm1_ready      ),      
               .std__pe32__lane9_strm1_cntl          ( std__pe32__lane9_strm1_cntl       ),      
               .std__pe32__lane9_strm1_data          ( std__pe32__lane9_strm1_data       ),      
               .std__pe32__lane9_strm1_data_valid    ( std__pe32__lane9_strm1_data_valid ),      
               .std__pe32__lane9_strm1_data_mask     ( std__pe32__lane9_strm1_data_mask  ),      

               // PE 32, Lane 10                 
               .pe32__std__lane10_strm0_ready         ( pe32__std__lane10_strm0_ready      ),      
               .std__pe32__lane10_strm0_cntl          ( std__pe32__lane10_strm0_cntl       ),      
               .std__pe32__lane10_strm0_data          ( std__pe32__lane10_strm0_data       ),      
               .std__pe32__lane10_strm0_data_valid    ( std__pe32__lane10_strm0_data_valid ),      
               .std__pe32__lane10_strm0_data_mask     ( std__pe32__lane10_strm0_data_mask  ),      

               .pe32__std__lane10_strm1_ready         ( pe32__std__lane10_strm1_ready      ),      
               .std__pe32__lane10_strm1_cntl          ( std__pe32__lane10_strm1_cntl       ),      
               .std__pe32__lane10_strm1_data          ( std__pe32__lane10_strm1_data       ),      
               .std__pe32__lane10_strm1_data_valid    ( std__pe32__lane10_strm1_data_valid ),      
               .std__pe32__lane10_strm1_data_mask     ( std__pe32__lane10_strm1_data_mask  ),      

               // PE 32, Lane 11                 
               .pe32__std__lane11_strm0_ready         ( pe32__std__lane11_strm0_ready      ),      
               .std__pe32__lane11_strm0_cntl          ( std__pe32__lane11_strm0_cntl       ),      
               .std__pe32__lane11_strm0_data          ( std__pe32__lane11_strm0_data       ),      
               .std__pe32__lane11_strm0_data_valid    ( std__pe32__lane11_strm0_data_valid ),      
               .std__pe32__lane11_strm0_data_mask     ( std__pe32__lane11_strm0_data_mask  ),      

               .pe32__std__lane11_strm1_ready         ( pe32__std__lane11_strm1_ready      ),      
               .std__pe32__lane11_strm1_cntl          ( std__pe32__lane11_strm1_cntl       ),      
               .std__pe32__lane11_strm1_data          ( std__pe32__lane11_strm1_data       ),      
               .std__pe32__lane11_strm1_data_valid    ( std__pe32__lane11_strm1_data_valid ),      
               .std__pe32__lane11_strm1_data_mask     ( std__pe32__lane11_strm1_data_mask  ),      

               // PE 32, Lane 12                 
               .pe32__std__lane12_strm0_ready         ( pe32__std__lane12_strm0_ready      ),      
               .std__pe32__lane12_strm0_cntl          ( std__pe32__lane12_strm0_cntl       ),      
               .std__pe32__lane12_strm0_data          ( std__pe32__lane12_strm0_data       ),      
               .std__pe32__lane12_strm0_data_valid    ( std__pe32__lane12_strm0_data_valid ),      
               .std__pe32__lane12_strm0_data_mask     ( std__pe32__lane12_strm0_data_mask  ),      

               .pe32__std__lane12_strm1_ready         ( pe32__std__lane12_strm1_ready      ),      
               .std__pe32__lane12_strm1_cntl          ( std__pe32__lane12_strm1_cntl       ),      
               .std__pe32__lane12_strm1_data          ( std__pe32__lane12_strm1_data       ),      
               .std__pe32__lane12_strm1_data_valid    ( std__pe32__lane12_strm1_data_valid ),      
               .std__pe32__lane12_strm1_data_mask     ( std__pe32__lane12_strm1_data_mask  ),      

               // PE 32, Lane 13                 
               .pe32__std__lane13_strm0_ready         ( pe32__std__lane13_strm0_ready      ),      
               .std__pe32__lane13_strm0_cntl          ( std__pe32__lane13_strm0_cntl       ),      
               .std__pe32__lane13_strm0_data          ( std__pe32__lane13_strm0_data       ),      
               .std__pe32__lane13_strm0_data_valid    ( std__pe32__lane13_strm0_data_valid ),      
               .std__pe32__lane13_strm0_data_mask     ( std__pe32__lane13_strm0_data_mask  ),      

               .pe32__std__lane13_strm1_ready         ( pe32__std__lane13_strm1_ready      ),      
               .std__pe32__lane13_strm1_cntl          ( std__pe32__lane13_strm1_cntl       ),      
               .std__pe32__lane13_strm1_data          ( std__pe32__lane13_strm1_data       ),      
               .std__pe32__lane13_strm1_data_valid    ( std__pe32__lane13_strm1_data_valid ),      
               .std__pe32__lane13_strm1_data_mask     ( std__pe32__lane13_strm1_data_mask  ),      

               // PE 32, Lane 14                 
               .pe32__std__lane14_strm0_ready         ( pe32__std__lane14_strm0_ready      ),      
               .std__pe32__lane14_strm0_cntl          ( std__pe32__lane14_strm0_cntl       ),      
               .std__pe32__lane14_strm0_data          ( std__pe32__lane14_strm0_data       ),      
               .std__pe32__lane14_strm0_data_valid    ( std__pe32__lane14_strm0_data_valid ),      
               .std__pe32__lane14_strm0_data_mask     ( std__pe32__lane14_strm0_data_mask  ),      

               .pe32__std__lane14_strm1_ready         ( pe32__std__lane14_strm1_ready      ),      
               .std__pe32__lane14_strm1_cntl          ( std__pe32__lane14_strm1_cntl       ),      
               .std__pe32__lane14_strm1_data          ( std__pe32__lane14_strm1_data       ),      
               .std__pe32__lane14_strm1_data_valid    ( std__pe32__lane14_strm1_data_valid ),      
               .std__pe32__lane14_strm1_data_mask     ( std__pe32__lane14_strm1_data_mask  ),      

               // PE 32, Lane 15                 
               .pe32__std__lane15_strm0_ready         ( pe32__std__lane15_strm0_ready      ),      
               .std__pe32__lane15_strm0_cntl          ( std__pe32__lane15_strm0_cntl       ),      
               .std__pe32__lane15_strm0_data          ( std__pe32__lane15_strm0_data       ),      
               .std__pe32__lane15_strm0_data_valid    ( std__pe32__lane15_strm0_data_valid ),      
               .std__pe32__lane15_strm0_data_mask     ( std__pe32__lane15_strm0_data_mask  ),      

               .pe32__std__lane15_strm1_ready         ( pe32__std__lane15_strm1_ready      ),      
               .std__pe32__lane15_strm1_cntl          ( std__pe32__lane15_strm1_cntl       ),      
               .std__pe32__lane15_strm1_data          ( std__pe32__lane15_strm1_data       ),      
               .std__pe32__lane15_strm1_data_valid    ( std__pe32__lane15_strm1_data_valid ),      
               .std__pe32__lane15_strm1_data_mask     ( std__pe32__lane15_strm1_data_mask  ),      

               // PE 32, Lane 16                 
               .pe32__std__lane16_strm0_ready         ( pe32__std__lane16_strm0_ready      ),      
               .std__pe32__lane16_strm0_cntl          ( std__pe32__lane16_strm0_cntl       ),      
               .std__pe32__lane16_strm0_data          ( std__pe32__lane16_strm0_data       ),      
               .std__pe32__lane16_strm0_data_valid    ( std__pe32__lane16_strm0_data_valid ),      
               .std__pe32__lane16_strm0_data_mask     ( std__pe32__lane16_strm0_data_mask  ),      

               .pe32__std__lane16_strm1_ready         ( pe32__std__lane16_strm1_ready      ),      
               .std__pe32__lane16_strm1_cntl          ( std__pe32__lane16_strm1_cntl       ),      
               .std__pe32__lane16_strm1_data          ( std__pe32__lane16_strm1_data       ),      
               .std__pe32__lane16_strm1_data_valid    ( std__pe32__lane16_strm1_data_valid ),      
               .std__pe32__lane16_strm1_data_mask     ( std__pe32__lane16_strm1_data_mask  ),      

               // PE 32, Lane 17                 
               .pe32__std__lane17_strm0_ready         ( pe32__std__lane17_strm0_ready      ),      
               .std__pe32__lane17_strm0_cntl          ( std__pe32__lane17_strm0_cntl       ),      
               .std__pe32__lane17_strm0_data          ( std__pe32__lane17_strm0_data       ),      
               .std__pe32__lane17_strm0_data_valid    ( std__pe32__lane17_strm0_data_valid ),      
               .std__pe32__lane17_strm0_data_mask     ( std__pe32__lane17_strm0_data_mask  ),      

               .pe32__std__lane17_strm1_ready         ( pe32__std__lane17_strm1_ready      ),      
               .std__pe32__lane17_strm1_cntl          ( std__pe32__lane17_strm1_cntl       ),      
               .std__pe32__lane17_strm1_data          ( std__pe32__lane17_strm1_data       ),      
               .std__pe32__lane17_strm1_data_valid    ( std__pe32__lane17_strm1_data_valid ),      
               .std__pe32__lane17_strm1_data_mask     ( std__pe32__lane17_strm1_data_mask  ),      

               // PE 32, Lane 18                 
               .pe32__std__lane18_strm0_ready         ( pe32__std__lane18_strm0_ready      ),      
               .std__pe32__lane18_strm0_cntl          ( std__pe32__lane18_strm0_cntl       ),      
               .std__pe32__lane18_strm0_data          ( std__pe32__lane18_strm0_data       ),      
               .std__pe32__lane18_strm0_data_valid    ( std__pe32__lane18_strm0_data_valid ),      
               .std__pe32__lane18_strm0_data_mask     ( std__pe32__lane18_strm0_data_mask  ),      

               .pe32__std__lane18_strm1_ready         ( pe32__std__lane18_strm1_ready      ),      
               .std__pe32__lane18_strm1_cntl          ( std__pe32__lane18_strm1_cntl       ),      
               .std__pe32__lane18_strm1_data          ( std__pe32__lane18_strm1_data       ),      
               .std__pe32__lane18_strm1_data_valid    ( std__pe32__lane18_strm1_data_valid ),      
               .std__pe32__lane18_strm1_data_mask     ( std__pe32__lane18_strm1_data_mask  ),      

               // PE 32, Lane 19                 
               .pe32__std__lane19_strm0_ready         ( pe32__std__lane19_strm0_ready      ),      
               .std__pe32__lane19_strm0_cntl          ( std__pe32__lane19_strm0_cntl       ),      
               .std__pe32__lane19_strm0_data          ( std__pe32__lane19_strm0_data       ),      
               .std__pe32__lane19_strm0_data_valid    ( std__pe32__lane19_strm0_data_valid ),      
               .std__pe32__lane19_strm0_data_mask     ( std__pe32__lane19_strm0_data_mask  ),      

               .pe32__std__lane19_strm1_ready         ( pe32__std__lane19_strm1_ready      ),      
               .std__pe32__lane19_strm1_cntl          ( std__pe32__lane19_strm1_cntl       ),      
               .std__pe32__lane19_strm1_data          ( std__pe32__lane19_strm1_data       ),      
               .std__pe32__lane19_strm1_data_valid    ( std__pe32__lane19_strm1_data_valid ),      
               .std__pe32__lane19_strm1_data_mask     ( std__pe32__lane19_strm1_data_mask  ),      

               // PE 32, Lane 20                 
               .pe32__std__lane20_strm0_ready         ( pe32__std__lane20_strm0_ready      ),      
               .std__pe32__lane20_strm0_cntl          ( std__pe32__lane20_strm0_cntl       ),      
               .std__pe32__lane20_strm0_data          ( std__pe32__lane20_strm0_data       ),      
               .std__pe32__lane20_strm0_data_valid    ( std__pe32__lane20_strm0_data_valid ),      
               .std__pe32__lane20_strm0_data_mask     ( std__pe32__lane20_strm0_data_mask  ),      

               .pe32__std__lane20_strm1_ready         ( pe32__std__lane20_strm1_ready      ),      
               .std__pe32__lane20_strm1_cntl          ( std__pe32__lane20_strm1_cntl       ),      
               .std__pe32__lane20_strm1_data          ( std__pe32__lane20_strm1_data       ),      
               .std__pe32__lane20_strm1_data_valid    ( std__pe32__lane20_strm1_data_valid ),      
               .std__pe32__lane20_strm1_data_mask     ( std__pe32__lane20_strm1_data_mask  ),      

               // PE 32, Lane 21                 
               .pe32__std__lane21_strm0_ready         ( pe32__std__lane21_strm0_ready      ),      
               .std__pe32__lane21_strm0_cntl          ( std__pe32__lane21_strm0_cntl       ),      
               .std__pe32__lane21_strm0_data          ( std__pe32__lane21_strm0_data       ),      
               .std__pe32__lane21_strm0_data_valid    ( std__pe32__lane21_strm0_data_valid ),      
               .std__pe32__lane21_strm0_data_mask     ( std__pe32__lane21_strm0_data_mask  ),      

               .pe32__std__lane21_strm1_ready         ( pe32__std__lane21_strm1_ready      ),      
               .std__pe32__lane21_strm1_cntl          ( std__pe32__lane21_strm1_cntl       ),      
               .std__pe32__lane21_strm1_data          ( std__pe32__lane21_strm1_data       ),      
               .std__pe32__lane21_strm1_data_valid    ( std__pe32__lane21_strm1_data_valid ),      
               .std__pe32__lane21_strm1_data_mask     ( std__pe32__lane21_strm1_data_mask  ),      

               // PE 32, Lane 22                 
               .pe32__std__lane22_strm0_ready         ( pe32__std__lane22_strm0_ready      ),      
               .std__pe32__lane22_strm0_cntl          ( std__pe32__lane22_strm0_cntl       ),      
               .std__pe32__lane22_strm0_data          ( std__pe32__lane22_strm0_data       ),      
               .std__pe32__lane22_strm0_data_valid    ( std__pe32__lane22_strm0_data_valid ),      
               .std__pe32__lane22_strm0_data_mask     ( std__pe32__lane22_strm0_data_mask  ),      

               .pe32__std__lane22_strm1_ready         ( pe32__std__lane22_strm1_ready      ),      
               .std__pe32__lane22_strm1_cntl          ( std__pe32__lane22_strm1_cntl       ),      
               .std__pe32__lane22_strm1_data          ( std__pe32__lane22_strm1_data       ),      
               .std__pe32__lane22_strm1_data_valid    ( std__pe32__lane22_strm1_data_valid ),      
               .std__pe32__lane22_strm1_data_mask     ( std__pe32__lane22_strm1_data_mask  ),      

               // PE 32, Lane 23                 
               .pe32__std__lane23_strm0_ready         ( pe32__std__lane23_strm0_ready      ),      
               .std__pe32__lane23_strm0_cntl          ( std__pe32__lane23_strm0_cntl       ),      
               .std__pe32__lane23_strm0_data          ( std__pe32__lane23_strm0_data       ),      
               .std__pe32__lane23_strm0_data_valid    ( std__pe32__lane23_strm0_data_valid ),      
               .std__pe32__lane23_strm0_data_mask     ( std__pe32__lane23_strm0_data_mask  ),      

               .pe32__std__lane23_strm1_ready         ( pe32__std__lane23_strm1_ready      ),      
               .std__pe32__lane23_strm1_cntl          ( std__pe32__lane23_strm1_cntl       ),      
               .std__pe32__lane23_strm1_data          ( std__pe32__lane23_strm1_data       ),      
               .std__pe32__lane23_strm1_data_valid    ( std__pe32__lane23_strm1_data_valid ),      
               .std__pe32__lane23_strm1_data_mask     ( std__pe32__lane23_strm1_data_mask  ),      

               // PE 32, Lane 24                 
               .pe32__std__lane24_strm0_ready         ( pe32__std__lane24_strm0_ready      ),      
               .std__pe32__lane24_strm0_cntl          ( std__pe32__lane24_strm0_cntl       ),      
               .std__pe32__lane24_strm0_data          ( std__pe32__lane24_strm0_data       ),      
               .std__pe32__lane24_strm0_data_valid    ( std__pe32__lane24_strm0_data_valid ),      
               .std__pe32__lane24_strm0_data_mask     ( std__pe32__lane24_strm0_data_mask  ),      

               .pe32__std__lane24_strm1_ready         ( pe32__std__lane24_strm1_ready      ),      
               .std__pe32__lane24_strm1_cntl          ( std__pe32__lane24_strm1_cntl       ),      
               .std__pe32__lane24_strm1_data          ( std__pe32__lane24_strm1_data       ),      
               .std__pe32__lane24_strm1_data_valid    ( std__pe32__lane24_strm1_data_valid ),      
               .std__pe32__lane24_strm1_data_mask     ( std__pe32__lane24_strm1_data_mask  ),      

               // PE 32, Lane 25                 
               .pe32__std__lane25_strm0_ready         ( pe32__std__lane25_strm0_ready      ),      
               .std__pe32__lane25_strm0_cntl          ( std__pe32__lane25_strm0_cntl       ),      
               .std__pe32__lane25_strm0_data          ( std__pe32__lane25_strm0_data       ),      
               .std__pe32__lane25_strm0_data_valid    ( std__pe32__lane25_strm0_data_valid ),      
               .std__pe32__lane25_strm0_data_mask     ( std__pe32__lane25_strm0_data_mask  ),      

               .pe32__std__lane25_strm1_ready         ( pe32__std__lane25_strm1_ready      ),      
               .std__pe32__lane25_strm1_cntl          ( std__pe32__lane25_strm1_cntl       ),      
               .std__pe32__lane25_strm1_data          ( std__pe32__lane25_strm1_data       ),      
               .std__pe32__lane25_strm1_data_valid    ( std__pe32__lane25_strm1_data_valid ),      
               .std__pe32__lane25_strm1_data_mask     ( std__pe32__lane25_strm1_data_mask  ),      

               // PE 32, Lane 26                 
               .pe32__std__lane26_strm0_ready         ( pe32__std__lane26_strm0_ready      ),      
               .std__pe32__lane26_strm0_cntl          ( std__pe32__lane26_strm0_cntl       ),      
               .std__pe32__lane26_strm0_data          ( std__pe32__lane26_strm0_data       ),      
               .std__pe32__lane26_strm0_data_valid    ( std__pe32__lane26_strm0_data_valid ),      
               .std__pe32__lane26_strm0_data_mask     ( std__pe32__lane26_strm0_data_mask  ),      

               .pe32__std__lane26_strm1_ready         ( pe32__std__lane26_strm1_ready      ),      
               .std__pe32__lane26_strm1_cntl          ( std__pe32__lane26_strm1_cntl       ),      
               .std__pe32__lane26_strm1_data          ( std__pe32__lane26_strm1_data       ),      
               .std__pe32__lane26_strm1_data_valid    ( std__pe32__lane26_strm1_data_valid ),      
               .std__pe32__lane26_strm1_data_mask     ( std__pe32__lane26_strm1_data_mask  ),      

               // PE 32, Lane 27                 
               .pe32__std__lane27_strm0_ready         ( pe32__std__lane27_strm0_ready      ),      
               .std__pe32__lane27_strm0_cntl          ( std__pe32__lane27_strm0_cntl       ),      
               .std__pe32__lane27_strm0_data          ( std__pe32__lane27_strm0_data       ),      
               .std__pe32__lane27_strm0_data_valid    ( std__pe32__lane27_strm0_data_valid ),      
               .std__pe32__lane27_strm0_data_mask     ( std__pe32__lane27_strm0_data_mask  ),      

               .pe32__std__lane27_strm1_ready         ( pe32__std__lane27_strm1_ready      ),      
               .std__pe32__lane27_strm1_cntl          ( std__pe32__lane27_strm1_cntl       ),      
               .std__pe32__lane27_strm1_data          ( std__pe32__lane27_strm1_data       ),      
               .std__pe32__lane27_strm1_data_valid    ( std__pe32__lane27_strm1_data_valid ),      
               .std__pe32__lane27_strm1_data_mask     ( std__pe32__lane27_strm1_data_mask  ),      

               // PE 32, Lane 28                 
               .pe32__std__lane28_strm0_ready         ( pe32__std__lane28_strm0_ready      ),      
               .std__pe32__lane28_strm0_cntl          ( std__pe32__lane28_strm0_cntl       ),      
               .std__pe32__lane28_strm0_data          ( std__pe32__lane28_strm0_data       ),      
               .std__pe32__lane28_strm0_data_valid    ( std__pe32__lane28_strm0_data_valid ),      
               .std__pe32__lane28_strm0_data_mask     ( std__pe32__lane28_strm0_data_mask  ),      

               .pe32__std__lane28_strm1_ready         ( pe32__std__lane28_strm1_ready      ),      
               .std__pe32__lane28_strm1_cntl          ( std__pe32__lane28_strm1_cntl       ),      
               .std__pe32__lane28_strm1_data          ( std__pe32__lane28_strm1_data       ),      
               .std__pe32__lane28_strm1_data_valid    ( std__pe32__lane28_strm1_data_valid ),      
               .std__pe32__lane28_strm1_data_mask     ( std__pe32__lane28_strm1_data_mask  ),      

               // PE 32, Lane 29                 
               .pe32__std__lane29_strm0_ready         ( pe32__std__lane29_strm0_ready      ),      
               .std__pe32__lane29_strm0_cntl          ( std__pe32__lane29_strm0_cntl       ),      
               .std__pe32__lane29_strm0_data          ( std__pe32__lane29_strm0_data       ),      
               .std__pe32__lane29_strm0_data_valid    ( std__pe32__lane29_strm0_data_valid ),      
               .std__pe32__lane29_strm0_data_mask     ( std__pe32__lane29_strm0_data_mask  ),      

               .pe32__std__lane29_strm1_ready         ( pe32__std__lane29_strm1_ready      ),      
               .std__pe32__lane29_strm1_cntl          ( std__pe32__lane29_strm1_cntl       ),      
               .std__pe32__lane29_strm1_data          ( std__pe32__lane29_strm1_data       ),      
               .std__pe32__lane29_strm1_data_valid    ( std__pe32__lane29_strm1_data_valid ),      
               .std__pe32__lane29_strm1_data_mask     ( std__pe32__lane29_strm1_data_mask  ),      

               // PE 32, Lane 30                 
               .pe32__std__lane30_strm0_ready         ( pe32__std__lane30_strm0_ready      ),      
               .std__pe32__lane30_strm0_cntl          ( std__pe32__lane30_strm0_cntl       ),      
               .std__pe32__lane30_strm0_data          ( std__pe32__lane30_strm0_data       ),      
               .std__pe32__lane30_strm0_data_valid    ( std__pe32__lane30_strm0_data_valid ),      
               .std__pe32__lane30_strm0_data_mask     ( std__pe32__lane30_strm0_data_mask  ),      

               .pe32__std__lane30_strm1_ready         ( pe32__std__lane30_strm1_ready      ),      
               .std__pe32__lane30_strm1_cntl          ( std__pe32__lane30_strm1_cntl       ),      
               .std__pe32__lane30_strm1_data          ( std__pe32__lane30_strm1_data       ),      
               .std__pe32__lane30_strm1_data_valid    ( std__pe32__lane30_strm1_data_valid ),      
               .std__pe32__lane30_strm1_data_mask     ( std__pe32__lane30_strm1_data_mask  ),      

               // PE 32, Lane 31                 
               .pe32__std__lane31_strm0_ready         ( pe32__std__lane31_strm0_ready      ),      
               .std__pe32__lane31_strm0_cntl          ( std__pe32__lane31_strm0_cntl       ),      
               .std__pe32__lane31_strm0_data          ( std__pe32__lane31_strm0_data       ),      
               .std__pe32__lane31_strm0_data_valid    ( std__pe32__lane31_strm0_data_valid ),      
               .std__pe32__lane31_strm0_data_mask     ( std__pe32__lane31_strm0_data_mask  ),      

               .pe32__std__lane31_strm1_ready         ( pe32__std__lane31_strm1_ready      ),      
               .std__pe32__lane31_strm1_cntl          ( std__pe32__lane31_strm1_cntl       ),      
               .std__pe32__lane31_strm1_data          ( std__pe32__lane31_strm1_data       ),      
               .std__pe32__lane31_strm1_data_valid    ( std__pe32__lane31_strm1_data_valid ),      
               .std__pe32__lane31_strm1_data_mask     ( std__pe32__lane31_strm1_data_mask  ),      

               // PE 33, Lane 0                 
               .pe33__std__lane0_strm0_ready         ( pe33__std__lane0_strm0_ready      ),      
               .std__pe33__lane0_strm0_cntl          ( std__pe33__lane0_strm0_cntl       ),      
               .std__pe33__lane0_strm0_data          ( std__pe33__lane0_strm0_data       ),      
               .std__pe33__lane0_strm0_data_valid    ( std__pe33__lane0_strm0_data_valid ),      
               .std__pe33__lane0_strm0_data_mask     ( std__pe33__lane0_strm0_data_mask  ),      

               .pe33__std__lane0_strm1_ready         ( pe33__std__lane0_strm1_ready      ),      
               .std__pe33__lane0_strm1_cntl          ( std__pe33__lane0_strm1_cntl       ),      
               .std__pe33__lane0_strm1_data          ( std__pe33__lane0_strm1_data       ),      
               .std__pe33__lane0_strm1_data_valid    ( std__pe33__lane0_strm1_data_valid ),      
               .std__pe33__lane0_strm1_data_mask     ( std__pe33__lane0_strm1_data_mask  ),      

               // PE 33, Lane 1                 
               .pe33__std__lane1_strm0_ready         ( pe33__std__lane1_strm0_ready      ),      
               .std__pe33__lane1_strm0_cntl          ( std__pe33__lane1_strm0_cntl       ),      
               .std__pe33__lane1_strm0_data          ( std__pe33__lane1_strm0_data       ),      
               .std__pe33__lane1_strm0_data_valid    ( std__pe33__lane1_strm0_data_valid ),      
               .std__pe33__lane1_strm0_data_mask     ( std__pe33__lane1_strm0_data_mask  ),      

               .pe33__std__lane1_strm1_ready         ( pe33__std__lane1_strm1_ready      ),      
               .std__pe33__lane1_strm1_cntl          ( std__pe33__lane1_strm1_cntl       ),      
               .std__pe33__lane1_strm1_data          ( std__pe33__lane1_strm1_data       ),      
               .std__pe33__lane1_strm1_data_valid    ( std__pe33__lane1_strm1_data_valid ),      
               .std__pe33__lane1_strm1_data_mask     ( std__pe33__lane1_strm1_data_mask  ),      

               // PE 33, Lane 2                 
               .pe33__std__lane2_strm0_ready         ( pe33__std__lane2_strm0_ready      ),      
               .std__pe33__lane2_strm0_cntl          ( std__pe33__lane2_strm0_cntl       ),      
               .std__pe33__lane2_strm0_data          ( std__pe33__lane2_strm0_data       ),      
               .std__pe33__lane2_strm0_data_valid    ( std__pe33__lane2_strm0_data_valid ),      
               .std__pe33__lane2_strm0_data_mask     ( std__pe33__lane2_strm0_data_mask  ),      

               .pe33__std__lane2_strm1_ready         ( pe33__std__lane2_strm1_ready      ),      
               .std__pe33__lane2_strm1_cntl          ( std__pe33__lane2_strm1_cntl       ),      
               .std__pe33__lane2_strm1_data          ( std__pe33__lane2_strm1_data       ),      
               .std__pe33__lane2_strm1_data_valid    ( std__pe33__lane2_strm1_data_valid ),      
               .std__pe33__lane2_strm1_data_mask     ( std__pe33__lane2_strm1_data_mask  ),      

               // PE 33, Lane 3                 
               .pe33__std__lane3_strm0_ready         ( pe33__std__lane3_strm0_ready      ),      
               .std__pe33__lane3_strm0_cntl          ( std__pe33__lane3_strm0_cntl       ),      
               .std__pe33__lane3_strm0_data          ( std__pe33__lane3_strm0_data       ),      
               .std__pe33__lane3_strm0_data_valid    ( std__pe33__lane3_strm0_data_valid ),      
               .std__pe33__lane3_strm0_data_mask     ( std__pe33__lane3_strm0_data_mask  ),      

               .pe33__std__lane3_strm1_ready         ( pe33__std__lane3_strm1_ready      ),      
               .std__pe33__lane3_strm1_cntl          ( std__pe33__lane3_strm1_cntl       ),      
               .std__pe33__lane3_strm1_data          ( std__pe33__lane3_strm1_data       ),      
               .std__pe33__lane3_strm1_data_valid    ( std__pe33__lane3_strm1_data_valid ),      
               .std__pe33__lane3_strm1_data_mask     ( std__pe33__lane3_strm1_data_mask  ),      

               // PE 33, Lane 4                 
               .pe33__std__lane4_strm0_ready         ( pe33__std__lane4_strm0_ready      ),      
               .std__pe33__lane4_strm0_cntl          ( std__pe33__lane4_strm0_cntl       ),      
               .std__pe33__lane4_strm0_data          ( std__pe33__lane4_strm0_data       ),      
               .std__pe33__lane4_strm0_data_valid    ( std__pe33__lane4_strm0_data_valid ),      
               .std__pe33__lane4_strm0_data_mask     ( std__pe33__lane4_strm0_data_mask  ),      

               .pe33__std__lane4_strm1_ready         ( pe33__std__lane4_strm1_ready      ),      
               .std__pe33__lane4_strm1_cntl          ( std__pe33__lane4_strm1_cntl       ),      
               .std__pe33__lane4_strm1_data          ( std__pe33__lane4_strm1_data       ),      
               .std__pe33__lane4_strm1_data_valid    ( std__pe33__lane4_strm1_data_valid ),      
               .std__pe33__lane4_strm1_data_mask     ( std__pe33__lane4_strm1_data_mask  ),      

               // PE 33, Lane 5                 
               .pe33__std__lane5_strm0_ready         ( pe33__std__lane5_strm0_ready      ),      
               .std__pe33__lane5_strm0_cntl          ( std__pe33__lane5_strm0_cntl       ),      
               .std__pe33__lane5_strm0_data          ( std__pe33__lane5_strm0_data       ),      
               .std__pe33__lane5_strm0_data_valid    ( std__pe33__lane5_strm0_data_valid ),      
               .std__pe33__lane5_strm0_data_mask     ( std__pe33__lane5_strm0_data_mask  ),      

               .pe33__std__lane5_strm1_ready         ( pe33__std__lane5_strm1_ready      ),      
               .std__pe33__lane5_strm1_cntl          ( std__pe33__lane5_strm1_cntl       ),      
               .std__pe33__lane5_strm1_data          ( std__pe33__lane5_strm1_data       ),      
               .std__pe33__lane5_strm1_data_valid    ( std__pe33__lane5_strm1_data_valid ),      
               .std__pe33__lane5_strm1_data_mask     ( std__pe33__lane5_strm1_data_mask  ),      

               // PE 33, Lane 6                 
               .pe33__std__lane6_strm0_ready         ( pe33__std__lane6_strm0_ready      ),      
               .std__pe33__lane6_strm0_cntl          ( std__pe33__lane6_strm0_cntl       ),      
               .std__pe33__lane6_strm0_data          ( std__pe33__lane6_strm0_data       ),      
               .std__pe33__lane6_strm0_data_valid    ( std__pe33__lane6_strm0_data_valid ),      
               .std__pe33__lane6_strm0_data_mask     ( std__pe33__lane6_strm0_data_mask  ),      

               .pe33__std__lane6_strm1_ready         ( pe33__std__lane6_strm1_ready      ),      
               .std__pe33__lane6_strm1_cntl          ( std__pe33__lane6_strm1_cntl       ),      
               .std__pe33__lane6_strm1_data          ( std__pe33__lane6_strm1_data       ),      
               .std__pe33__lane6_strm1_data_valid    ( std__pe33__lane6_strm1_data_valid ),      
               .std__pe33__lane6_strm1_data_mask     ( std__pe33__lane6_strm1_data_mask  ),      

               // PE 33, Lane 7                 
               .pe33__std__lane7_strm0_ready         ( pe33__std__lane7_strm0_ready      ),      
               .std__pe33__lane7_strm0_cntl          ( std__pe33__lane7_strm0_cntl       ),      
               .std__pe33__lane7_strm0_data          ( std__pe33__lane7_strm0_data       ),      
               .std__pe33__lane7_strm0_data_valid    ( std__pe33__lane7_strm0_data_valid ),      
               .std__pe33__lane7_strm0_data_mask     ( std__pe33__lane7_strm0_data_mask  ),      

               .pe33__std__lane7_strm1_ready         ( pe33__std__lane7_strm1_ready      ),      
               .std__pe33__lane7_strm1_cntl          ( std__pe33__lane7_strm1_cntl       ),      
               .std__pe33__lane7_strm1_data          ( std__pe33__lane7_strm1_data       ),      
               .std__pe33__lane7_strm1_data_valid    ( std__pe33__lane7_strm1_data_valid ),      
               .std__pe33__lane7_strm1_data_mask     ( std__pe33__lane7_strm1_data_mask  ),      

               // PE 33, Lane 8                 
               .pe33__std__lane8_strm0_ready         ( pe33__std__lane8_strm0_ready      ),      
               .std__pe33__lane8_strm0_cntl          ( std__pe33__lane8_strm0_cntl       ),      
               .std__pe33__lane8_strm0_data          ( std__pe33__lane8_strm0_data       ),      
               .std__pe33__lane8_strm0_data_valid    ( std__pe33__lane8_strm0_data_valid ),      
               .std__pe33__lane8_strm0_data_mask     ( std__pe33__lane8_strm0_data_mask  ),      

               .pe33__std__lane8_strm1_ready         ( pe33__std__lane8_strm1_ready      ),      
               .std__pe33__lane8_strm1_cntl          ( std__pe33__lane8_strm1_cntl       ),      
               .std__pe33__lane8_strm1_data          ( std__pe33__lane8_strm1_data       ),      
               .std__pe33__lane8_strm1_data_valid    ( std__pe33__lane8_strm1_data_valid ),      
               .std__pe33__lane8_strm1_data_mask     ( std__pe33__lane8_strm1_data_mask  ),      

               // PE 33, Lane 9                 
               .pe33__std__lane9_strm0_ready         ( pe33__std__lane9_strm0_ready      ),      
               .std__pe33__lane9_strm0_cntl          ( std__pe33__lane9_strm0_cntl       ),      
               .std__pe33__lane9_strm0_data          ( std__pe33__lane9_strm0_data       ),      
               .std__pe33__lane9_strm0_data_valid    ( std__pe33__lane9_strm0_data_valid ),      
               .std__pe33__lane9_strm0_data_mask     ( std__pe33__lane9_strm0_data_mask  ),      

               .pe33__std__lane9_strm1_ready         ( pe33__std__lane9_strm1_ready      ),      
               .std__pe33__lane9_strm1_cntl          ( std__pe33__lane9_strm1_cntl       ),      
               .std__pe33__lane9_strm1_data          ( std__pe33__lane9_strm1_data       ),      
               .std__pe33__lane9_strm1_data_valid    ( std__pe33__lane9_strm1_data_valid ),      
               .std__pe33__lane9_strm1_data_mask     ( std__pe33__lane9_strm1_data_mask  ),      

               // PE 33, Lane 10                 
               .pe33__std__lane10_strm0_ready         ( pe33__std__lane10_strm0_ready      ),      
               .std__pe33__lane10_strm0_cntl          ( std__pe33__lane10_strm0_cntl       ),      
               .std__pe33__lane10_strm0_data          ( std__pe33__lane10_strm0_data       ),      
               .std__pe33__lane10_strm0_data_valid    ( std__pe33__lane10_strm0_data_valid ),      
               .std__pe33__lane10_strm0_data_mask     ( std__pe33__lane10_strm0_data_mask  ),      

               .pe33__std__lane10_strm1_ready         ( pe33__std__lane10_strm1_ready      ),      
               .std__pe33__lane10_strm1_cntl          ( std__pe33__lane10_strm1_cntl       ),      
               .std__pe33__lane10_strm1_data          ( std__pe33__lane10_strm1_data       ),      
               .std__pe33__lane10_strm1_data_valid    ( std__pe33__lane10_strm1_data_valid ),      
               .std__pe33__lane10_strm1_data_mask     ( std__pe33__lane10_strm1_data_mask  ),      

               // PE 33, Lane 11                 
               .pe33__std__lane11_strm0_ready         ( pe33__std__lane11_strm0_ready      ),      
               .std__pe33__lane11_strm0_cntl          ( std__pe33__lane11_strm0_cntl       ),      
               .std__pe33__lane11_strm0_data          ( std__pe33__lane11_strm0_data       ),      
               .std__pe33__lane11_strm0_data_valid    ( std__pe33__lane11_strm0_data_valid ),      
               .std__pe33__lane11_strm0_data_mask     ( std__pe33__lane11_strm0_data_mask  ),      

               .pe33__std__lane11_strm1_ready         ( pe33__std__lane11_strm1_ready      ),      
               .std__pe33__lane11_strm1_cntl          ( std__pe33__lane11_strm1_cntl       ),      
               .std__pe33__lane11_strm1_data          ( std__pe33__lane11_strm1_data       ),      
               .std__pe33__lane11_strm1_data_valid    ( std__pe33__lane11_strm1_data_valid ),      
               .std__pe33__lane11_strm1_data_mask     ( std__pe33__lane11_strm1_data_mask  ),      

               // PE 33, Lane 12                 
               .pe33__std__lane12_strm0_ready         ( pe33__std__lane12_strm0_ready      ),      
               .std__pe33__lane12_strm0_cntl          ( std__pe33__lane12_strm0_cntl       ),      
               .std__pe33__lane12_strm0_data          ( std__pe33__lane12_strm0_data       ),      
               .std__pe33__lane12_strm0_data_valid    ( std__pe33__lane12_strm0_data_valid ),      
               .std__pe33__lane12_strm0_data_mask     ( std__pe33__lane12_strm0_data_mask  ),      

               .pe33__std__lane12_strm1_ready         ( pe33__std__lane12_strm1_ready      ),      
               .std__pe33__lane12_strm1_cntl          ( std__pe33__lane12_strm1_cntl       ),      
               .std__pe33__lane12_strm1_data          ( std__pe33__lane12_strm1_data       ),      
               .std__pe33__lane12_strm1_data_valid    ( std__pe33__lane12_strm1_data_valid ),      
               .std__pe33__lane12_strm1_data_mask     ( std__pe33__lane12_strm1_data_mask  ),      

               // PE 33, Lane 13                 
               .pe33__std__lane13_strm0_ready         ( pe33__std__lane13_strm0_ready      ),      
               .std__pe33__lane13_strm0_cntl          ( std__pe33__lane13_strm0_cntl       ),      
               .std__pe33__lane13_strm0_data          ( std__pe33__lane13_strm0_data       ),      
               .std__pe33__lane13_strm0_data_valid    ( std__pe33__lane13_strm0_data_valid ),      
               .std__pe33__lane13_strm0_data_mask     ( std__pe33__lane13_strm0_data_mask  ),      

               .pe33__std__lane13_strm1_ready         ( pe33__std__lane13_strm1_ready      ),      
               .std__pe33__lane13_strm1_cntl          ( std__pe33__lane13_strm1_cntl       ),      
               .std__pe33__lane13_strm1_data          ( std__pe33__lane13_strm1_data       ),      
               .std__pe33__lane13_strm1_data_valid    ( std__pe33__lane13_strm1_data_valid ),      
               .std__pe33__lane13_strm1_data_mask     ( std__pe33__lane13_strm1_data_mask  ),      

               // PE 33, Lane 14                 
               .pe33__std__lane14_strm0_ready         ( pe33__std__lane14_strm0_ready      ),      
               .std__pe33__lane14_strm0_cntl          ( std__pe33__lane14_strm0_cntl       ),      
               .std__pe33__lane14_strm0_data          ( std__pe33__lane14_strm0_data       ),      
               .std__pe33__lane14_strm0_data_valid    ( std__pe33__lane14_strm0_data_valid ),      
               .std__pe33__lane14_strm0_data_mask     ( std__pe33__lane14_strm0_data_mask  ),      

               .pe33__std__lane14_strm1_ready         ( pe33__std__lane14_strm1_ready      ),      
               .std__pe33__lane14_strm1_cntl          ( std__pe33__lane14_strm1_cntl       ),      
               .std__pe33__lane14_strm1_data          ( std__pe33__lane14_strm1_data       ),      
               .std__pe33__lane14_strm1_data_valid    ( std__pe33__lane14_strm1_data_valid ),      
               .std__pe33__lane14_strm1_data_mask     ( std__pe33__lane14_strm1_data_mask  ),      

               // PE 33, Lane 15                 
               .pe33__std__lane15_strm0_ready         ( pe33__std__lane15_strm0_ready      ),      
               .std__pe33__lane15_strm0_cntl          ( std__pe33__lane15_strm0_cntl       ),      
               .std__pe33__lane15_strm0_data          ( std__pe33__lane15_strm0_data       ),      
               .std__pe33__lane15_strm0_data_valid    ( std__pe33__lane15_strm0_data_valid ),      
               .std__pe33__lane15_strm0_data_mask     ( std__pe33__lane15_strm0_data_mask  ),      

               .pe33__std__lane15_strm1_ready         ( pe33__std__lane15_strm1_ready      ),      
               .std__pe33__lane15_strm1_cntl          ( std__pe33__lane15_strm1_cntl       ),      
               .std__pe33__lane15_strm1_data          ( std__pe33__lane15_strm1_data       ),      
               .std__pe33__lane15_strm1_data_valid    ( std__pe33__lane15_strm1_data_valid ),      
               .std__pe33__lane15_strm1_data_mask     ( std__pe33__lane15_strm1_data_mask  ),      

               // PE 33, Lane 16                 
               .pe33__std__lane16_strm0_ready         ( pe33__std__lane16_strm0_ready      ),      
               .std__pe33__lane16_strm0_cntl          ( std__pe33__lane16_strm0_cntl       ),      
               .std__pe33__lane16_strm0_data          ( std__pe33__lane16_strm0_data       ),      
               .std__pe33__lane16_strm0_data_valid    ( std__pe33__lane16_strm0_data_valid ),      
               .std__pe33__lane16_strm0_data_mask     ( std__pe33__lane16_strm0_data_mask  ),      

               .pe33__std__lane16_strm1_ready         ( pe33__std__lane16_strm1_ready      ),      
               .std__pe33__lane16_strm1_cntl          ( std__pe33__lane16_strm1_cntl       ),      
               .std__pe33__lane16_strm1_data          ( std__pe33__lane16_strm1_data       ),      
               .std__pe33__lane16_strm1_data_valid    ( std__pe33__lane16_strm1_data_valid ),      
               .std__pe33__lane16_strm1_data_mask     ( std__pe33__lane16_strm1_data_mask  ),      

               // PE 33, Lane 17                 
               .pe33__std__lane17_strm0_ready         ( pe33__std__lane17_strm0_ready      ),      
               .std__pe33__lane17_strm0_cntl          ( std__pe33__lane17_strm0_cntl       ),      
               .std__pe33__lane17_strm0_data          ( std__pe33__lane17_strm0_data       ),      
               .std__pe33__lane17_strm0_data_valid    ( std__pe33__lane17_strm0_data_valid ),      
               .std__pe33__lane17_strm0_data_mask     ( std__pe33__lane17_strm0_data_mask  ),      

               .pe33__std__lane17_strm1_ready         ( pe33__std__lane17_strm1_ready      ),      
               .std__pe33__lane17_strm1_cntl          ( std__pe33__lane17_strm1_cntl       ),      
               .std__pe33__lane17_strm1_data          ( std__pe33__lane17_strm1_data       ),      
               .std__pe33__lane17_strm1_data_valid    ( std__pe33__lane17_strm1_data_valid ),      
               .std__pe33__lane17_strm1_data_mask     ( std__pe33__lane17_strm1_data_mask  ),      

               // PE 33, Lane 18                 
               .pe33__std__lane18_strm0_ready         ( pe33__std__lane18_strm0_ready      ),      
               .std__pe33__lane18_strm0_cntl          ( std__pe33__lane18_strm0_cntl       ),      
               .std__pe33__lane18_strm0_data          ( std__pe33__lane18_strm0_data       ),      
               .std__pe33__lane18_strm0_data_valid    ( std__pe33__lane18_strm0_data_valid ),      
               .std__pe33__lane18_strm0_data_mask     ( std__pe33__lane18_strm0_data_mask  ),      

               .pe33__std__lane18_strm1_ready         ( pe33__std__lane18_strm1_ready      ),      
               .std__pe33__lane18_strm1_cntl          ( std__pe33__lane18_strm1_cntl       ),      
               .std__pe33__lane18_strm1_data          ( std__pe33__lane18_strm1_data       ),      
               .std__pe33__lane18_strm1_data_valid    ( std__pe33__lane18_strm1_data_valid ),      
               .std__pe33__lane18_strm1_data_mask     ( std__pe33__lane18_strm1_data_mask  ),      

               // PE 33, Lane 19                 
               .pe33__std__lane19_strm0_ready         ( pe33__std__lane19_strm0_ready      ),      
               .std__pe33__lane19_strm0_cntl          ( std__pe33__lane19_strm0_cntl       ),      
               .std__pe33__lane19_strm0_data          ( std__pe33__lane19_strm0_data       ),      
               .std__pe33__lane19_strm0_data_valid    ( std__pe33__lane19_strm0_data_valid ),      
               .std__pe33__lane19_strm0_data_mask     ( std__pe33__lane19_strm0_data_mask  ),      

               .pe33__std__lane19_strm1_ready         ( pe33__std__lane19_strm1_ready      ),      
               .std__pe33__lane19_strm1_cntl          ( std__pe33__lane19_strm1_cntl       ),      
               .std__pe33__lane19_strm1_data          ( std__pe33__lane19_strm1_data       ),      
               .std__pe33__lane19_strm1_data_valid    ( std__pe33__lane19_strm1_data_valid ),      
               .std__pe33__lane19_strm1_data_mask     ( std__pe33__lane19_strm1_data_mask  ),      

               // PE 33, Lane 20                 
               .pe33__std__lane20_strm0_ready         ( pe33__std__lane20_strm0_ready      ),      
               .std__pe33__lane20_strm0_cntl          ( std__pe33__lane20_strm0_cntl       ),      
               .std__pe33__lane20_strm0_data          ( std__pe33__lane20_strm0_data       ),      
               .std__pe33__lane20_strm0_data_valid    ( std__pe33__lane20_strm0_data_valid ),      
               .std__pe33__lane20_strm0_data_mask     ( std__pe33__lane20_strm0_data_mask  ),      

               .pe33__std__lane20_strm1_ready         ( pe33__std__lane20_strm1_ready      ),      
               .std__pe33__lane20_strm1_cntl          ( std__pe33__lane20_strm1_cntl       ),      
               .std__pe33__lane20_strm1_data          ( std__pe33__lane20_strm1_data       ),      
               .std__pe33__lane20_strm1_data_valid    ( std__pe33__lane20_strm1_data_valid ),      
               .std__pe33__lane20_strm1_data_mask     ( std__pe33__lane20_strm1_data_mask  ),      

               // PE 33, Lane 21                 
               .pe33__std__lane21_strm0_ready         ( pe33__std__lane21_strm0_ready      ),      
               .std__pe33__lane21_strm0_cntl          ( std__pe33__lane21_strm0_cntl       ),      
               .std__pe33__lane21_strm0_data          ( std__pe33__lane21_strm0_data       ),      
               .std__pe33__lane21_strm0_data_valid    ( std__pe33__lane21_strm0_data_valid ),      
               .std__pe33__lane21_strm0_data_mask     ( std__pe33__lane21_strm0_data_mask  ),      

               .pe33__std__lane21_strm1_ready         ( pe33__std__lane21_strm1_ready      ),      
               .std__pe33__lane21_strm1_cntl          ( std__pe33__lane21_strm1_cntl       ),      
               .std__pe33__lane21_strm1_data          ( std__pe33__lane21_strm1_data       ),      
               .std__pe33__lane21_strm1_data_valid    ( std__pe33__lane21_strm1_data_valid ),      
               .std__pe33__lane21_strm1_data_mask     ( std__pe33__lane21_strm1_data_mask  ),      

               // PE 33, Lane 22                 
               .pe33__std__lane22_strm0_ready         ( pe33__std__lane22_strm0_ready      ),      
               .std__pe33__lane22_strm0_cntl          ( std__pe33__lane22_strm0_cntl       ),      
               .std__pe33__lane22_strm0_data          ( std__pe33__lane22_strm0_data       ),      
               .std__pe33__lane22_strm0_data_valid    ( std__pe33__lane22_strm0_data_valid ),      
               .std__pe33__lane22_strm0_data_mask     ( std__pe33__lane22_strm0_data_mask  ),      

               .pe33__std__lane22_strm1_ready         ( pe33__std__lane22_strm1_ready      ),      
               .std__pe33__lane22_strm1_cntl          ( std__pe33__lane22_strm1_cntl       ),      
               .std__pe33__lane22_strm1_data          ( std__pe33__lane22_strm1_data       ),      
               .std__pe33__lane22_strm1_data_valid    ( std__pe33__lane22_strm1_data_valid ),      
               .std__pe33__lane22_strm1_data_mask     ( std__pe33__lane22_strm1_data_mask  ),      

               // PE 33, Lane 23                 
               .pe33__std__lane23_strm0_ready         ( pe33__std__lane23_strm0_ready      ),      
               .std__pe33__lane23_strm0_cntl          ( std__pe33__lane23_strm0_cntl       ),      
               .std__pe33__lane23_strm0_data          ( std__pe33__lane23_strm0_data       ),      
               .std__pe33__lane23_strm0_data_valid    ( std__pe33__lane23_strm0_data_valid ),      
               .std__pe33__lane23_strm0_data_mask     ( std__pe33__lane23_strm0_data_mask  ),      

               .pe33__std__lane23_strm1_ready         ( pe33__std__lane23_strm1_ready      ),      
               .std__pe33__lane23_strm1_cntl          ( std__pe33__lane23_strm1_cntl       ),      
               .std__pe33__lane23_strm1_data          ( std__pe33__lane23_strm1_data       ),      
               .std__pe33__lane23_strm1_data_valid    ( std__pe33__lane23_strm1_data_valid ),      
               .std__pe33__lane23_strm1_data_mask     ( std__pe33__lane23_strm1_data_mask  ),      

               // PE 33, Lane 24                 
               .pe33__std__lane24_strm0_ready         ( pe33__std__lane24_strm0_ready      ),      
               .std__pe33__lane24_strm0_cntl          ( std__pe33__lane24_strm0_cntl       ),      
               .std__pe33__lane24_strm0_data          ( std__pe33__lane24_strm0_data       ),      
               .std__pe33__lane24_strm0_data_valid    ( std__pe33__lane24_strm0_data_valid ),      
               .std__pe33__lane24_strm0_data_mask     ( std__pe33__lane24_strm0_data_mask  ),      

               .pe33__std__lane24_strm1_ready         ( pe33__std__lane24_strm1_ready      ),      
               .std__pe33__lane24_strm1_cntl          ( std__pe33__lane24_strm1_cntl       ),      
               .std__pe33__lane24_strm1_data          ( std__pe33__lane24_strm1_data       ),      
               .std__pe33__lane24_strm1_data_valid    ( std__pe33__lane24_strm1_data_valid ),      
               .std__pe33__lane24_strm1_data_mask     ( std__pe33__lane24_strm1_data_mask  ),      

               // PE 33, Lane 25                 
               .pe33__std__lane25_strm0_ready         ( pe33__std__lane25_strm0_ready      ),      
               .std__pe33__lane25_strm0_cntl          ( std__pe33__lane25_strm0_cntl       ),      
               .std__pe33__lane25_strm0_data          ( std__pe33__lane25_strm0_data       ),      
               .std__pe33__lane25_strm0_data_valid    ( std__pe33__lane25_strm0_data_valid ),      
               .std__pe33__lane25_strm0_data_mask     ( std__pe33__lane25_strm0_data_mask  ),      

               .pe33__std__lane25_strm1_ready         ( pe33__std__lane25_strm1_ready      ),      
               .std__pe33__lane25_strm1_cntl          ( std__pe33__lane25_strm1_cntl       ),      
               .std__pe33__lane25_strm1_data          ( std__pe33__lane25_strm1_data       ),      
               .std__pe33__lane25_strm1_data_valid    ( std__pe33__lane25_strm1_data_valid ),      
               .std__pe33__lane25_strm1_data_mask     ( std__pe33__lane25_strm1_data_mask  ),      

               // PE 33, Lane 26                 
               .pe33__std__lane26_strm0_ready         ( pe33__std__lane26_strm0_ready      ),      
               .std__pe33__lane26_strm0_cntl          ( std__pe33__lane26_strm0_cntl       ),      
               .std__pe33__lane26_strm0_data          ( std__pe33__lane26_strm0_data       ),      
               .std__pe33__lane26_strm0_data_valid    ( std__pe33__lane26_strm0_data_valid ),      
               .std__pe33__lane26_strm0_data_mask     ( std__pe33__lane26_strm0_data_mask  ),      

               .pe33__std__lane26_strm1_ready         ( pe33__std__lane26_strm1_ready      ),      
               .std__pe33__lane26_strm1_cntl          ( std__pe33__lane26_strm1_cntl       ),      
               .std__pe33__lane26_strm1_data          ( std__pe33__lane26_strm1_data       ),      
               .std__pe33__lane26_strm1_data_valid    ( std__pe33__lane26_strm1_data_valid ),      
               .std__pe33__lane26_strm1_data_mask     ( std__pe33__lane26_strm1_data_mask  ),      

               // PE 33, Lane 27                 
               .pe33__std__lane27_strm0_ready         ( pe33__std__lane27_strm0_ready      ),      
               .std__pe33__lane27_strm0_cntl          ( std__pe33__lane27_strm0_cntl       ),      
               .std__pe33__lane27_strm0_data          ( std__pe33__lane27_strm0_data       ),      
               .std__pe33__lane27_strm0_data_valid    ( std__pe33__lane27_strm0_data_valid ),      
               .std__pe33__lane27_strm0_data_mask     ( std__pe33__lane27_strm0_data_mask  ),      

               .pe33__std__lane27_strm1_ready         ( pe33__std__lane27_strm1_ready      ),      
               .std__pe33__lane27_strm1_cntl          ( std__pe33__lane27_strm1_cntl       ),      
               .std__pe33__lane27_strm1_data          ( std__pe33__lane27_strm1_data       ),      
               .std__pe33__lane27_strm1_data_valid    ( std__pe33__lane27_strm1_data_valid ),      
               .std__pe33__lane27_strm1_data_mask     ( std__pe33__lane27_strm1_data_mask  ),      

               // PE 33, Lane 28                 
               .pe33__std__lane28_strm0_ready         ( pe33__std__lane28_strm0_ready      ),      
               .std__pe33__lane28_strm0_cntl          ( std__pe33__lane28_strm0_cntl       ),      
               .std__pe33__lane28_strm0_data          ( std__pe33__lane28_strm0_data       ),      
               .std__pe33__lane28_strm0_data_valid    ( std__pe33__lane28_strm0_data_valid ),      
               .std__pe33__lane28_strm0_data_mask     ( std__pe33__lane28_strm0_data_mask  ),      

               .pe33__std__lane28_strm1_ready         ( pe33__std__lane28_strm1_ready      ),      
               .std__pe33__lane28_strm1_cntl          ( std__pe33__lane28_strm1_cntl       ),      
               .std__pe33__lane28_strm1_data          ( std__pe33__lane28_strm1_data       ),      
               .std__pe33__lane28_strm1_data_valid    ( std__pe33__lane28_strm1_data_valid ),      
               .std__pe33__lane28_strm1_data_mask     ( std__pe33__lane28_strm1_data_mask  ),      

               // PE 33, Lane 29                 
               .pe33__std__lane29_strm0_ready         ( pe33__std__lane29_strm0_ready      ),      
               .std__pe33__lane29_strm0_cntl          ( std__pe33__lane29_strm0_cntl       ),      
               .std__pe33__lane29_strm0_data          ( std__pe33__lane29_strm0_data       ),      
               .std__pe33__lane29_strm0_data_valid    ( std__pe33__lane29_strm0_data_valid ),      
               .std__pe33__lane29_strm0_data_mask     ( std__pe33__lane29_strm0_data_mask  ),      

               .pe33__std__lane29_strm1_ready         ( pe33__std__lane29_strm1_ready      ),      
               .std__pe33__lane29_strm1_cntl          ( std__pe33__lane29_strm1_cntl       ),      
               .std__pe33__lane29_strm1_data          ( std__pe33__lane29_strm1_data       ),      
               .std__pe33__lane29_strm1_data_valid    ( std__pe33__lane29_strm1_data_valid ),      
               .std__pe33__lane29_strm1_data_mask     ( std__pe33__lane29_strm1_data_mask  ),      

               // PE 33, Lane 30                 
               .pe33__std__lane30_strm0_ready         ( pe33__std__lane30_strm0_ready      ),      
               .std__pe33__lane30_strm0_cntl          ( std__pe33__lane30_strm0_cntl       ),      
               .std__pe33__lane30_strm0_data          ( std__pe33__lane30_strm0_data       ),      
               .std__pe33__lane30_strm0_data_valid    ( std__pe33__lane30_strm0_data_valid ),      
               .std__pe33__lane30_strm0_data_mask     ( std__pe33__lane30_strm0_data_mask  ),      

               .pe33__std__lane30_strm1_ready         ( pe33__std__lane30_strm1_ready      ),      
               .std__pe33__lane30_strm1_cntl          ( std__pe33__lane30_strm1_cntl       ),      
               .std__pe33__lane30_strm1_data          ( std__pe33__lane30_strm1_data       ),      
               .std__pe33__lane30_strm1_data_valid    ( std__pe33__lane30_strm1_data_valid ),      
               .std__pe33__lane30_strm1_data_mask     ( std__pe33__lane30_strm1_data_mask  ),      

               // PE 33, Lane 31                 
               .pe33__std__lane31_strm0_ready         ( pe33__std__lane31_strm0_ready      ),      
               .std__pe33__lane31_strm0_cntl          ( std__pe33__lane31_strm0_cntl       ),      
               .std__pe33__lane31_strm0_data          ( std__pe33__lane31_strm0_data       ),      
               .std__pe33__lane31_strm0_data_valid    ( std__pe33__lane31_strm0_data_valid ),      
               .std__pe33__lane31_strm0_data_mask     ( std__pe33__lane31_strm0_data_mask  ),      

               .pe33__std__lane31_strm1_ready         ( pe33__std__lane31_strm1_ready      ),      
               .std__pe33__lane31_strm1_cntl          ( std__pe33__lane31_strm1_cntl       ),      
               .std__pe33__lane31_strm1_data          ( std__pe33__lane31_strm1_data       ),      
               .std__pe33__lane31_strm1_data_valid    ( std__pe33__lane31_strm1_data_valid ),      
               .std__pe33__lane31_strm1_data_mask     ( std__pe33__lane31_strm1_data_mask  ),      

               // PE 34, Lane 0                 
               .pe34__std__lane0_strm0_ready         ( pe34__std__lane0_strm0_ready      ),      
               .std__pe34__lane0_strm0_cntl          ( std__pe34__lane0_strm0_cntl       ),      
               .std__pe34__lane0_strm0_data          ( std__pe34__lane0_strm0_data       ),      
               .std__pe34__lane0_strm0_data_valid    ( std__pe34__lane0_strm0_data_valid ),      
               .std__pe34__lane0_strm0_data_mask     ( std__pe34__lane0_strm0_data_mask  ),      

               .pe34__std__lane0_strm1_ready         ( pe34__std__lane0_strm1_ready      ),      
               .std__pe34__lane0_strm1_cntl          ( std__pe34__lane0_strm1_cntl       ),      
               .std__pe34__lane0_strm1_data          ( std__pe34__lane0_strm1_data       ),      
               .std__pe34__lane0_strm1_data_valid    ( std__pe34__lane0_strm1_data_valid ),      
               .std__pe34__lane0_strm1_data_mask     ( std__pe34__lane0_strm1_data_mask  ),      

               // PE 34, Lane 1                 
               .pe34__std__lane1_strm0_ready         ( pe34__std__lane1_strm0_ready      ),      
               .std__pe34__lane1_strm0_cntl          ( std__pe34__lane1_strm0_cntl       ),      
               .std__pe34__lane1_strm0_data          ( std__pe34__lane1_strm0_data       ),      
               .std__pe34__lane1_strm0_data_valid    ( std__pe34__lane1_strm0_data_valid ),      
               .std__pe34__lane1_strm0_data_mask     ( std__pe34__lane1_strm0_data_mask  ),      

               .pe34__std__lane1_strm1_ready         ( pe34__std__lane1_strm1_ready      ),      
               .std__pe34__lane1_strm1_cntl          ( std__pe34__lane1_strm1_cntl       ),      
               .std__pe34__lane1_strm1_data          ( std__pe34__lane1_strm1_data       ),      
               .std__pe34__lane1_strm1_data_valid    ( std__pe34__lane1_strm1_data_valid ),      
               .std__pe34__lane1_strm1_data_mask     ( std__pe34__lane1_strm1_data_mask  ),      

               // PE 34, Lane 2                 
               .pe34__std__lane2_strm0_ready         ( pe34__std__lane2_strm0_ready      ),      
               .std__pe34__lane2_strm0_cntl          ( std__pe34__lane2_strm0_cntl       ),      
               .std__pe34__lane2_strm0_data          ( std__pe34__lane2_strm0_data       ),      
               .std__pe34__lane2_strm0_data_valid    ( std__pe34__lane2_strm0_data_valid ),      
               .std__pe34__lane2_strm0_data_mask     ( std__pe34__lane2_strm0_data_mask  ),      

               .pe34__std__lane2_strm1_ready         ( pe34__std__lane2_strm1_ready      ),      
               .std__pe34__lane2_strm1_cntl          ( std__pe34__lane2_strm1_cntl       ),      
               .std__pe34__lane2_strm1_data          ( std__pe34__lane2_strm1_data       ),      
               .std__pe34__lane2_strm1_data_valid    ( std__pe34__lane2_strm1_data_valid ),      
               .std__pe34__lane2_strm1_data_mask     ( std__pe34__lane2_strm1_data_mask  ),      

               // PE 34, Lane 3                 
               .pe34__std__lane3_strm0_ready         ( pe34__std__lane3_strm0_ready      ),      
               .std__pe34__lane3_strm0_cntl          ( std__pe34__lane3_strm0_cntl       ),      
               .std__pe34__lane3_strm0_data          ( std__pe34__lane3_strm0_data       ),      
               .std__pe34__lane3_strm0_data_valid    ( std__pe34__lane3_strm0_data_valid ),      
               .std__pe34__lane3_strm0_data_mask     ( std__pe34__lane3_strm0_data_mask  ),      

               .pe34__std__lane3_strm1_ready         ( pe34__std__lane3_strm1_ready      ),      
               .std__pe34__lane3_strm1_cntl          ( std__pe34__lane3_strm1_cntl       ),      
               .std__pe34__lane3_strm1_data          ( std__pe34__lane3_strm1_data       ),      
               .std__pe34__lane3_strm1_data_valid    ( std__pe34__lane3_strm1_data_valid ),      
               .std__pe34__lane3_strm1_data_mask     ( std__pe34__lane3_strm1_data_mask  ),      

               // PE 34, Lane 4                 
               .pe34__std__lane4_strm0_ready         ( pe34__std__lane4_strm0_ready      ),      
               .std__pe34__lane4_strm0_cntl          ( std__pe34__lane4_strm0_cntl       ),      
               .std__pe34__lane4_strm0_data          ( std__pe34__lane4_strm0_data       ),      
               .std__pe34__lane4_strm0_data_valid    ( std__pe34__lane4_strm0_data_valid ),      
               .std__pe34__lane4_strm0_data_mask     ( std__pe34__lane4_strm0_data_mask  ),      

               .pe34__std__lane4_strm1_ready         ( pe34__std__lane4_strm1_ready      ),      
               .std__pe34__lane4_strm1_cntl          ( std__pe34__lane4_strm1_cntl       ),      
               .std__pe34__lane4_strm1_data          ( std__pe34__lane4_strm1_data       ),      
               .std__pe34__lane4_strm1_data_valid    ( std__pe34__lane4_strm1_data_valid ),      
               .std__pe34__lane4_strm1_data_mask     ( std__pe34__lane4_strm1_data_mask  ),      

               // PE 34, Lane 5                 
               .pe34__std__lane5_strm0_ready         ( pe34__std__lane5_strm0_ready      ),      
               .std__pe34__lane5_strm0_cntl          ( std__pe34__lane5_strm0_cntl       ),      
               .std__pe34__lane5_strm0_data          ( std__pe34__lane5_strm0_data       ),      
               .std__pe34__lane5_strm0_data_valid    ( std__pe34__lane5_strm0_data_valid ),      
               .std__pe34__lane5_strm0_data_mask     ( std__pe34__lane5_strm0_data_mask  ),      

               .pe34__std__lane5_strm1_ready         ( pe34__std__lane5_strm1_ready      ),      
               .std__pe34__lane5_strm1_cntl          ( std__pe34__lane5_strm1_cntl       ),      
               .std__pe34__lane5_strm1_data          ( std__pe34__lane5_strm1_data       ),      
               .std__pe34__lane5_strm1_data_valid    ( std__pe34__lane5_strm1_data_valid ),      
               .std__pe34__lane5_strm1_data_mask     ( std__pe34__lane5_strm1_data_mask  ),      

               // PE 34, Lane 6                 
               .pe34__std__lane6_strm0_ready         ( pe34__std__lane6_strm0_ready      ),      
               .std__pe34__lane6_strm0_cntl          ( std__pe34__lane6_strm0_cntl       ),      
               .std__pe34__lane6_strm0_data          ( std__pe34__lane6_strm0_data       ),      
               .std__pe34__lane6_strm0_data_valid    ( std__pe34__lane6_strm0_data_valid ),      
               .std__pe34__lane6_strm0_data_mask     ( std__pe34__lane6_strm0_data_mask  ),      

               .pe34__std__lane6_strm1_ready         ( pe34__std__lane6_strm1_ready      ),      
               .std__pe34__lane6_strm1_cntl          ( std__pe34__lane6_strm1_cntl       ),      
               .std__pe34__lane6_strm1_data          ( std__pe34__lane6_strm1_data       ),      
               .std__pe34__lane6_strm1_data_valid    ( std__pe34__lane6_strm1_data_valid ),      
               .std__pe34__lane6_strm1_data_mask     ( std__pe34__lane6_strm1_data_mask  ),      

               // PE 34, Lane 7                 
               .pe34__std__lane7_strm0_ready         ( pe34__std__lane7_strm0_ready      ),      
               .std__pe34__lane7_strm0_cntl          ( std__pe34__lane7_strm0_cntl       ),      
               .std__pe34__lane7_strm0_data          ( std__pe34__lane7_strm0_data       ),      
               .std__pe34__lane7_strm0_data_valid    ( std__pe34__lane7_strm0_data_valid ),      
               .std__pe34__lane7_strm0_data_mask     ( std__pe34__lane7_strm0_data_mask  ),      

               .pe34__std__lane7_strm1_ready         ( pe34__std__lane7_strm1_ready      ),      
               .std__pe34__lane7_strm1_cntl          ( std__pe34__lane7_strm1_cntl       ),      
               .std__pe34__lane7_strm1_data          ( std__pe34__lane7_strm1_data       ),      
               .std__pe34__lane7_strm1_data_valid    ( std__pe34__lane7_strm1_data_valid ),      
               .std__pe34__lane7_strm1_data_mask     ( std__pe34__lane7_strm1_data_mask  ),      

               // PE 34, Lane 8                 
               .pe34__std__lane8_strm0_ready         ( pe34__std__lane8_strm0_ready      ),      
               .std__pe34__lane8_strm0_cntl          ( std__pe34__lane8_strm0_cntl       ),      
               .std__pe34__lane8_strm0_data          ( std__pe34__lane8_strm0_data       ),      
               .std__pe34__lane8_strm0_data_valid    ( std__pe34__lane8_strm0_data_valid ),      
               .std__pe34__lane8_strm0_data_mask     ( std__pe34__lane8_strm0_data_mask  ),      

               .pe34__std__lane8_strm1_ready         ( pe34__std__lane8_strm1_ready      ),      
               .std__pe34__lane8_strm1_cntl          ( std__pe34__lane8_strm1_cntl       ),      
               .std__pe34__lane8_strm1_data          ( std__pe34__lane8_strm1_data       ),      
               .std__pe34__lane8_strm1_data_valid    ( std__pe34__lane8_strm1_data_valid ),      
               .std__pe34__lane8_strm1_data_mask     ( std__pe34__lane8_strm1_data_mask  ),      

               // PE 34, Lane 9                 
               .pe34__std__lane9_strm0_ready         ( pe34__std__lane9_strm0_ready      ),      
               .std__pe34__lane9_strm0_cntl          ( std__pe34__lane9_strm0_cntl       ),      
               .std__pe34__lane9_strm0_data          ( std__pe34__lane9_strm0_data       ),      
               .std__pe34__lane9_strm0_data_valid    ( std__pe34__lane9_strm0_data_valid ),      
               .std__pe34__lane9_strm0_data_mask     ( std__pe34__lane9_strm0_data_mask  ),      

               .pe34__std__lane9_strm1_ready         ( pe34__std__lane9_strm1_ready      ),      
               .std__pe34__lane9_strm1_cntl          ( std__pe34__lane9_strm1_cntl       ),      
               .std__pe34__lane9_strm1_data          ( std__pe34__lane9_strm1_data       ),      
               .std__pe34__lane9_strm1_data_valid    ( std__pe34__lane9_strm1_data_valid ),      
               .std__pe34__lane9_strm1_data_mask     ( std__pe34__lane9_strm1_data_mask  ),      

               // PE 34, Lane 10                 
               .pe34__std__lane10_strm0_ready         ( pe34__std__lane10_strm0_ready      ),      
               .std__pe34__lane10_strm0_cntl          ( std__pe34__lane10_strm0_cntl       ),      
               .std__pe34__lane10_strm0_data          ( std__pe34__lane10_strm0_data       ),      
               .std__pe34__lane10_strm0_data_valid    ( std__pe34__lane10_strm0_data_valid ),      
               .std__pe34__lane10_strm0_data_mask     ( std__pe34__lane10_strm0_data_mask  ),      

               .pe34__std__lane10_strm1_ready         ( pe34__std__lane10_strm1_ready      ),      
               .std__pe34__lane10_strm1_cntl          ( std__pe34__lane10_strm1_cntl       ),      
               .std__pe34__lane10_strm1_data          ( std__pe34__lane10_strm1_data       ),      
               .std__pe34__lane10_strm1_data_valid    ( std__pe34__lane10_strm1_data_valid ),      
               .std__pe34__lane10_strm1_data_mask     ( std__pe34__lane10_strm1_data_mask  ),      

               // PE 34, Lane 11                 
               .pe34__std__lane11_strm0_ready         ( pe34__std__lane11_strm0_ready      ),      
               .std__pe34__lane11_strm0_cntl          ( std__pe34__lane11_strm0_cntl       ),      
               .std__pe34__lane11_strm0_data          ( std__pe34__lane11_strm0_data       ),      
               .std__pe34__lane11_strm0_data_valid    ( std__pe34__lane11_strm0_data_valid ),      
               .std__pe34__lane11_strm0_data_mask     ( std__pe34__lane11_strm0_data_mask  ),      

               .pe34__std__lane11_strm1_ready         ( pe34__std__lane11_strm1_ready      ),      
               .std__pe34__lane11_strm1_cntl          ( std__pe34__lane11_strm1_cntl       ),      
               .std__pe34__lane11_strm1_data          ( std__pe34__lane11_strm1_data       ),      
               .std__pe34__lane11_strm1_data_valid    ( std__pe34__lane11_strm1_data_valid ),      
               .std__pe34__lane11_strm1_data_mask     ( std__pe34__lane11_strm1_data_mask  ),      

               // PE 34, Lane 12                 
               .pe34__std__lane12_strm0_ready         ( pe34__std__lane12_strm0_ready      ),      
               .std__pe34__lane12_strm0_cntl          ( std__pe34__lane12_strm0_cntl       ),      
               .std__pe34__lane12_strm0_data          ( std__pe34__lane12_strm0_data       ),      
               .std__pe34__lane12_strm0_data_valid    ( std__pe34__lane12_strm0_data_valid ),      
               .std__pe34__lane12_strm0_data_mask     ( std__pe34__lane12_strm0_data_mask  ),      

               .pe34__std__lane12_strm1_ready         ( pe34__std__lane12_strm1_ready      ),      
               .std__pe34__lane12_strm1_cntl          ( std__pe34__lane12_strm1_cntl       ),      
               .std__pe34__lane12_strm1_data          ( std__pe34__lane12_strm1_data       ),      
               .std__pe34__lane12_strm1_data_valid    ( std__pe34__lane12_strm1_data_valid ),      
               .std__pe34__lane12_strm1_data_mask     ( std__pe34__lane12_strm1_data_mask  ),      

               // PE 34, Lane 13                 
               .pe34__std__lane13_strm0_ready         ( pe34__std__lane13_strm0_ready      ),      
               .std__pe34__lane13_strm0_cntl          ( std__pe34__lane13_strm0_cntl       ),      
               .std__pe34__lane13_strm0_data          ( std__pe34__lane13_strm0_data       ),      
               .std__pe34__lane13_strm0_data_valid    ( std__pe34__lane13_strm0_data_valid ),      
               .std__pe34__lane13_strm0_data_mask     ( std__pe34__lane13_strm0_data_mask  ),      

               .pe34__std__lane13_strm1_ready         ( pe34__std__lane13_strm1_ready      ),      
               .std__pe34__lane13_strm1_cntl          ( std__pe34__lane13_strm1_cntl       ),      
               .std__pe34__lane13_strm1_data          ( std__pe34__lane13_strm1_data       ),      
               .std__pe34__lane13_strm1_data_valid    ( std__pe34__lane13_strm1_data_valid ),      
               .std__pe34__lane13_strm1_data_mask     ( std__pe34__lane13_strm1_data_mask  ),      

               // PE 34, Lane 14                 
               .pe34__std__lane14_strm0_ready         ( pe34__std__lane14_strm0_ready      ),      
               .std__pe34__lane14_strm0_cntl          ( std__pe34__lane14_strm0_cntl       ),      
               .std__pe34__lane14_strm0_data          ( std__pe34__lane14_strm0_data       ),      
               .std__pe34__lane14_strm0_data_valid    ( std__pe34__lane14_strm0_data_valid ),      
               .std__pe34__lane14_strm0_data_mask     ( std__pe34__lane14_strm0_data_mask  ),      

               .pe34__std__lane14_strm1_ready         ( pe34__std__lane14_strm1_ready      ),      
               .std__pe34__lane14_strm1_cntl          ( std__pe34__lane14_strm1_cntl       ),      
               .std__pe34__lane14_strm1_data          ( std__pe34__lane14_strm1_data       ),      
               .std__pe34__lane14_strm1_data_valid    ( std__pe34__lane14_strm1_data_valid ),      
               .std__pe34__lane14_strm1_data_mask     ( std__pe34__lane14_strm1_data_mask  ),      

               // PE 34, Lane 15                 
               .pe34__std__lane15_strm0_ready         ( pe34__std__lane15_strm0_ready      ),      
               .std__pe34__lane15_strm0_cntl          ( std__pe34__lane15_strm0_cntl       ),      
               .std__pe34__lane15_strm0_data          ( std__pe34__lane15_strm0_data       ),      
               .std__pe34__lane15_strm0_data_valid    ( std__pe34__lane15_strm0_data_valid ),      
               .std__pe34__lane15_strm0_data_mask     ( std__pe34__lane15_strm0_data_mask  ),      

               .pe34__std__lane15_strm1_ready         ( pe34__std__lane15_strm1_ready      ),      
               .std__pe34__lane15_strm1_cntl          ( std__pe34__lane15_strm1_cntl       ),      
               .std__pe34__lane15_strm1_data          ( std__pe34__lane15_strm1_data       ),      
               .std__pe34__lane15_strm1_data_valid    ( std__pe34__lane15_strm1_data_valid ),      
               .std__pe34__lane15_strm1_data_mask     ( std__pe34__lane15_strm1_data_mask  ),      

               // PE 34, Lane 16                 
               .pe34__std__lane16_strm0_ready         ( pe34__std__lane16_strm0_ready      ),      
               .std__pe34__lane16_strm0_cntl          ( std__pe34__lane16_strm0_cntl       ),      
               .std__pe34__lane16_strm0_data          ( std__pe34__lane16_strm0_data       ),      
               .std__pe34__lane16_strm0_data_valid    ( std__pe34__lane16_strm0_data_valid ),      
               .std__pe34__lane16_strm0_data_mask     ( std__pe34__lane16_strm0_data_mask  ),      

               .pe34__std__lane16_strm1_ready         ( pe34__std__lane16_strm1_ready      ),      
               .std__pe34__lane16_strm1_cntl          ( std__pe34__lane16_strm1_cntl       ),      
               .std__pe34__lane16_strm1_data          ( std__pe34__lane16_strm1_data       ),      
               .std__pe34__lane16_strm1_data_valid    ( std__pe34__lane16_strm1_data_valid ),      
               .std__pe34__lane16_strm1_data_mask     ( std__pe34__lane16_strm1_data_mask  ),      

               // PE 34, Lane 17                 
               .pe34__std__lane17_strm0_ready         ( pe34__std__lane17_strm0_ready      ),      
               .std__pe34__lane17_strm0_cntl          ( std__pe34__lane17_strm0_cntl       ),      
               .std__pe34__lane17_strm0_data          ( std__pe34__lane17_strm0_data       ),      
               .std__pe34__lane17_strm0_data_valid    ( std__pe34__lane17_strm0_data_valid ),      
               .std__pe34__lane17_strm0_data_mask     ( std__pe34__lane17_strm0_data_mask  ),      

               .pe34__std__lane17_strm1_ready         ( pe34__std__lane17_strm1_ready      ),      
               .std__pe34__lane17_strm1_cntl          ( std__pe34__lane17_strm1_cntl       ),      
               .std__pe34__lane17_strm1_data          ( std__pe34__lane17_strm1_data       ),      
               .std__pe34__lane17_strm1_data_valid    ( std__pe34__lane17_strm1_data_valid ),      
               .std__pe34__lane17_strm1_data_mask     ( std__pe34__lane17_strm1_data_mask  ),      

               // PE 34, Lane 18                 
               .pe34__std__lane18_strm0_ready         ( pe34__std__lane18_strm0_ready      ),      
               .std__pe34__lane18_strm0_cntl          ( std__pe34__lane18_strm0_cntl       ),      
               .std__pe34__lane18_strm0_data          ( std__pe34__lane18_strm0_data       ),      
               .std__pe34__lane18_strm0_data_valid    ( std__pe34__lane18_strm0_data_valid ),      
               .std__pe34__lane18_strm0_data_mask     ( std__pe34__lane18_strm0_data_mask  ),      

               .pe34__std__lane18_strm1_ready         ( pe34__std__lane18_strm1_ready      ),      
               .std__pe34__lane18_strm1_cntl          ( std__pe34__lane18_strm1_cntl       ),      
               .std__pe34__lane18_strm1_data          ( std__pe34__lane18_strm1_data       ),      
               .std__pe34__lane18_strm1_data_valid    ( std__pe34__lane18_strm1_data_valid ),      
               .std__pe34__lane18_strm1_data_mask     ( std__pe34__lane18_strm1_data_mask  ),      

               // PE 34, Lane 19                 
               .pe34__std__lane19_strm0_ready         ( pe34__std__lane19_strm0_ready      ),      
               .std__pe34__lane19_strm0_cntl          ( std__pe34__lane19_strm0_cntl       ),      
               .std__pe34__lane19_strm0_data          ( std__pe34__lane19_strm0_data       ),      
               .std__pe34__lane19_strm0_data_valid    ( std__pe34__lane19_strm0_data_valid ),      
               .std__pe34__lane19_strm0_data_mask     ( std__pe34__lane19_strm0_data_mask  ),      

               .pe34__std__lane19_strm1_ready         ( pe34__std__lane19_strm1_ready      ),      
               .std__pe34__lane19_strm1_cntl          ( std__pe34__lane19_strm1_cntl       ),      
               .std__pe34__lane19_strm1_data          ( std__pe34__lane19_strm1_data       ),      
               .std__pe34__lane19_strm1_data_valid    ( std__pe34__lane19_strm1_data_valid ),      
               .std__pe34__lane19_strm1_data_mask     ( std__pe34__lane19_strm1_data_mask  ),      

               // PE 34, Lane 20                 
               .pe34__std__lane20_strm0_ready         ( pe34__std__lane20_strm0_ready      ),      
               .std__pe34__lane20_strm0_cntl          ( std__pe34__lane20_strm0_cntl       ),      
               .std__pe34__lane20_strm0_data          ( std__pe34__lane20_strm0_data       ),      
               .std__pe34__lane20_strm0_data_valid    ( std__pe34__lane20_strm0_data_valid ),      
               .std__pe34__lane20_strm0_data_mask     ( std__pe34__lane20_strm0_data_mask  ),      

               .pe34__std__lane20_strm1_ready         ( pe34__std__lane20_strm1_ready      ),      
               .std__pe34__lane20_strm1_cntl          ( std__pe34__lane20_strm1_cntl       ),      
               .std__pe34__lane20_strm1_data          ( std__pe34__lane20_strm1_data       ),      
               .std__pe34__lane20_strm1_data_valid    ( std__pe34__lane20_strm1_data_valid ),      
               .std__pe34__lane20_strm1_data_mask     ( std__pe34__lane20_strm1_data_mask  ),      

               // PE 34, Lane 21                 
               .pe34__std__lane21_strm0_ready         ( pe34__std__lane21_strm0_ready      ),      
               .std__pe34__lane21_strm0_cntl          ( std__pe34__lane21_strm0_cntl       ),      
               .std__pe34__lane21_strm0_data          ( std__pe34__lane21_strm0_data       ),      
               .std__pe34__lane21_strm0_data_valid    ( std__pe34__lane21_strm0_data_valid ),      
               .std__pe34__lane21_strm0_data_mask     ( std__pe34__lane21_strm0_data_mask  ),      

               .pe34__std__lane21_strm1_ready         ( pe34__std__lane21_strm1_ready      ),      
               .std__pe34__lane21_strm1_cntl          ( std__pe34__lane21_strm1_cntl       ),      
               .std__pe34__lane21_strm1_data          ( std__pe34__lane21_strm1_data       ),      
               .std__pe34__lane21_strm1_data_valid    ( std__pe34__lane21_strm1_data_valid ),      
               .std__pe34__lane21_strm1_data_mask     ( std__pe34__lane21_strm1_data_mask  ),      

               // PE 34, Lane 22                 
               .pe34__std__lane22_strm0_ready         ( pe34__std__lane22_strm0_ready      ),      
               .std__pe34__lane22_strm0_cntl          ( std__pe34__lane22_strm0_cntl       ),      
               .std__pe34__lane22_strm0_data          ( std__pe34__lane22_strm0_data       ),      
               .std__pe34__lane22_strm0_data_valid    ( std__pe34__lane22_strm0_data_valid ),      
               .std__pe34__lane22_strm0_data_mask     ( std__pe34__lane22_strm0_data_mask  ),      

               .pe34__std__lane22_strm1_ready         ( pe34__std__lane22_strm1_ready      ),      
               .std__pe34__lane22_strm1_cntl          ( std__pe34__lane22_strm1_cntl       ),      
               .std__pe34__lane22_strm1_data          ( std__pe34__lane22_strm1_data       ),      
               .std__pe34__lane22_strm1_data_valid    ( std__pe34__lane22_strm1_data_valid ),      
               .std__pe34__lane22_strm1_data_mask     ( std__pe34__lane22_strm1_data_mask  ),      

               // PE 34, Lane 23                 
               .pe34__std__lane23_strm0_ready         ( pe34__std__lane23_strm0_ready      ),      
               .std__pe34__lane23_strm0_cntl          ( std__pe34__lane23_strm0_cntl       ),      
               .std__pe34__lane23_strm0_data          ( std__pe34__lane23_strm0_data       ),      
               .std__pe34__lane23_strm0_data_valid    ( std__pe34__lane23_strm0_data_valid ),      
               .std__pe34__lane23_strm0_data_mask     ( std__pe34__lane23_strm0_data_mask  ),      

               .pe34__std__lane23_strm1_ready         ( pe34__std__lane23_strm1_ready      ),      
               .std__pe34__lane23_strm1_cntl          ( std__pe34__lane23_strm1_cntl       ),      
               .std__pe34__lane23_strm1_data          ( std__pe34__lane23_strm1_data       ),      
               .std__pe34__lane23_strm1_data_valid    ( std__pe34__lane23_strm1_data_valid ),      
               .std__pe34__lane23_strm1_data_mask     ( std__pe34__lane23_strm1_data_mask  ),      

               // PE 34, Lane 24                 
               .pe34__std__lane24_strm0_ready         ( pe34__std__lane24_strm0_ready      ),      
               .std__pe34__lane24_strm0_cntl          ( std__pe34__lane24_strm0_cntl       ),      
               .std__pe34__lane24_strm0_data          ( std__pe34__lane24_strm0_data       ),      
               .std__pe34__lane24_strm0_data_valid    ( std__pe34__lane24_strm0_data_valid ),      
               .std__pe34__lane24_strm0_data_mask     ( std__pe34__lane24_strm0_data_mask  ),      

               .pe34__std__lane24_strm1_ready         ( pe34__std__lane24_strm1_ready      ),      
               .std__pe34__lane24_strm1_cntl          ( std__pe34__lane24_strm1_cntl       ),      
               .std__pe34__lane24_strm1_data          ( std__pe34__lane24_strm1_data       ),      
               .std__pe34__lane24_strm1_data_valid    ( std__pe34__lane24_strm1_data_valid ),      
               .std__pe34__lane24_strm1_data_mask     ( std__pe34__lane24_strm1_data_mask  ),      

               // PE 34, Lane 25                 
               .pe34__std__lane25_strm0_ready         ( pe34__std__lane25_strm0_ready      ),      
               .std__pe34__lane25_strm0_cntl          ( std__pe34__lane25_strm0_cntl       ),      
               .std__pe34__lane25_strm0_data          ( std__pe34__lane25_strm0_data       ),      
               .std__pe34__lane25_strm0_data_valid    ( std__pe34__lane25_strm0_data_valid ),      
               .std__pe34__lane25_strm0_data_mask     ( std__pe34__lane25_strm0_data_mask  ),      

               .pe34__std__lane25_strm1_ready         ( pe34__std__lane25_strm1_ready      ),      
               .std__pe34__lane25_strm1_cntl          ( std__pe34__lane25_strm1_cntl       ),      
               .std__pe34__lane25_strm1_data          ( std__pe34__lane25_strm1_data       ),      
               .std__pe34__lane25_strm1_data_valid    ( std__pe34__lane25_strm1_data_valid ),      
               .std__pe34__lane25_strm1_data_mask     ( std__pe34__lane25_strm1_data_mask  ),      

               // PE 34, Lane 26                 
               .pe34__std__lane26_strm0_ready         ( pe34__std__lane26_strm0_ready      ),      
               .std__pe34__lane26_strm0_cntl          ( std__pe34__lane26_strm0_cntl       ),      
               .std__pe34__lane26_strm0_data          ( std__pe34__lane26_strm0_data       ),      
               .std__pe34__lane26_strm0_data_valid    ( std__pe34__lane26_strm0_data_valid ),      
               .std__pe34__lane26_strm0_data_mask     ( std__pe34__lane26_strm0_data_mask  ),      

               .pe34__std__lane26_strm1_ready         ( pe34__std__lane26_strm1_ready      ),      
               .std__pe34__lane26_strm1_cntl          ( std__pe34__lane26_strm1_cntl       ),      
               .std__pe34__lane26_strm1_data          ( std__pe34__lane26_strm1_data       ),      
               .std__pe34__lane26_strm1_data_valid    ( std__pe34__lane26_strm1_data_valid ),      
               .std__pe34__lane26_strm1_data_mask     ( std__pe34__lane26_strm1_data_mask  ),      

               // PE 34, Lane 27                 
               .pe34__std__lane27_strm0_ready         ( pe34__std__lane27_strm0_ready      ),      
               .std__pe34__lane27_strm0_cntl          ( std__pe34__lane27_strm0_cntl       ),      
               .std__pe34__lane27_strm0_data          ( std__pe34__lane27_strm0_data       ),      
               .std__pe34__lane27_strm0_data_valid    ( std__pe34__lane27_strm0_data_valid ),      
               .std__pe34__lane27_strm0_data_mask     ( std__pe34__lane27_strm0_data_mask  ),      

               .pe34__std__lane27_strm1_ready         ( pe34__std__lane27_strm1_ready      ),      
               .std__pe34__lane27_strm1_cntl          ( std__pe34__lane27_strm1_cntl       ),      
               .std__pe34__lane27_strm1_data          ( std__pe34__lane27_strm1_data       ),      
               .std__pe34__lane27_strm1_data_valid    ( std__pe34__lane27_strm1_data_valid ),      
               .std__pe34__lane27_strm1_data_mask     ( std__pe34__lane27_strm1_data_mask  ),      

               // PE 34, Lane 28                 
               .pe34__std__lane28_strm0_ready         ( pe34__std__lane28_strm0_ready      ),      
               .std__pe34__lane28_strm0_cntl          ( std__pe34__lane28_strm0_cntl       ),      
               .std__pe34__lane28_strm0_data          ( std__pe34__lane28_strm0_data       ),      
               .std__pe34__lane28_strm0_data_valid    ( std__pe34__lane28_strm0_data_valid ),      
               .std__pe34__lane28_strm0_data_mask     ( std__pe34__lane28_strm0_data_mask  ),      

               .pe34__std__lane28_strm1_ready         ( pe34__std__lane28_strm1_ready      ),      
               .std__pe34__lane28_strm1_cntl          ( std__pe34__lane28_strm1_cntl       ),      
               .std__pe34__lane28_strm1_data          ( std__pe34__lane28_strm1_data       ),      
               .std__pe34__lane28_strm1_data_valid    ( std__pe34__lane28_strm1_data_valid ),      
               .std__pe34__lane28_strm1_data_mask     ( std__pe34__lane28_strm1_data_mask  ),      

               // PE 34, Lane 29                 
               .pe34__std__lane29_strm0_ready         ( pe34__std__lane29_strm0_ready      ),      
               .std__pe34__lane29_strm0_cntl          ( std__pe34__lane29_strm0_cntl       ),      
               .std__pe34__lane29_strm0_data          ( std__pe34__lane29_strm0_data       ),      
               .std__pe34__lane29_strm0_data_valid    ( std__pe34__lane29_strm0_data_valid ),      
               .std__pe34__lane29_strm0_data_mask     ( std__pe34__lane29_strm0_data_mask  ),      

               .pe34__std__lane29_strm1_ready         ( pe34__std__lane29_strm1_ready      ),      
               .std__pe34__lane29_strm1_cntl          ( std__pe34__lane29_strm1_cntl       ),      
               .std__pe34__lane29_strm1_data          ( std__pe34__lane29_strm1_data       ),      
               .std__pe34__lane29_strm1_data_valid    ( std__pe34__lane29_strm1_data_valid ),      
               .std__pe34__lane29_strm1_data_mask     ( std__pe34__lane29_strm1_data_mask  ),      

               // PE 34, Lane 30                 
               .pe34__std__lane30_strm0_ready         ( pe34__std__lane30_strm0_ready      ),      
               .std__pe34__lane30_strm0_cntl          ( std__pe34__lane30_strm0_cntl       ),      
               .std__pe34__lane30_strm0_data          ( std__pe34__lane30_strm0_data       ),      
               .std__pe34__lane30_strm0_data_valid    ( std__pe34__lane30_strm0_data_valid ),      
               .std__pe34__lane30_strm0_data_mask     ( std__pe34__lane30_strm0_data_mask  ),      

               .pe34__std__lane30_strm1_ready         ( pe34__std__lane30_strm1_ready      ),      
               .std__pe34__lane30_strm1_cntl          ( std__pe34__lane30_strm1_cntl       ),      
               .std__pe34__lane30_strm1_data          ( std__pe34__lane30_strm1_data       ),      
               .std__pe34__lane30_strm1_data_valid    ( std__pe34__lane30_strm1_data_valid ),      
               .std__pe34__lane30_strm1_data_mask     ( std__pe34__lane30_strm1_data_mask  ),      

               // PE 34, Lane 31                 
               .pe34__std__lane31_strm0_ready         ( pe34__std__lane31_strm0_ready      ),      
               .std__pe34__lane31_strm0_cntl          ( std__pe34__lane31_strm0_cntl       ),      
               .std__pe34__lane31_strm0_data          ( std__pe34__lane31_strm0_data       ),      
               .std__pe34__lane31_strm0_data_valid    ( std__pe34__lane31_strm0_data_valid ),      
               .std__pe34__lane31_strm0_data_mask     ( std__pe34__lane31_strm0_data_mask  ),      

               .pe34__std__lane31_strm1_ready         ( pe34__std__lane31_strm1_ready      ),      
               .std__pe34__lane31_strm1_cntl          ( std__pe34__lane31_strm1_cntl       ),      
               .std__pe34__lane31_strm1_data          ( std__pe34__lane31_strm1_data       ),      
               .std__pe34__lane31_strm1_data_valid    ( std__pe34__lane31_strm1_data_valid ),      
               .std__pe34__lane31_strm1_data_mask     ( std__pe34__lane31_strm1_data_mask  ),      

               // PE 35, Lane 0                 
               .pe35__std__lane0_strm0_ready         ( pe35__std__lane0_strm0_ready      ),      
               .std__pe35__lane0_strm0_cntl          ( std__pe35__lane0_strm0_cntl       ),      
               .std__pe35__lane0_strm0_data          ( std__pe35__lane0_strm0_data       ),      
               .std__pe35__lane0_strm0_data_valid    ( std__pe35__lane0_strm0_data_valid ),      
               .std__pe35__lane0_strm0_data_mask     ( std__pe35__lane0_strm0_data_mask  ),      

               .pe35__std__lane0_strm1_ready         ( pe35__std__lane0_strm1_ready      ),      
               .std__pe35__lane0_strm1_cntl          ( std__pe35__lane0_strm1_cntl       ),      
               .std__pe35__lane0_strm1_data          ( std__pe35__lane0_strm1_data       ),      
               .std__pe35__lane0_strm1_data_valid    ( std__pe35__lane0_strm1_data_valid ),      
               .std__pe35__lane0_strm1_data_mask     ( std__pe35__lane0_strm1_data_mask  ),      

               // PE 35, Lane 1                 
               .pe35__std__lane1_strm0_ready         ( pe35__std__lane1_strm0_ready      ),      
               .std__pe35__lane1_strm0_cntl          ( std__pe35__lane1_strm0_cntl       ),      
               .std__pe35__lane1_strm0_data          ( std__pe35__lane1_strm0_data       ),      
               .std__pe35__lane1_strm0_data_valid    ( std__pe35__lane1_strm0_data_valid ),      
               .std__pe35__lane1_strm0_data_mask     ( std__pe35__lane1_strm0_data_mask  ),      

               .pe35__std__lane1_strm1_ready         ( pe35__std__lane1_strm1_ready      ),      
               .std__pe35__lane1_strm1_cntl          ( std__pe35__lane1_strm1_cntl       ),      
               .std__pe35__lane1_strm1_data          ( std__pe35__lane1_strm1_data       ),      
               .std__pe35__lane1_strm1_data_valid    ( std__pe35__lane1_strm1_data_valid ),      
               .std__pe35__lane1_strm1_data_mask     ( std__pe35__lane1_strm1_data_mask  ),      

               // PE 35, Lane 2                 
               .pe35__std__lane2_strm0_ready         ( pe35__std__lane2_strm0_ready      ),      
               .std__pe35__lane2_strm0_cntl          ( std__pe35__lane2_strm0_cntl       ),      
               .std__pe35__lane2_strm0_data          ( std__pe35__lane2_strm0_data       ),      
               .std__pe35__lane2_strm0_data_valid    ( std__pe35__lane2_strm0_data_valid ),      
               .std__pe35__lane2_strm0_data_mask     ( std__pe35__lane2_strm0_data_mask  ),      

               .pe35__std__lane2_strm1_ready         ( pe35__std__lane2_strm1_ready      ),      
               .std__pe35__lane2_strm1_cntl          ( std__pe35__lane2_strm1_cntl       ),      
               .std__pe35__lane2_strm1_data          ( std__pe35__lane2_strm1_data       ),      
               .std__pe35__lane2_strm1_data_valid    ( std__pe35__lane2_strm1_data_valid ),      
               .std__pe35__lane2_strm1_data_mask     ( std__pe35__lane2_strm1_data_mask  ),      

               // PE 35, Lane 3                 
               .pe35__std__lane3_strm0_ready         ( pe35__std__lane3_strm0_ready      ),      
               .std__pe35__lane3_strm0_cntl          ( std__pe35__lane3_strm0_cntl       ),      
               .std__pe35__lane3_strm0_data          ( std__pe35__lane3_strm0_data       ),      
               .std__pe35__lane3_strm0_data_valid    ( std__pe35__lane3_strm0_data_valid ),      
               .std__pe35__lane3_strm0_data_mask     ( std__pe35__lane3_strm0_data_mask  ),      

               .pe35__std__lane3_strm1_ready         ( pe35__std__lane3_strm1_ready      ),      
               .std__pe35__lane3_strm1_cntl          ( std__pe35__lane3_strm1_cntl       ),      
               .std__pe35__lane3_strm1_data          ( std__pe35__lane3_strm1_data       ),      
               .std__pe35__lane3_strm1_data_valid    ( std__pe35__lane3_strm1_data_valid ),      
               .std__pe35__lane3_strm1_data_mask     ( std__pe35__lane3_strm1_data_mask  ),      

               // PE 35, Lane 4                 
               .pe35__std__lane4_strm0_ready         ( pe35__std__lane4_strm0_ready      ),      
               .std__pe35__lane4_strm0_cntl          ( std__pe35__lane4_strm0_cntl       ),      
               .std__pe35__lane4_strm0_data          ( std__pe35__lane4_strm0_data       ),      
               .std__pe35__lane4_strm0_data_valid    ( std__pe35__lane4_strm0_data_valid ),      
               .std__pe35__lane4_strm0_data_mask     ( std__pe35__lane4_strm0_data_mask  ),      

               .pe35__std__lane4_strm1_ready         ( pe35__std__lane4_strm1_ready      ),      
               .std__pe35__lane4_strm1_cntl          ( std__pe35__lane4_strm1_cntl       ),      
               .std__pe35__lane4_strm1_data          ( std__pe35__lane4_strm1_data       ),      
               .std__pe35__lane4_strm1_data_valid    ( std__pe35__lane4_strm1_data_valid ),      
               .std__pe35__lane4_strm1_data_mask     ( std__pe35__lane4_strm1_data_mask  ),      

               // PE 35, Lane 5                 
               .pe35__std__lane5_strm0_ready         ( pe35__std__lane5_strm0_ready      ),      
               .std__pe35__lane5_strm0_cntl          ( std__pe35__lane5_strm0_cntl       ),      
               .std__pe35__lane5_strm0_data          ( std__pe35__lane5_strm0_data       ),      
               .std__pe35__lane5_strm0_data_valid    ( std__pe35__lane5_strm0_data_valid ),      
               .std__pe35__lane5_strm0_data_mask     ( std__pe35__lane5_strm0_data_mask  ),      

               .pe35__std__lane5_strm1_ready         ( pe35__std__lane5_strm1_ready      ),      
               .std__pe35__lane5_strm1_cntl          ( std__pe35__lane5_strm1_cntl       ),      
               .std__pe35__lane5_strm1_data          ( std__pe35__lane5_strm1_data       ),      
               .std__pe35__lane5_strm1_data_valid    ( std__pe35__lane5_strm1_data_valid ),      
               .std__pe35__lane5_strm1_data_mask     ( std__pe35__lane5_strm1_data_mask  ),      

               // PE 35, Lane 6                 
               .pe35__std__lane6_strm0_ready         ( pe35__std__lane6_strm0_ready      ),      
               .std__pe35__lane6_strm0_cntl          ( std__pe35__lane6_strm0_cntl       ),      
               .std__pe35__lane6_strm0_data          ( std__pe35__lane6_strm0_data       ),      
               .std__pe35__lane6_strm0_data_valid    ( std__pe35__lane6_strm0_data_valid ),      
               .std__pe35__lane6_strm0_data_mask     ( std__pe35__lane6_strm0_data_mask  ),      

               .pe35__std__lane6_strm1_ready         ( pe35__std__lane6_strm1_ready      ),      
               .std__pe35__lane6_strm1_cntl          ( std__pe35__lane6_strm1_cntl       ),      
               .std__pe35__lane6_strm1_data          ( std__pe35__lane6_strm1_data       ),      
               .std__pe35__lane6_strm1_data_valid    ( std__pe35__lane6_strm1_data_valid ),      
               .std__pe35__lane6_strm1_data_mask     ( std__pe35__lane6_strm1_data_mask  ),      

               // PE 35, Lane 7                 
               .pe35__std__lane7_strm0_ready         ( pe35__std__lane7_strm0_ready      ),      
               .std__pe35__lane7_strm0_cntl          ( std__pe35__lane7_strm0_cntl       ),      
               .std__pe35__lane7_strm0_data          ( std__pe35__lane7_strm0_data       ),      
               .std__pe35__lane7_strm0_data_valid    ( std__pe35__lane7_strm0_data_valid ),      
               .std__pe35__lane7_strm0_data_mask     ( std__pe35__lane7_strm0_data_mask  ),      

               .pe35__std__lane7_strm1_ready         ( pe35__std__lane7_strm1_ready      ),      
               .std__pe35__lane7_strm1_cntl          ( std__pe35__lane7_strm1_cntl       ),      
               .std__pe35__lane7_strm1_data          ( std__pe35__lane7_strm1_data       ),      
               .std__pe35__lane7_strm1_data_valid    ( std__pe35__lane7_strm1_data_valid ),      
               .std__pe35__lane7_strm1_data_mask     ( std__pe35__lane7_strm1_data_mask  ),      

               // PE 35, Lane 8                 
               .pe35__std__lane8_strm0_ready         ( pe35__std__lane8_strm0_ready      ),      
               .std__pe35__lane8_strm0_cntl          ( std__pe35__lane8_strm0_cntl       ),      
               .std__pe35__lane8_strm0_data          ( std__pe35__lane8_strm0_data       ),      
               .std__pe35__lane8_strm0_data_valid    ( std__pe35__lane8_strm0_data_valid ),      
               .std__pe35__lane8_strm0_data_mask     ( std__pe35__lane8_strm0_data_mask  ),      

               .pe35__std__lane8_strm1_ready         ( pe35__std__lane8_strm1_ready      ),      
               .std__pe35__lane8_strm1_cntl          ( std__pe35__lane8_strm1_cntl       ),      
               .std__pe35__lane8_strm1_data          ( std__pe35__lane8_strm1_data       ),      
               .std__pe35__lane8_strm1_data_valid    ( std__pe35__lane8_strm1_data_valid ),      
               .std__pe35__lane8_strm1_data_mask     ( std__pe35__lane8_strm1_data_mask  ),      

               // PE 35, Lane 9                 
               .pe35__std__lane9_strm0_ready         ( pe35__std__lane9_strm0_ready      ),      
               .std__pe35__lane9_strm0_cntl          ( std__pe35__lane9_strm0_cntl       ),      
               .std__pe35__lane9_strm0_data          ( std__pe35__lane9_strm0_data       ),      
               .std__pe35__lane9_strm0_data_valid    ( std__pe35__lane9_strm0_data_valid ),      
               .std__pe35__lane9_strm0_data_mask     ( std__pe35__lane9_strm0_data_mask  ),      

               .pe35__std__lane9_strm1_ready         ( pe35__std__lane9_strm1_ready      ),      
               .std__pe35__lane9_strm1_cntl          ( std__pe35__lane9_strm1_cntl       ),      
               .std__pe35__lane9_strm1_data          ( std__pe35__lane9_strm1_data       ),      
               .std__pe35__lane9_strm1_data_valid    ( std__pe35__lane9_strm1_data_valid ),      
               .std__pe35__lane9_strm1_data_mask     ( std__pe35__lane9_strm1_data_mask  ),      

               // PE 35, Lane 10                 
               .pe35__std__lane10_strm0_ready         ( pe35__std__lane10_strm0_ready      ),      
               .std__pe35__lane10_strm0_cntl          ( std__pe35__lane10_strm0_cntl       ),      
               .std__pe35__lane10_strm0_data          ( std__pe35__lane10_strm0_data       ),      
               .std__pe35__lane10_strm0_data_valid    ( std__pe35__lane10_strm0_data_valid ),      
               .std__pe35__lane10_strm0_data_mask     ( std__pe35__lane10_strm0_data_mask  ),      

               .pe35__std__lane10_strm1_ready         ( pe35__std__lane10_strm1_ready      ),      
               .std__pe35__lane10_strm1_cntl          ( std__pe35__lane10_strm1_cntl       ),      
               .std__pe35__lane10_strm1_data          ( std__pe35__lane10_strm1_data       ),      
               .std__pe35__lane10_strm1_data_valid    ( std__pe35__lane10_strm1_data_valid ),      
               .std__pe35__lane10_strm1_data_mask     ( std__pe35__lane10_strm1_data_mask  ),      

               // PE 35, Lane 11                 
               .pe35__std__lane11_strm0_ready         ( pe35__std__lane11_strm0_ready      ),      
               .std__pe35__lane11_strm0_cntl          ( std__pe35__lane11_strm0_cntl       ),      
               .std__pe35__lane11_strm0_data          ( std__pe35__lane11_strm0_data       ),      
               .std__pe35__lane11_strm0_data_valid    ( std__pe35__lane11_strm0_data_valid ),      
               .std__pe35__lane11_strm0_data_mask     ( std__pe35__lane11_strm0_data_mask  ),      

               .pe35__std__lane11_strm1_ready         ( pe35__std__lane11_strm1_ready      ),      
               .std__pe35__lane11_strm1_cntl          ( std__pe35__lane11_strm1_cntl       ),      
               .std__pe35__lane11_strm1_data          ( std__pe35__lane11_strm1_data       ),      
               .std__pe35__lane11_strm1_data_valid    ( std__pe35__lane11_strm1_data_valid ),      
               .std__pe35__lane11_strm1_data_mask     ( std__pe35__lane11_strm1_data_mask  ),      

               // PE 35, Lane 12                 
               .pe35__std__lane12_strm0_ready         ( pe35__std__lane12_strm0_ready      ),      
               .std__pe35__lane12_strm0_cntl          ( std__pe35__lane12_strm0_cntl       ),      
               .std__pe35__lane12_strm0_data          ( std__pe35__lane12_strm0_data       ),      
               .std__pe35__lane12_strm0_data_valid    ( std__pe35__lane12_strm0_data_valid ),      
               .std__pe35__lane12_strm0_data_mask     ( std__pe35__lane12_strm0_data_mask  ),      

               .pe35__std__lane12_strm1_ready         ( pe35__std__lane12_strm1_ready      ),      
               .std__pe35__lane12_strm1_cntl          ( std__pe35__lane12_strm1_cntl       ),      
               .std__pe35__lane12_strm1_data          ( std__pe35__lane12_strm1_data       ),      
               .std__pe35__lane12_strm1_data_valid    ( std__pe35__lane12_strm1_data_valid ),      
               .std__pe35__lane12_strm1_data_mask     ( std__pe35__lane12_strm1_data_mask  ),      

               // PE 35, Lane 13                 
               .pe35__std__lane13_strm0_ready         ( pe35__std__lane13_strm0_ready      ),      
               .std__pe35__lane13_strm0_cntl          ( std__pe35__lane13_strm0_cntl       ),      
               .std__pe35__lane13_strm0_data          ( std__pe35__lane13_strm0_data       ),      
               .std__pe35__lane13_strm0_data_valid    ( std__pe35__lane13_strm0_data_valid ),      
               .std__pe35__lane13_strm0_data_mask     ( std__pe35__lane13_strm0_data_mask  ),      

               .pe35__std__lane13_strm1_ready         ( pe35__std__lane13_strm1_ready      ),      
               .std__pe35__lane13_strm1_cntl          ( std__pe35__lane13_strm1_cntl       ),      
               .std__pe35__lane13_strm1_data          ( std__pe35__lane13_strm1_data       ),      
               .std__pe35__lane13_strm1_data_valid    ( std__pe35__lane13_strm1_data_valid ),      
               .std__pe35__lane13_strm1_data_mask     ( std__pe35__lane13_strm1_data_mask  ),      

               // PE 35, Lane 14                 
               .pe35__std__lane14_strm0_ready         ( pe35__std__lane14_strm0_ready      ),      
               .std__pe35__lane14_strm0_cntl          ( std__pe35__lane14_strm0_cntl       ),      
               .std__pe35__lane14_strm0_data          ( std__pe35__lane14_strm0_data       ),      
               .std__pe35__lane14_strm0_data_valid    ( std__pe35__lane14_strm0_data_valid ),      
               .std__pe35__lane14_strm0_data_mask     ( std__pe35__lane14_strm0_data_mask  ),      

               .pe35__std__lane14_strm1_ready         ( pe35__std__lane14_strm1_ready      ),      
               .std__pe35__lane14_strm1_cntl          ( std__pe35__lane14_strm1_cntl       ),      
               .std__pe35__lane14_strm1_data          ( std__pe35__lane14_strm1_data       ),      
               .std__pe35__lane14_strm1_data_valid    ( std__pe35__lane14_strm1_data_valid ),      
               .std__pe35__lane14_strm1_data_mask     ( std__pe35__lane14_strm1_data_mask  ),      

               // PE 35, Lane 15                 
               .pe35__std__lane15_strm0_ready         ( pe35__std__lane15_strm0_ready      ),      
               .std__pe35__lane15_strm0_cntl          ( std__pe35__lane15_strm0_cntl       ),      
               .std__pe35__lane15_strm0_data          ( std__pe35__lane15_strm0_data       ),      
               .std__pe35__lane15_strm0_data_valid    ( std__pe35__lane15_strm0_data_valid ),      
               .std__pe35__lane15_strm0_data_mask     ( std__pe35__lane15_strm0_data_mask  ),      

               .pe35__std__lane15_strm1_ready         ( pe35__std__lane15_strm1_ready      ),      
               .std__pe35__lane15_strm1_cntl          ( std__pe35__lane15_strm1_cntl       ),      
               .std__pe35__lane15_strm1_data          ( std__pe35__lane15_strm1_data       ),      
               .std__pe35__lane15_strm1_data_valid    ( std__pe35__lane15_strm1_data_valid ),      
               .std__pe35__lane15_strm1_data_mask     ( std__pe35__lane15_strm1_data_mask  ),      

               // PE 35, Lane 16                 
               .pe35__std__lane16_strm0_ready         ( pe35__std__lane16_strm0_ready      ),      
               .std__pe35__lane16_strm0_cntl          ( std__pe35__lane16_strm0_cntl       ),      
               .std__pe35__lane16_strm0_data          ( std__pe35__lane16_strm0_data       ),      
               .std__pe35__lane16_strm0_data_valid    ( std__pe35__lane16_strm0_data_valid ),      
               .std__pe35__lane16_strm0_data_mask     ( std__pe35__lane16_strm0_data_mask  ),      

               .pe35__std__lane16_strm1_ready         ( pe35__std__lane16_strm1_ready      ),      
               .std__pe35__lane16_strm1_cntl          ( std__pe35__lane16_strm1_cntl       ),      
               .std__pe35__lane16_strm1_data          ( std__pe35__lane16_strm1_data       ),      
               .std__pe35__lane16_strm1_data_valid    ( std__pe35__lane16_strm1_data_valid ),      
               .std__pe35__lane16_strm1_data_mask     ( std__pe35__lane16_strm1_data_mask  ),      

               // PE 35, Lane 17                 
               .pe35__std__lane17_strm0_ready         ( pe35__std__lane17_strm0_ready      ),      
               .std__pe35__lane17_strm0_cntl          ( std__pe35__lane17_strm0_cntl       ),      
               .std__pe35__lane17_strm0_data          ( std__pe35__lane17_strm0_data       ),      
               .std__pe35__lane17_strm0_data_valid    ( std__pe35__lane17_strm0_data_valid ),      
               .std__pe35__lane17_strm0_data_mask     ( std__pe35__lane17_strm0_data_mask  ),      

               .pe35__std__lane17_strm1_ready         ( pe35__std__lane17_strm1_ready      ),      
               .std__pe35__lane17_strm1_cntl          ( std__pe35__lane17_strm1_cntl       ),      
               .std__pe35__lane17_strm1_data          ( std__pe35__lane17_strm1_data       ),      
               .std__pe35__lane17_strm1_data_valid    ( std__pe35__lane17_strm1_data_valid ),      
               .std__pe35__lane17_strm1_data_mask     ( std__pe35__lane17_strm1_data_mask  ),      

               // PE 35, Lane 18                 
               .pe35__std__lane18_strm0_ready         ( pe35__std__lane18_strm0_ready      ),      
               .std__pe35__lane18_strm0_cntl          ( std__pe35__lane18_strm0_cntl       ),      
               .std__pe35__lane18_strm0_data          ( std__pe35__lane18_strm0_data       ),      
               .std__pe35__lane18_strm0_data_valid    ( std__pe35__lane18_strm0_data_valid ),      
               .std__pe35__lane18_strm0_data_mask     ( std__pe35__lane18_strm0_data_mask  ),      

               .pe35__std__lane18_strm1_ready         ( pe35__std__lane18_strm1_ready      ),      
               .std__pe35__lane18_strm1_cntl          ( std__pe35__lane18_strm1_cntl       ),      
               .std__pe35__lane18_strm1_data          ( std__pe35__lane18_strm1_data       ),      
               .std__pe35__lane18_strm1_data_valid    ( std__pe35__lane18_strm1_data_valid ),      
               .std__pe35__lane18_strm1_data_mask     ( std__pe35__lane18_strm1_data_mask  ),      

               // PE 35, Lane 19                 
               .pe35__std__lane19_strm0_ready         ( pe35__std__lane19_strm0_ready      ),      
               .std__pe35__lane19_strm0_cntl          ( std__pe35__lane19_strm0_cntl       ),      
               .std__pe35__lane19_strm0_data          ( std__pe35__lane19_strm0_data       ),      
               .std__pe35__lane19_strm0_data_valid    ( std__pe35__lane19_strm0_data_valid ),      
               .std__pe35__lane19_strm0_data_mask     ( std__pe35__lane19_strm0_data_mask  ),      

               .pe35__std__lane19_strm1_ready         ( pe35__std__lane19_strm1_ready      ),      
               .std__pe35__lane19_strm1_cntl          ( std__pe35__lane19_strm1_cntl       ),      
               .std__pe35__lane19_strm1_data          ( std__pe35__lane19_strm1_data       ),      
               .std__pe35__lane19_strm1_data_valid    ( std__pe35__lane19_strm1_data_valid ),      
               .std__pe35__lane19_strm1_data_mask     ( std__pe35__lane19_strm1_data_mask  ),      

               // PE 35, Lane 20                 
               .pe35__std__lane20_strm0_ready         ( pe35__std__lane20_strm0_ready      ),      
               .std__pe35__lane20_strm0_cntl          ( std__pe35__lane20_strm0_cntl       ),      
               .std__pe35__lane20_strm0_data          ( std__pe35__lane20_strm0_data       ),      
               .std__pe35__lane20_strm0_data_valid    ( std__pe35__lane20_strm0_data_valid ),      
               .std__pe35__lane20_strm0_data_mask     ( std__pe35__lane20_strm0_data_mask  ),      

               .pe35__std__lane20_strm1_ready         ( pe35__std__lane20_strm1_ready      ),      
               .std__pe35__lane20_strm1_cntl          ( std__pe35__lane20_strm1_cntl       ),      
               .std__pe35__lane20_strm1_data          ( std__pe35__lane20_strm1_data       ),      
               .std__pe35__lane20_strm1_data_valid    ( std__pe35__lane20_strm1_data_valid ),      
               .std__pe35__lane20_strm1_data_mask     ( std__pe35__lane20_strm1_data_mask  ),      

               // PE 35, Lane 21                 
               .pe35__std__lane21_strm0_ready         ( pe35__std__lane21_strm0_ready      ),      
               .std__pe35__lane21_strm0_cntl          ( std__pe35__lane21_strm0_cntl       ),      
               .std__pe35__lane21_strm0_data          ( std__pe35__lane21_strm0_data       ),      
               .std__pe35__lane21_strm0_data_valid    ( std__pe35__lane21_strm0_data_valid ),      
               .std__pe35__lane21_strm0_data_mask     ( std__pe35__lane21_strm0_data_mask  ),      

               .pe35__std__lane21_strm1_ready         ( pe35__std__lane21_strm1_ready      ),      
               .std__pe35__lane21_strm1_cntl          ( std__pe35__lane21_strm1_cntl       ),      
               .std__pe35__lane21_strm1_data          ( std__pe35__lane21_strm1_data       ),      
               .std__pe35__lane21_strm1_data_valid    ( std__pe35__lane21_strm1_data_valid ),      
               .std__pe35__lane21_strm1_data_mask     ( std__pe35__lane21_strm1_data_mask  ),      

               // PE 35, Lane 22                 
               .pe35__std__lane22_strm0_ready         ( pe35__std__lane22_strm0_ready      ),      
               .std__pe35__lane22_strm0_cntl          ( std__pe35__lane22_strm0_cntl       ),      
               .std__pe35__lane22_strm0_data          ( std__pe35__lane22_strm0_data       ),      
               .std__pe35__lane22_strm0_data_valid    ( std__pe35__lane22_strm0_data_valid ),      
               .std__pe35__lane22_strm0_data_mask     ( std__pe35__lane22_strm0_data_mask  ),      

               .pe35__std__lane22_strm1_ready         ( pe35__std__lane22_strm1_ready      ),      
               .std__pe35__lane22_strm1_cntl          ( std__pe35__lane22_strm1_cntl       ),      
               .std__pe35__lane22_strm1_data          ( std__pe35__lane22_strm1_data       ),      
               .std__pe35__lane22_strm1_data_valid    ( std__pe35__lane22_strm1_data_valid ),      
               .std__pe35__lane22_strm1_data_mask     ( std__pe35__lane22_strm1_data_mask  ),      

               // PE 35, Lane 23                 
               .pe35__std__lane23_strm0_ready         ( pe35__std__lane23_strm0_ready      ),      
               .std__pe35__lane23_strm0_cntl          ( std__pe35__lane23_strm0_cntl       ),      
               .std__pe35__lane23_strm0_data          ( std__pe35__lane23_strm0_data       ),      
               .std__pe35__lane23_strm0_data_valid    ( std__pe35__lane23_strm0_data_valid ),      
               .std__pe35__lane23_strm0_data_mask     ( std__pe35__lane23_strm0_data_mask  ),      

               .pe35__std__lane23_strm1_ready         ( pe35__std__lane23_strm1_ready      ),      
               .std__pe35__lane23_strm1_cntl          ( std__pe35__lane23_strm1_cntl       ),      
               .std__pe35__lane23_strm1_data          ( std__pe35__lane23_strm1_data       ),      
               .std__pe35__lane23_strm1_data_valid    ( std__pe35__lane23_strm1_data_valid ),      
               .std__pe35__lane23_strm1_data_mask     ( std__pe35__lane23_strm1_data_mask  ),      

               // PE 35, Lane 24                 
               .pe35__std__lane24_strm0_ready         ( pe35__std__lane24_strm0_ready      ),      
               .std__pe35__lane24_strm0_cntl          ( std__pe35__lane24_strm0_cntl       ),      
               .std__pe35__lane24_strm0_data          ( std__pe35__lane24_strm0_data       ),      
               .std__pe35__lane24_strm0_data_valid    ( std__pe35__lane24_strm0_data_valid ),      
               .std__pe35__lane24_strm0_data_mask     ( std__pe35__lane24_strm0_data_mask  ),      

               .pe35__std__lane24_strm1_ready         ( pe35__std__lane24_strm1_ready      ),      
               .std__pe35__lane24_strm1_cntl          ( std__pe35__lane24_strm1_cntl       ),      
               .std__pe35__lane24_strm1_data          ( std__pe35__lane24_strm1_data       ),      
               .std__pe35__lane24_strm1_data_valid    ( std__pe35__lane24_strm1_data_valid ),      
               .std__pe35__lane24_strm1_data_mask     ( std__pe35__lane24_strm1_data_mask  ),      

               // PE 35, Lane 25                 
               .pe35__std__lane25_strm0_ready         ( pe35__std__lane25_strm0_ready      ),      
               .std__pe35__lane25_strm0_cntl          ( std__pe35__lane25_strm0_cntl       ),      
               .std__pe35__lane25_strm0_data          ( std__pe35__lane25_strm0_data       ),      
               .std__pe35__lane25_strm0_data_valid    ( std__pe35__lane25_strm0_data_valid ),      
               .std__pe35__lane25_strm0_data_mask     ( std__pe35__lane25_strm0_data_mask  ),      

               .pe35__std__lane25_strm1_ready         ( pe35__std__lane25_strm1_ready      ),      
               .std__pe35__lane25_strm1_cntl          ( std__pe35__lane25_strm1_cntl       ),      
               .std__pe35__lane25_strm1_data          ( std__pe35__lane25_strm1_data       ),      
               .std__pe35__lane25_strm1_data_valid    ( std__pe35__lane25_strm1_data_valid ),      
               .std__pe35__lane25_strm1_data_mask     ( std__pe35__lane25_strm1_data_mask  ),      

               // PE 35, Lane 26                 
               .pe35__std__lane26_strm0_ready         ( pe35__std__lane26_strm0_ready      ),      
               .std__pe35__lane26_strm0_cntl          ( std__pe35__lane26_strm0_cntl       ),      
               .std__pe35__lane26_strm0_data          ( std__pe35__lane26_strm0_data       ),      
               .std__pe35__lane26_strm0_data_valid    ( std__pe35__lane26_strm0_data_valid ),      
               .std__pe35__lane26_strm0_data_mask     ( std__pe35__lane26_strm0_data_mask  ),      

               .pe35__std__lane26_strm1_ready         ( pe35__std__lane26_strm1_ready      ),      
               .std__pe35__lane26_strm1_cntl          ( std__pe35__lane26_strm1_cntl       ),      
               .std__pe35__lane26_strm1_data          ( std__pe35__lane26_strm1_data       ),      
               .std__pe35__lane26_strm1_data_valid    ( std__pe35__lane26_strm1_data_valid ),      
               .std__pe35__lane26_strm1_data_mask     ( std__pe35__lane26_strm1_data_mask  ),      

               // PE 35, Lane 27                 
               .pe35__std__lane27_strm0_ready         ( pe35__std__lane27_strm0_ready      ),      
               .std__pe35__lane27_strm0_cntl          ( std__pe35__lane27_strm0_cntl       ),      
               .std__pe35__lane27_strm0_data          ( std__pe35__lane27_strm0_data       ),      
               .std__pe35__lane27_strm0_data_valid    ( std__pe35__lane27_strm0_data_valid ),      
               .std__pe35__lane27_strm0_data_mask     ( std__pe35__lane27_strm0_data_mask  ),      

               .pe35__std__lane27_strm1_ready         ( pe35__std__lane27_strm1_ready      ),      
               .std__pe35__lane27_strm1_cntl          ( std__pe35__lane27_strm1_cntl       ),      
               .std__pe35__lane27_strm1_data          ( std__pe35__lane27_strm1_data       ),      
               .std__pe35__lane27_strm1_data_valid    ( std__pe35__lane27_strm1_data_valid ),      
               .std__pe35__lane27_strm1_data_mask     ( std__pe35__lane27_strm1_data_mask  ),      

               // PE 35, Lane 28                 
               .pe35__std__lane28_strm0_ready         ( pe35__std__lane28_strm0_ready      ),      
               .std__pe35__lane28_strm0_cntl          ( std__pe35__lane28_strm0_cntl       ),      
               .std__pe35__lane28_strm0_data          ( std__pe35__lane28_strm0_data       ),      
               .std__pe35__lane28_strm0_data_valid    ( std__pe35__lane28_strm0_data_valid ),      
               .std__pe35__lane28_strm0_data_mask     ( std__pe35__lane28_strm0_data_mask  ),      

               .pe35__std__lane28_strm1_ready         ( pe35__std__lane28_strm1_ready      ),      
               .std__pe35__lane28_strm1_cntl          ( std__pe35__lane28_strm1_cntl       ),      
               .std__pe35__lane28_strm1_data          ( std__pe35__lane28_strm1_data       ),      
               .std__pe35__lane28_strm1_data_valid    ( std__pe35__lane28_strm1_data_valid ),      
               .std__pe35__lane28_strm1_data_mask     ( std__pe35__lane28_strm1_data_mask  ),      

               // PE 35, Lane 29                 
               .pe35__std__lane29_strm0_ready         ( pe35__std__lane29_strm0_ready      ),      
               .std__pe35__lane29_strm0_cntl          ( std__pe35__lane29_strm0_cntl       ),      
               .std__pe35__lane29_strm0_data          ( std__pe35__lane29_strm0_data       ),      
               .std__pe35__lane29_strm0_data_valid    ( std__pe35__lane29_strm0_data_valid ),      
               .std__pe35__lane29_strm0_data_mask     ( std__pe35__lane29_strm0_data_mask  ),      

               .pe35__std__lane29_strm1_ready         ( pe35__std__lane29_strm1_ready      ),      
               .std__pe35__lane29_strm1_cntl          ( std__pe35__lane29_strm1_cntl       ),      
               .std__pe35__lane29_strm1_data          ( std__pe35__lane29_strm1_data       ),      
               .std__pe35__lane29_strm1_data_valid    ( std__pe35__lane29_strm1_data_valid ),      
               .std__pe35__lane29_strm1_data_mask     ( std__pe35__lane29_strm1_data_mask  ),      

               // PE 35, Lane 30                 
               .pe35__std__lane30_strm0_ready         ( pe35__std__lane30_strm0_ready      ),      
               .std__pe35__lane30_strm0_cntl          ( std__pe35__lane30_strm0_cntl       ),      
               .std__pe35__lane30_strm0_data          ( std__pe35__lane30_strm0_data       ),      
               .std__pe35__lane30_strm0_data_valid    ( std__pe35__lane30_strm0_data_valid ),      
               .std__pe35__lane30_strm0_data_mask     ( std__pe35__lane30_strm0_data_mask  ),      

               .pe35__std__lane30_strm1_ready         ( pe35__std__lane30_strm1_ready      ),      
               .std__pe35__lane30_strm1_cntl          ( std__pe35__lane30_strm1_cntl       ),      
               .std__pe35__lane30_strm1_data          ( std__pe35__lane30_strm1_data       ),      
               .std__pe35__lane30_strm1_data_valid    ( std__pe35__lane30_strm1_data_valid ),      
               .std__pe35__lane30_strm1_data_mask     ( std__pe35__lane30_strm1_data_mask  ),      

               // PE 35, Lane 31                 
               .pe35__std__lane31_strm0_ready         ( pe35__std__lane31_strm0_ready      ),      
               .std__pe35__lane31_strm0_cntl          ( std__pe35__lane31_strm0_cntl       ),      
               .std__pe35__lane31_strm0_data          ( std__pe35__lane31_strm0_data       ),      
               .std__pe35__lane31_strm0_data_valid    ( std__pe35__lane31_strm0_data_valid ),      
               .std__pe35__lane31_strm0_data_mask     ( std__pe35__lane31_strm0_data_mask  ),      

               .pe35__std__lane31_strm1_ready         ( pe35__std__lane31_strm1_ready      ),      
               .std__pe35__lane31_strm1_cntl          ( std__pe35__lane31_strm1_cntl       ),      
               .std__pe35__lane31_strm1_data          ( std__pe35__lane31_strm1_data       ),      
               .std__pe35__lane31_strm1_data_valid    ( std__pe35__lane31_strm1_data_valid ),      
               .std__pe35__lane31_strm1_data_mask     ( std__pe35__lane31_strm1_data_mask  ),      

               // PE 36, Lane 0                 
               .pe36__std__lane0_strm0_ready         ( pe36__std__lane0_strm0_ready      ),      
               .std__pe36__lane0_strm0_cntl          ( std__pe36__lane0_strm0_cntl       ),      
               .std__pe36__lane0_strm0_data          ( std__pe36__lane0_strm0_data       ),      
               .std__pe36__lane0_strm0_data_valid    ( std__pe36__lane0_strm0_data_valid ),      
               .std__pe36__lane0_strm0_data_mask     ( std__pe36__lane0_strm0_data_mask  ),      

               .pe36__std__lane0_strm1_ready         ( pe36__std__lane0_strm1_ready      ),      
               .std__pe36__lane0_strm1_cntl          ( std__pe36__lane0_strm1_cntl       ),      
               .std__pe36__lane0_strm1_data          ( std__pe36__lane0_strm1_data       ),      
               .std__pe36__lane0_strm1_data_valid    ( std__pe36__lane0_strm1_data_valid ),      
               .std__pe36__lane0_strm1_data_mask     ( std__pe36__lane0_strm1_data_mask  ),      

               // PE 36, Lane 1                 
               .pe36__std__lane1_strm0_ready         ( pe36__std__lane1_strm0_ready      ),      
               .std__pe36__lane1_strm0_cntl          ( std__pe36__lane1_strm0_cntl       ),      
               .std__pe36__lane1_strm0_data          ( std__pe36__lane1_strm0_data       ),      
               .std__pe36__lane1_strm0_data_valid    ( std__pe36__lane1_strm0_data_valid ),      
               .std__pe36__lane1_strm0_data_mask     ( std__pe36__lane1_strm0_data_mask  ),      

               .pe36__std__lane1_strm1_ready         ( pe36__std__lane1_strm1_ready      ),      
               .std__pe36__lane1_strm1_cntl          ( std__pe36__lane1_strm1_cntl       ),      
               .std__pe36__lane1_strm1_data          ( std__pe36__lane1_strm1_data       ),      
               .std__pe36__lane1_strm1_data_valid    ( std__pe36__lane1_strm1_data_valid ),      
               .std__pe36__lane1_strm1_data_mask     ( std__pe36__lane1_strm1_data_mask  ),      

               // PE 36, Lane 2                 
               .pe36__std__lane2_strm0_ready         ( pe36__std__lane2_strm0_ready      ),      
               .std__pe36__lane2_strm0_cntl          ( std__pe36__lane2_strm0_cntl       ),      
               .std__pe36__lane2_strm0_data          ( std__pe36__lane2_strm0_data       ),      
               .std__pe36__lane2_strm0_data_valid    ( std__pe36__lane2_strm0_data_valid ),      
               .std__pe36__lane2_strm0_data_mask     ( std__pe36__lane2_strm0_data_mask  ),      

               .pe36__std__lane2_strm1_ready         ( pe36__std__lane2_strm1_ready      ),      
               .std__pe36__lane2_strm1_cntl          ( std__pe36__lane2_strm1_cntl       ),      
               .std__pe36__lane2_strm1_data          ( std__pe36__lane2_strm1_data       ),      
               .std__pe36__lane2_strm1_data_valid    ( std__pe36__lane2_strm1_data_valid ),      
               .std__pe36__lane2_strm1_data_mask     ( std__pe36__lane2_strm1_data_mask  ),      

               // PE 36, Lane 3                 
               .pe36__std__lane3_strm0_ready         ( pe36__std__lane3_strm0_ready      ),      
               .std__pe36__lane3_strm0_cntl          ( std__pe36__lane3_strm0_cntl       ),      
               .std__pe36__lane3_strm0_data          ( std__pe36__lane3_strm0_data       ),      
               .std__pe36__lane3_strm0_data_valid    ( std__pe36__lane3_strm0_data_valid ),      
               .std__pe36__lane3_strm0_data_mask     ( std__pe36__lane3_strm0_data_mask  ),      

               .pe36__std__lane3_strm1_ready         ( pe36__std__lane3_strm1_ready      ),      
               .std__pe36__lane3_strm1_cntl          ( std__pe36__lane3_strm1_cntl       ),      
               .std__pe36__lane3_strm1_data          ( std__pe36__lane3_strm1_data       ),      
               .std__pe36__lane3_strm1_data_valid    ( std__pe36__lane3_strm1_data_valid ),      
               .std__pe36__lane3_strm1_data_mask     ( std__pe36__lane3_strm1_data_mask  ),      

               // PE 36, Lane 4                 
               .pe36__std__lane4_strm0_ready         ( pe36__std__lane4_strm0_ready      ),      
               .std__pe36__lane4_strm0_cntl          ( std__pe36__lane4_strm0_cntl       ),      
               .std__pe36__lane4_strm0_data          ( std__pe36__lane4_strm0_data       ),      
               .std__pe36__lane4_strm0_data_valid    ( std__pe36__lane4_strm0_data_valid ),      
               .std__pe36__lane4_strm0_data_mask     ( std__pe36__lane4_strm0_data_mask  ),      

               .pe36__std__lane4_strm1_ready         ( pe36__std__lane4_strm1_ready      ),      
               .std__pe36__lane4_strm1_cntl          ( std__pe36__lane4_strm1_cntl       ),      
               .std__pe36__lane4_strm1_data          ( std__pe36__lane4_strm1_data       ),      
               .std__pe36__lane4_strm1_data_valid    ( std__pe36__lane4_strm1_data_valid ),      
               .std__pe36__lane4_strm1_data_mask     ( std__pe36__lane4_strm1_data_mask  ),      

               // PE 36, Lane 5                 
               .pe36__std__lane5_strm0_ready         ( pe36__std__lane5_strm0_ready      ),      
               .std__pe36__lane5_strm0_cntl          ( std__pe36__lane5_strm0_cntl       ),      
               .std__pe36__lane5_strm0_data          ( std__pe36__lane5_strm0_data       ),      
               .std__pe36__lane5_strm0_data_valid    ( std__pe36__lane5_strm0_data_valid ),      
               .std__pe36__lane5_strm0_data_mask     ( std__pe36__lane5_strm0_data_mask  ),      

               .pe36__std__lane5_strm1_ready         ( pe36__std__lane5_strm1_ready      ),      
               .std__pe36__lane5_strm1_cntl          ( std__pe36__lane5_strm1_cntl       ),      
               .std__pe36__lane5_strm1_data          ( std__pe36__lane5_strm1_data       ),      
               .std__pe36__lane5_strm1_data_valid    ( std__pe36__lane5_strm1_data_valid ),      
               .std__pe36__lane5_strm1_data_mask     ( std__pe36__lane5_strm1_data_mask  ),      

               // PE 36, Lane 6                 
               .pe36__std__lane6_strm0_ready         ( pe36__std__lane6_strm0_ready      ),      
               .std__pe36__lane6_strm0_cntl          ( std__pe36__lane6_strm0_cntl       ),      
               .std__pe36__lane6_strm0_data          ( std__pe36__lane6_strm0_data       ),      
               .std__pe36__lane6_strm0_data_valid    ( std__pe36__lane6_strm0_data_valid ),      
               .std__pe36__lane6_strm0_data_mask     ( std__pe36__lane6_strm0_data_mask  ),      

               .pe36__std__lane6_strm1_ready         ( pe36__std__lane6_strm1_ready      ),      
               .std__pe36__lane6_strm1_cntl          ( std__pe36__lane6_strm1_cntl       ),      
               .std__pe36__lane6_strm1_data          ( std__pe36__lane6_strm1_data       ),      
               .std__pe36__lane6_strm1_data_valid    ( std__pe36__lane6_strm1_data_valid ),      
               .std__pe36__lane6_strm1_data_mask     ( std__pe36__lane6_strm1_data_mask  ),      

               // PE 36, Lane 7                 
               .pe36__std__lane7_strm0_ready         ( pe36__std__lane7_strm0_ready      ),      
               .std__pe36__lane7_strm0_cntl          ( std__pe36__lane7_strm0_cntl       ),      
               .std__pe36__lane7_strm0_data          ( std__pe36__lane7_strm0_data       ),      
               .std__pe36__lane7_strm0_data_valid    ( std__pe36__lane7_strm0_data_valid ),      
               .std__pe36__lane7_strm0_data_mask     ( std__pe36__lane7_strm0_data_mask  ),      

               .pe36__std__lane7_strm1_ready         ( pe36__std__lane7_strm1_ready      ),      
               .std__pe36__lane7_strm1_cntl          ( std__pe36__lane7_strm1_cntl       ),      
               .std__pe36__lane7_strm1_data          ( std__pe36__lane7_strm1_data       ),      
               .std__pe36__lane7_strm1_data_valid    ( std__pe36__lane7_strm1_data_valid ),      
               .std__pe36__lane7_strm1_data_mask     ( std__pe36__lane7_strm1_data_mask  ),      

               // PE 36, Lane 8                 
               .pe36__std__lane8_strm0_ready         ( pe36__std__lane8_strm0_ready      ),      
               .std__pe36__lane8_strm0_cntl          ( std__pe36__lane8_strm0_cntl       ),      
               .std__pe36__lane8_strm0_data          ( std__pe36__lane8_strm0_data       ),      
               .std__pe36__lane8_strm0_data_valid    ( std__pe36__lane8_strm0_data_valid ),      
               .std__pe36__lane8_strm0_data_mask     ( std__pe36__lane8_strm0_data_mask  ),      

               .pe36__std__lane8_strm1_ready         ( pe36__std__lane8_strm1_ready      ),      
               .std__pe36__lane8_strm1_cntl          ( std__pe36__lane8_strm1_cntl       ),      
               .std__pe36__lane8_strm1_data          ( std__pe36__lane8_strm1_data       ),      
               .std__pe36__lane8_strm1_data_valid    ( std__pe36__lane8_strm1_data_valid ),      
               .std__pe36__lane8_strm1_data_mask     ( std__pe36__lane8_strm1_data_mask  ),      

               // PE 36, Lane 9                 
               .pe36__std__lane9_strm0_ready         ( pe36__std__lane9_strm0_ready      ),      
               .std__pe36__lane9_strm0_cntl          ( std__pe36__lane9_strm0_cntl       ),      
               .std__pe36__lane9_strm0_data          ( std__pe36__lane9_strm0_data       ),      
               .std__pe36__lane9_strm0_data_valid    ( std__pe36__lane9_strm0_data_valid ),      
               .std__pe36__lane9_strm0_data_mask     ( std__pe36__lane9_strm0_data_mask  ),      

               .pe36__std__lane9_strm1_ready         ( pe36__std__lane9_strm1_ready      ),      
               .std__pe36__lane9_strm1_cntl          ( std__pe36__lane9_strm1_cntl       ),      
               .std__pe36__lane9_strm1_data          ( std__pe36__lane9_strm1_data       ),      
               .std__pe36__lane9_strm1_data_valid    ( std__pe36__lane9_strm1_data_valid ),      
               .std__pe36__lane9_strm1_data_mask     ( std__pe36__lane9_strm1_data_mask  ),      

               // PE 36, Lane 10                 
               .pe36__std__lane10_strm0_ready         ( pe36__std__lane10_strm0_ready      ),      
               .std__pe36__lane10_strm0_cntl          ( std__pe36__lane10_strm0_cntl       ),      
               .std__pe36__lane10_strm0_data          ( std__pe36__lane10_strm0_data       ),      
               .std__pe36__lane10_strm0_data_valid    ( std__pe36__lane10_strm0_data_valid ),      
               .std__pe36__lane10_strm0_data_mask     ( std__pe36__lane10_strm0_data_mask  ),      

               .pe36__std__lane10_strm1_ready         ( pe36__std__lane10_strm1_ready      ),      
               .std__pe36__lane10_strm1_cntl          ( std__pe36__lane10_strm1_cntl       ),      
               .std__pe36__lane10_strm1_data          ( std__pe36__lane10_strm1_data       ),      
               .std__pe36__lane10_strm1_data_valid    ( std__pe36__lane10_strm1_data_valid ),      
               .std__pe36__lane10_strm1_data_mask     ( std__pe36__lane10_strm1_data_mask  ),      

               // PE 36, Lane 11                 
               .pe36__std__lane11_strm0_ready         ( pe36__std__lane11_strm0_ready      ),      
               .std__pe36__lane11_strm0_cntl          ( std__pe36__lane11_strm0_cntl       ),      
               .std__pe36__lane11_strm0_data          ( std__pe36__lane11_strm0_data       ),      
               .std__pe36__lane11_strm0_data_valid    ( std__pe36__lane11_strm0_data_valid ),      
               .std__pe36__lane11_strm0_data_mask     ( std__pe36__lane11_strm0_data_mask  ),      

               .pe36__std__lane11_strm1_ready         ( pe36__std__lane11_strm1_ready      ),      
               .std__pe36__lane11_strm1_cntl          ( std__pe36__lane11_strm1_cntl       ),      
               .std__pe36__lane11_strm1_data          ( std__pe36__lane11_strm1_data       ),      
               .std__pe36__lane11_strm1_data_valid    ( std__pe36__lane11_strm1_data_valid ),      
               .std__pe36__lane11_strm1_data_mask     ( std__pe36__lane11_strm1_data_mask  ),      

               // PE 36, Lane 12                 
               .pe36__std__lane12_strm0_ready         ( pe36__std__lane12_strm0_ready      ),      
               .std__pe36__lane12_strm0_cntl          ( std__pe36__lane12_strm0_cntl       ),      
               .std__pe36__lane12_strm0_data          ( std__pe36__lane12_strm0_data       ),      
               .std__pe36__lane12_strm0_data_valid    ( std__pe36__lane12_strm0_data_valid ),      
               .std__pe36__lane12_strm0_data_mask     ( std__pe36__lane12_strm0_data_mask  ),      

               .pe36__std__lane12_strm1_ready         ( pe36__std__lane12_strm1_ready      ),      
               .std__pe36__lane12_strm1_cntl          ( std__pe36__lane12_strm1_cntl       ),      
               .std__pe36__lane12_strm1_data          ( std__pe36__lane12_strm1_data       ),      
               .std__pe36__lane12_strm1_data_valid    ( std__pe36__lane12_strm1_data_valid ),      
               .std__pe36__lane12_strm1_data_mask     ( std__pe36__lane12_strm1_data_mask  ),      

               // PE 36, Lane 13                 
               .pe36__std__lane13_strm0_ready         ( pe36__std__lane13_strm0_ready      ),      
               .std__pe36__lane13_strm0_cntl          ( std__pe36__lane13_strm0_cntl       ),      
               .std__pe36__lane13_strm0_data          ( std__pe36__lane13_strm0_data       ),      
               .std__pe36__lane13_strm0_data_valid    ( std__pe36__lane13_strm0_data_valid ),      
               .std__pe36__lane13_strm0_data_mask     ( std__pe36__lane13_strm0_data_mask  ),      

               .pe36__std__lane13_strm1_ready         ( pe36__std__lane13_strm1_ready      ),      
               .std__pe36__lane13_strm1_cntl          ( std__pe36__lane13_strm1_cntl       ),      
               .std__pe36__lane13_strm1_data          ( std__pe36__lane13_strm1_data       ),      
               .std__pe36__lane13_strm1_data_valid    ( std__pe36__lane13_strm1_data_valid ),      
               .std__pe36__lane13_strm1_data_mask     ( std__pe36__lane13_strm1_data_mask  ),      

               // PE 36, Lane 14                 
               .pe36__std__lane14_strm0_ready         ( pe36__std__lane14_strm0_ready      ),      
               .std__pe36__lane14_strm0_cntl          ( std__pe36__lane14_strm0_cntl       ),      
               .std__pe36__lane14_strm0_data          ( std__pe36__lane14_strm0_data       ),      
               .std__pe36__lane14_strm0_data_valid    ( std__pe36__lane14_strm0_data_valid ),      
               .std__pe36__lane14_strm0_data_mask     ( std__pe36__lane14_strm0_data_mask  ),      

               .pe36__std__lane14_strm1_ready         ( pe36__std__lane14_strm1_ready      ),      
               .std__pe36__lane14_strm1_cntl          ( std__pe36__lane14_strm1_cntl       ),      
               .std__pe36__lane14_strm1_data          ( std__pe36__lane14_strm1_data       ),      
               .std__pe36__lane14_strm1_data_valid    ( std__pe36__lane14_strm1_data_valid ),      
               .std__pe36__lane14_strm1_data_mask     ( std__pe36__lane14_strm1_data_mask  ),      

               // PE 36, Lane 15                 
               .pe36__std__lane15_strm0_ready         ( pe36__std__lane15_strm0_ready      ),      
               .std__pe36__lane15_strm0_cntl          ( std__pe36__lane15_strm0_cntl       ),      
               .std__pe36__lane15_strm0_data          ( std__pe36__lane15_strm0_data       ),      
               .std__pe36__lane15_strm0_data_valid    ( std__pe36__lane15_strm0_data_valid ),      
               .std__pe36__lane15_strm0_data_mask     ( std__pe36__lane15_strm0_data_mask  ),      

               .pe36__std__lane15_strm1_ready         ( pe36__std__lane15_strm1_ready      ),      
               .std__pe36__lane15_strm1_cntl          ( std__pe36__lane15_strm1_cntl       ),      
               .std__pe36__lane15_strm1_data          ( std__pe36__lane15_strm1_data       ),      
               .std__pe36__lane15_strm1_data_valid    ( std__pe36__lane15_strm1_data_valid ),      
               .std__pe36__lane15_strm1_data_mask     ( std__pe36__lane15_strm1_data_mask  ),      

               // PE 36, Lane 16                 
               .pe36__std__lane16_strm0_ready         ( pe36__std__lane16_strm0_ready      ),      
               .std__pe36__lane16_strm0_cntl          ( std__pe36__lane16_strm0_cntl       ),      
               .std__pe36__lane16_strm0_data          ( std__pe36__lane16_strm0_data       ),      
               .std__pe36__lane16_strm0_data_valid    ( std__pe36__lane16_strm0_data_valid ),      
               .std__pe36__lane16_strm0_data_mask     ( std__pe36__lane16_strm0_data_mask  ),      

               .pe36__std__lane16_strm1_ready         ( pe36__std__lane16_strm1_ready      ),      
               .std__pe36__lane16_strm1_cntl          ( std__pe36__lane16_strm1_cntl       ),      
               .std__pe36__lane16_strm1_data          ( std__pe36__lane16_strm1_data       ),      
               .std__pe36__lane16_strm1_data_valid    ( std__pe36__lane16_strm1_data_valid ),      
               .std__pe36__lane16_strm1_data_mask     ( std__pe36__lane16_strm1_data_mask  ),      

               // PE 36, Lane 17                 
               .pe36__std__lane17_strm0_ready         ( pe36__std__lane17_strm0_ready      ),      
               .std__pe36__lane17_strm0_cntl          ( std__pe36__lane17_strm0_cntl       ),      
               .std__pe36__lane17_strm0_data          ( std__pe36__lane17_strm0_data       ),      
               .std__pe36__lane17_strm0_data_valid    ( std__pe36__lane17_strm0_data_valid ),      
               .std__pe36__lane17_strm0_data_mask     ( std__pe36__lane17_strm0_data_mask  ),      

               .pe36__std__lane17_strm1_ready         ( pe36__std__lane17_strm1_ready      ),      
               .std__pe36__lane17_strm1_cntl          ( std__pe36__lane17_strm1_cntl       ),      
               .std__pe36__lane17_strm1_data          ( std__pe36__lane17_strm1_data       ),      
               .std__pe36__lane17_strm1_data_valid    ( std__pe36__lane17_strm1_data_valid ),      
               .std__pe36__lane17_strm1_data_mask     ( std__pe36__lane17_strm1_data_mask  ),      

               // PE 36, Lane 18                 
               .pe36__std__lane18_strm0_ready         ( pe36__std__lane18_strm0_ready      ),      
               .std__pe36__lane18_strm0_cntl          ( std__pe36__lane18_strm0_cntl       ),      
               .std__pe36__lane18_strm0_data          ( std__pe36__lane18_strm0_data       ),      
               .std__pe36__lane18_strm0_data_valid    ( std__pe36__lane18_strm0_data_valid ),      
               .std__pe36__lane18_strm0_data_mask     ( std__pe36__lane18_strm0_data_mask  ),      

               .pe36__std__lane18_strm1_ready         ( pe36__std__lane18_strm1_ready      ),      
               .std__pe36__lane18_strm1_cntl          ( std__pe36__lane18_strm1_cntl       ),      
               .std__pe36__lane18_strm1_data          ( std__pe36__lane18_strm1_data       ),      
               .std__pe36__lane18_strm1_data_valid    ( std__pe36__lane18_strm1_data_valid ),      
               .std__pe36__lane18_strm1_data_mask     ( std__pe36__lane18_strm1_data_mask  ),      

               // PE 36, Lane 19                 
               .pe36__std__lane19_strm0_ready         ( pe36__std__lane19_strm0_ready      ),      
               .std__pe36__lane19_strm0_cntl          ( std__pe36__lane19_strm0_cntl       ),      
               .std__pe36__lane19_strm0_data          ( std__pe36__lane19_strm0_data       ),      
               .std__pe36__lane19_strm0_data_valid    ( std__pe36__lane19_strm0_data_valid ),      
               .std__pe36__lane19_strm0_data_mask     ( std__pe36__lane19_strm0_data_mask  ),      

               .pe36__std__lane19_strm1_ready         ( pe36__std__lane19_strm1_ready      ),      
               .std__pe36__lane19_strm1_cntl          ( std__pe36__lane19_strm1_cntl       ),      
               .std__pe36__lane19_strm1_data          ( std__pe36__lane19_strm1_data       ),      
               .std__pe36__lane19_strm1_data_valid    ( std__pe36__lane19_strm1_data_valid ),      
               .std__pe36__lane19_strm1_data_mask     ( std__pe36__lane19_strm1_data_mask  ),      

               // PE 36, Lane 20                 
               .pe36__std__lane20_strm0_ready         ( pe36__std__lane20_strm0_ready      ),      
               .std__pe36__lane20_strm0_cntl          ( std__pe36__lane20_strm0_cntl       ),      
               .std__pe36__lane20_strm0_data          ( std__pe36__lane20_strm0_data       ),      
               .std__pe36__lane20_strm0_data_valid    ( std__pe36__lane20_strm0_data_valid ),      
               .std__pe36__lane20_strm0_data_mask     ( std__pe36__lane20_strm0_data_mask  ),      

               .pe36__std__lane20_strm1_ready         ( pe36__std__lane20_strm1_ready      ),      
               .std__pe36__lane20_strm1_cntl          ( std__pe36__lane20_strm1_cntl       ),      
               .std__pe36__lane20_strm1_data          ( std__pe36__lane20_strm1_data       ),      
               .std__pe36__lane20_strm1_data_valid    ( std__pe36__lane20_strm1_data_valid ),      
               .std__pe36__lane20_strm1_data_mask     ( std__pe36__lane20_strm1_data_mask  ),      

               // PE 36, Lane 21                 
               .pe36__std__lane21_strm0_ready         ( pe36__std__lane21_strm0_ready      ),      
               .std__pe36__lane21_strm0_cntl          ( std__pe36__lane21_strm0_cntl       ),      
               .std__pe36__lane21_strm0_data          ( std__pe36__lane21_strm0_data       ),      
               .std__pe36__lane21_strm0_data_valid    ( std__pe36__lane21_strm0_data_valid ),      
               .std__pe36__lane21_strm0_data_mask     ( std__pe36__lane21_strm0_data_mask  ),      

               .pe36__std__lane21_strm1_ready         ( pe36__std__lane21_strm1_ready      ),      
               .std__pe36__lane21_strm1_cntl          ( std__pe36__lane21_strm1_cntl       ),      
               .std__pe36__lane21_strm1_data          ( std__pe36__lane21_strm1_data       ),      
               .std__pe36__lane21_strm1_data_valid    ( std__pe36__lane21_strm1_data_valid ),      
               .std__pe36__lane21_strm1_data_mask     ( std__pe36__lane21_strm1_data_mask  ),      

               // PE 36, Lane 22                 
               .pe36__std__lane22_strm0_ready         ( pe36__std__lane22_strm0_ready      ),      
               .std__pe36__lane22_strm0_cntl          ( std__pe36__lane22_strm0_cntl       ),      
               .std__pe36__lane22_strm0_data          ( std__pe36__lane22_strm0_data       ),      
               .std__pe36__lane22_strm0_data_valid    ( std__pe36__lane22_strm0_data_valid ),      
               .std__pe36__lane22_strm0_data_mask     ( std__pe36__lane22_strm0_data_mask  ),      

               .pe36__std__lane22_strm1_ready         ( pe36__std__lane22_strm1_ready      ),      
               .std__pe36__lane22_strm1_cntl          ( std__pe36__lane22_strm1_cntl       ),      
               .std__pe36__lane22_strm1_data          ( std__pe36__lane22_strm1_data       ),      
               .std__pe36__lane22_strm1_data_valid    ( std__pe36__lane22_strm1_data_valid ),      
               .std__pe36__lane22_strm1_data_mask     ( std__pe36__lane22_strm1_data_mask  ),      

               // PE 36, Lane 23                 
               .pe36__std__lane23_strm0_ready         ( pe36__std__lane23_strm0_ready      ),      
               .std__pe36__lane23_strm0_cntl          ( std__pe36__lane23_strm0_cntl       ),      
               .std__pe36__lane23_strm0_data          ( std__pe36__lane23_strm0_data       ),      
               .std__pe36__lane23_strm0_data_valid    ( std__pe36__lane23_strm0_data_valid ),      
               .std__pe36__lane23_strm0_data_mask     ( std__pe36__lane23_strm0_data_mask  ),      

               .pe36__std__lane23_strm1_ready         ( pe36__std__lane23_strm1_ready      ),      
               .std__pe36__lane23_strm1_cntl          ( std__pe36__lane23_strm1_cntl       ),      
               .std__pe36__lane23_strm1_data          ( std__pe36__lane23_strm1_data       ),      
               .std__pe36__lane23_strm1_data_valid    ( std__pe36__lane23_strm1_data_valid ),      
               .std__pe36__lane23_strm1_data_mask     ( std__pe36__lane23_strm1_data_mask  ),      

               // PE 36, Lane 24                 
               .pe36__std__lane24_strm0_ready         ( pe36__std__lane24_strm0_ready      ),      
               .std__pe36__lane24_strm0_cntl          ( std__pe36__lane24_strm0_cntl       ),      
               .std__pe36__lane24_strm0_data          ( std__pe36__lane24_strm0_data       ),      
               .std__pe36__lane24_strm0_data_valid    ( std__pe36__lane24_strm0_data_valid ),      
               .std__pe36__lane24_strm0_data_mask     ( std__pe36__lane24_strm0_data_mask  ),      

               .pe36__std__lane24_strm1_ready         ( pe36__std__lane24_strm1_ready      ),      
               .std__pe36__lane24_strm1_cntl          ( std__pe36__lane24_strm1_cntl       ),      
               .std__pe36__lane24_strm1_data          ( std__pe36__lane24_strm1_data       ),      
               .std__pe36__lane24_strm1_data_valid    ( std__pe36__lane24_strm1_data_valid ),      
               .std__pe36__lane24_strm1_data_mask     ( std__pe36__lane24_strm1_data_mask  ),      

               // PE 36, Lane 25                 
               .pe36__std__lane25_strm0_ready         ( pe36__std__lane25_strm0_ready      ),      
               .std__pe36__lane25_strm0_cntl          ( std__pe36__lane25_strm0_cntl       ),      
               .std__pe36__lane25_strm0_data          ( std__pe36__lane25_strm0_data       ),      
               .std__pe36__lane25_strm0_data_valid    ( std__pe36__lane25_strm0_data_valid ),      
               .std__pe36__lane25_strm0_data_mask     ( std__pe36__lane25_strm0_data_mask  ),      

               .pe36__std__lane25_strm1_ready         ( pe36__std__lane25_strm1_ready      ),      
               .std__pe36__lane25_strm1_cntl          ( std__pe36__lane25_strm1_cntl       ),      
               .std__pe36__lane25_strm1_data          ( std__pe36__lane25_strm1_data       ),      
               .std__pe36__lane25_strm1_data_valid    ( std__pe36__lane25_strm1_data_valid ),      
               .std__pe36__lane25_strm1_data_mask     ( std__pe36__lane25_strm1_data_mask  ),      

               // PE 36, Lane 26                 
               .pe36__std__lane26_strm0_ready         ( pe36__std__lane26_strm0_ready      ),      
               .std__pe36__lane26_strm0_cntl          ( std__pe36__lane26_strm0_cntl       ),      
               .std__pe36__lane26_strm0_data          ( std__pe36__lane26_strm0_data       ),      
               .std__pe36__lane26_strm0_data_valid    ( std__pe36__lane26_strm0_data_valid ),      
               .std__pe36__lane26_strm0_data_mask     ( std__pe36__lane26_strm0_data_mask  ),      

               .pe36__std__lane26_strm1_ready         ( pe36__std__lane26_strm1_ready      ),      
               .std__pe36__lane26_strm1_cntl          ( std__pe36__lane26_strm1_cntl       ),      
               .std__pe36__lane26_strm1_data          ( std__pe36__lane26_strm1_data       ),      
               .std__pe36__lane26_strm1_data_valid    ( std__pe36__lane26_strm1_data_valid ),      
               .std__pe36__lane26_strm1_data_mask     ( std__pe36__lane26_strm1_data_mask  ),      

               // PE 36, Lane 27                 
               .pe36__std__lane27_strm0_ready         ( pe36__std__lane27_strm0_ready      ),      
               .std__pe36__lane27_strm0_cntl          ( std__pe36__lane27_strm0_cntl       ),      
               .std__pe36__lane27_strm0_data          ( std__pe36__lane27_strm0_data       ),      
               .std__pe36__lane27_strm0_data_valid    ( std__pe36__lane27_strm0_data_valid ),      
               .std__pe36__lane27_strm0_data_mask     ( std__pe36__lane27_strm0_data_mask  ),      

               .pe36__std__lane27_strm1_ready         ( pe36__std__lane27_strm1_ready      ),      
               .std__pe36__lane27_strm1_cntl          ( std__pe36__lane27_strm1_cntl       ),      
               .std__pe36__lane27_strm1_data          ( std__pe36__lane27_strm1_data       ),      
               .std__pe36__lane27_strm1_data_valid    ( std__pe36__lane27_strm1_data_valid ),      
               .std__pe36__lane27_strm1_data_mask     ( std__pe36__lane27_strm1_data_mask  ),      

               // PE 36, Lane 28                 
               .pe36__std__lane28_strm0_ready         ( pe36__std__lane28_strm0_ready      ),      
               .std__pe36__lane28_strm0_cntl          ( std__pe36__lane28_strm0_cntl       ),      
               .std__pe36__lane28_strm0_data          ( std__pe36__lane28_strm0_data       ),      
               .std__pe36__lane28_strm0_data_valid    ( std__pe36__lane28_strm0_data_valid ),      
               .std__pe36__lane28_strm0_data_mask     ( std__pe36__lane28_strm0_data_mask  ),      

               .pe36__std__lane28_strm1_ready         ( pe36__std__lane28_strm1_ready      ),      
               .std__pe36__lane28_strm1_cntl          ( std__pe36__lane28_strm1_cntl       ),      
               .std__pe36__lane28_strm1_data          ( std__pe36__lane28_strm1_data       ),      
               .std__pe36__lane28_strm1_data_valid    ( std__pe36__lane28_strm1_data_valid ),      
               .std__pe36__lane28_strm1_data_mask     ( std__pe36__lane28_strm1_data_mask  ),      

               // PE 36, Lane 29                 
               .pe36__std__lane29_strm0_ready         ( pe36__std__lane29_strm0_ready      ),      
               .std__pe36__lane29_strm0_cntl          ( std__pe36__lane29_strm0_cntl       ),      
               .std__pe36__lane29_strm0_data          ( std__pe36__lane29_strm0_data       ),      
               .std__pe36__lane29_strm0_data_valid    ( std__pe36__lane29_strm0_data_valid ),      
               .std__pe36__lane29_strm0_data_mask     ( std__pe36__lane29_strm0_data_mask  ),      

               .pe36__std__lane29_strm1_ready         ( pe36__std__lane29_strm1_ready      ),      
               .std__pe36__lane29_strm1_cntl          ( std__pe36__lane29_strm1_cntl       ),      
               .std__pe36__lane29_strm1_data          ( std__pe36__lane29_strm1_data       ),      
               .std__pe36__lane29_strm1_data_valid    ( std__pe36__lane29_strm1_data_valid ),      
               .std__pe36__lane29_strm1_data_mask     ( std__pe36__lane29_strm1_data_mask  ),      

               // PE 36, Lane 30                 
               .pe36__std__lane30_strm0_ready         ( pe36__std__lane30_strm0_ready      ),      
               .std__pe36__lane30_strm0_cntl          ( std__pe36__lane30_strm0_cntl       ),      
               .std__pe36__lane30_strm0_data          ( std__pe36__lane30_strm0_data       ),      
               .std__pe36__lane30_strm0_data_valid    ( std__pe36__lane30_strm0_data_valid ),      
               .std__pe36__lane30_strm0_data_mask     ( std__pe36__lane30_strm0_data_mask  ),      

               .pe36__std__lane30_strm1_ready         ( pe36__std__lane30_strm1_ready      ),      
               .std__pe36__lane30_strm1_cntl          ( std__pe36__lane30_strm1_cntl       ),      
               .std__pe36__lane30_strm1_data          ( std__pe36__lane30_strm1_data       ),      
               .std__pe36__lane30_strm1_data_valid    ( std__pe36__lane30_strm1_data_valid ),      
               .std__pe36__lane30_strm1_data_mask     ( std__pe36__lane30_strm1_data_mask  ),      

               // PE 36, Lane 31                 
               .pe36__std__lane31_strm0_ready         ( pe36__std__lane31_strm0_ready      ),      
               .std__pe36__lane31_strm0_cntl          ( std__pe36__lane31_strm0_cntl       ),      
               .std__pe36__lane31_strm0_data          ( std__pe36__lane31_strm0_data       ),      
               .std__pe36__lane31_strm0_data_valid    ( std__pe36__lane31_strm0_data_valid ),      
               .std__pe36__lane31_strm0_data_mask     ( std__pe36__lane31_strm0_data_mask  ),      

               .pe36__std__lane31_strm1_ready         ( pe36__std__lane31_strm1_ready      ),      
               .std__pe36__lane31_strm1_cntl          ( std__pe36__lane31_strm1_cntl       ),      
               .std__pe36__lane31_strm1_data          ( std__pe36__lane31_strm1_data       ),      
               .std__pe36__lane31_strm1_data_valid    ( std__pe36__lane31_strm1_data_valid ),      
               .std__pe36__lane31_strm1_data_mask     ( std__pe36__lane31_strm1_data_mask  ),      

               // PE 37, Lane 0                 
               .pe37__std__lane0_strm0_ready         ( pe37__std__lane0_strm0_ready      ),      
               .std__pe37__lane0_strm0_cntl          ( std__pe37__lane0_strm0_cntl       ),      
               .std__pe37__lane0_strm0_data          ( std__pe37__lane0_strm0_data       ),      
               .std__pe37__lane0_strm0_data_valid    ( std__pe37__lane0_strm0_data_valid ),      
               .std__pe37__lane0_strm0_data_mask     ( std__pe37__lane0_strm0_data_mask  ),      

               .pe37__std__lane0_strm1_ready         ( pe37__std__lane0_strm1_ready      ),      
               .std__pe37__lane0_strm1_cntl          ( std__pe37__lane0_strm1_cntl       ),      
               .std__pe37__lane0_strm1_data          ( std__pe37__lane0_strm1_data       ),      
               .std__pe37__lane0_strm1_data_valid    ( std__pe37__lane0_strm1_data_valid ),      
               .std__pe37__lane0_strm1_data_mask     ( std__pe37__lane0_strm1_data_mask  ),      

               // PE 37, Lane 1                 
               .pe37__std__lane1_strm0_ready         ( pe37__std__lane1_strm0_ready      ),      
               .std__pe37__lane1_strm0_cntl          ( std__pe37__lane1_strm0_cntl       ),      
               .std__pe37__lane1_strm0_data          ( std__pe37__lane1_strm0_data       ),      
               .std__pe37__lane1_strm0_data_valid    ( std__pe37__lane1_strm0_data_valid ),      
               .std__pe37__lane1_strm0_data_mask     ( std__pe37__lane1_strm0_data_mask  ),      

               .pe37__std__lane1_strm1_ready         ( pe37__std__lane1_strm1_ready      ),      
               .std__pe37__lane1_strm1_cntl          ( std__pe37__lane1_strm1_cntl       ),      
               .std__pe37__lane1_strm1_data          ( std__pe37__lane1_strm1_data       ),      
               .std__pe37__lane1_strm1_data_valid    ( std__pe37__lane1_strm1_data_valid ),      
               .std__pe37__lane1_strm1_data_mask     ( std__pe37__lane1_strm1_data_mask  ),      

               // PE 37, Lane 2                 
               .pe37__std__lane2_strm0_ready         ( pe37__std__lane2_strm0_ready      ),      
               .std__pe37__lane2_strm0_cntl          ( std__pe37__lane2_strm0_cntl       ),      
               .std__pe37__lane2_strm0_data          ( std__pe37__lane2_strm0_data       ),      
               .std__pe37__lane2_strm0_data_valid    ( std__pe37__lane2_strm0_data_valid ),      
               .std__pe37__lane2_strm0_data_mask     ( std__pe37__lane2_strm0_data_mask  ),      

               .pe37__std__lane2_strm1_ready         ( pe37__std__lane2_strm1_ready      ),      
               .std__pe37__lane2_strm1_cntl          ( std__pe37__lane2_strm1_cntl       ),      
               .std__pe37__lane2_strm1_data          ( std__pe37__lane2_strm1_data       ),      
               .std__pe37__lane2_strm1_data_valid    ( std__pe37__lane2_strm1_data_valid ),      
               .std__pe37__lane2_strm1_data_mask     ( std__pe37__lane2_strm1_data_mask  ),      

               // PE 37, Lane 3                 
               .pe37__std__lane3_strm0_ready         ( pe37__std__lane3_strm0_ready      ),      
               .std__pe37__lane3_strm0_cntl          ( std__pe37__lane3_strm0_cntl       ),      
               .std__pe37__lane3_strm0_data          ( std__pe37__lane3_strm0_data       ),      
               .std__pe37__lane3_strm0_data_valid    ( std__pe37__lane3_strm0_data_valid ),      
               .std__pe37__lane3_strm0_data_mask     ( std__pe37__lane3_strm0_data_mask  ),      

               .pe37__std__lane3_strm1_ready         ( pe37__std__lane3_strm1_ready      ),      
               .std__pe37__lane3_strm1_cntl          ( std__pe37__lane3_strm1_cntl       ),      
               .std__pe37__lane3_strm1_data          ( std__pe37__lane3_strm1_data       ),      
               .std__pe37__lane3_strm1_data_valid    ( std__pe37__lane3_strm1_data_valid ),      
               .std__pe37__lane3_strm1_data_mask     ( std__pe37__lane3_strm1_data_mask  ),      

               // PE 37, Lane 4                 
               .pe37__std__lane4_strm0_ready         ( pe37__std__lane4_strm0_ready      ),      
               .std__pe37__lane4_strm0_cntl          ( std__pe37__lane4_strm0_cntl       ),      
               .std__pe37__lane4_strm0_data          ( std__pe37__lane4_strm0_data       ),      
               .std__pe37__lane4_strm0_data_valid    ( std__pe37__lane4_strm0_data_valid ),      
               .std__pe37__lane4_strm0_data_mask     ( std__pe37__lane4_strm0_data_mask  ),      

               .pe37__std__lane4_strm1_ready         ( pe37__std__lane4_strm1_ready      ),      
               .std__pe37__lane4_strm1_cntl          ( std__pe37__lane4_strm1_cntl       ),      
               .std__pe37__lane4_strm1_data          ( std__pe37__lane4_strm1_data       ),      
               .std__pe37__lane4_strm1_data_valid    ( std__pe37__lane4_strm1_data_valid ),      
               .std__pe37__lane4_strm1_data_mask     ( std__pe37__lane4_strm1_data_mask  ),      

               // PE 37, Lane 5                 
               .pe37__std__lane5_strm0_ready         ( pe37__std__lane5_strm0_ready      ),      
               .std__pe37__lane5_strm0_cntl          ( std__pe37__lane5_strm0_cntl       ),      
               .std__pe37__lane5_strm0_data          ( std__pe37__lane5_strm0_data       ),      
               .std__pe37__lane5_strm0_data_valid    ( std__pe37__lane5_strm0_data_valid ),      
               .std__pe37__lane5_strm0_data_mask     ( std__pe37__lane5_strm0_data_mask  ),      

               .pe37__std__lane5_strm1_ready         ( pe37__std__lane5_strm1_ready      ),      
               .std__pe37__lane5_strm1_cntl          ( std__pe37__lane5_strm1_cntl       ),      
               .std__pe37__lane5_strm1_data          ( std__pe37__lane5_strm1_data       ),      
               .std__pe37__lane5_strm1_data_valid    ( std__pe37__lane5_strm1_data_valid ),      
               .std__pe37__lane5_strm1_data_mask     ( std__pe37__lane5_strm1_data_mask  ),      

               // PE 37, Lane 6                 
               .pe37__std__lane6_strm0_ready         ( pe37__std__lane6_strm0_ready      ),      
               .std__pe37__lane6_strm0_cntl          ( std__pe37__lane6_strm0_cntl       ),      
               .std__pe37__lane6_strm0_data          ( std__pe37__lane6_strm0_data       ),      
               .std__pe37__lane6_strm0_data_valid    ( std__pe37__lane6_strm0_data_valid ),      
               .std__pe37__lane6_strm0_data_mask     ( std__pe37__lane6_strm0_data_mask  ),      

               .pe37__std__lane6_strm1_ready         ( pe37__std__lane6_strm1_ready      ),      
               .std__pe37__lane6_strm1_cntl          ( std__pe37__lane6_strm1_cntl       ),      
               .std__pe37__lane6_strm1_data          ( std__pe37__lane6_strm1_data       ),      
               .std__pe37__lane6_strm1_data_valid    ( std__pe37__lane6_strm1_data_valid ),      
               .std__pe37__lane6_strm1_data_mask     ( std__pe37__lane6_strm1_data_mask  ),      

               // PE 37, Lane 7                 
               .pe37__std__lane7_strm0_ready         ( pe37__std__lane7_strm0_ready      ),      
               .std__pe37__lane7_strm0_cntl          ( std__pe37__lane7_strm0_cntl       ),      
               .std__pe37__lane7_strm0_data          ( std__pe37__lane7_strm0_data       ),      
               .std__pe37__lane7_strm0_data_valid    ( std__pe37__lane7_strm0_data_valid ),      
               .std__pe37__lane7_strm0_data_mask     ( std__pe37__lane7_strm0_data_mask  ),      

               .pe37__std__lane7_strm1_ready         ( pe37__std__lane7_strm1_ready      ),      
               .std__pe37__lane7_strm1_cntl          ( std__pe37__lane7_strm1_cntl       ),      
               .std__pe37__lane7_strm1_data          ( std__pe37__lane7_strm1_data       ),      
               .std__pe37__lane7_strm1_data_valid    ( std__pe37__lane7_strm1_data_valid ),      
               .std__pe37__lane7_strm1_data_mask     ( std__pe37__lane7_strm1_data_mask  ),      

               // PE 37, Lane 8                 
               .pe37__std__lane8_strm0_ready         ( pe37__std__lane8_strm0_ready      ),      
               .std__pe37__lane8_strm0_cntl          ( std__pe37__lane8_strm0_cntl       ),      
               .std__pe37__lane8_strm0_data          ( std__pe37__lane8_strm0_data       ),      
               .std__pe37__lane8_strm0_data_valid    ( std__pe37__lane8_strm0_data_valid ),      
               .std__pe37__lane8_strm0_data_mask     ( std__pe37__lane8_strm0_data_mask  ),      

               .pe37__std__lane8_strm1_ready         ( pe37__std__lane8_strm1_ready      ),      
               .std__pe37__lane8_strm1_cntl          ( std__pe37__lane8_strm1_cntl       ),      
               .std__pe37__lane8_strm1_data          ( std__pe37__lane8_strm1_data       ),      
               .std__pe37__lane8_strm1_data_valid    ( std__pe37__lane8_strm1_data_valid ),      
               .std__pe37__lane8_strm1_data_mask     ( std__pe37__lane8_strm1_data_mask  ),      

               // PE 37, Lane 9                 
               .pe37__std__lane9_strm0_ready         ( pe37__std__lane9_strm0_ready      ),      
               .std__pe37__lane9_strm0_cntl          ( std__pe37__lane9_strm0_cntl       ),      
               .std__pe37__lane9_strm0_data          ( std__pe37__lane9_strm0_data       ),      
               .std__pe37__lane9_strm0_data_valid    ( std__pe37__lane9_strm0_data_valid ),      
               .std__pe37__lane9_strm0_data_mask     ( std__pe37__lane9_strm0_data_mask  ),      

               .pe37__std__lane9_strm1_ready         ( pe37__std__lane9_strm1_ready      ),      
               .std__pe37__lane9_strm1_cntl          ( std__pe37__lane9_strm1_cntl       ),      
               .std__pe37__lane9_strm1_data          ( std__pe37__lane9_strm1_data       ),      
               .std__pe37__lane9_strm1_data_valid    ( std__pe37__lane9_strm1_data_valid ),      
               .std__pe37__lane9_strm1_data_mask     ( std__pe37__lane9_strm1_data_mask  ),      

               // PE 37, Lane 10                 
               .pe37__std__lane10_strm0_ready         ( pe37__std__lane10_strm0_ready      ),      
               .std__pe37__lane10_strm0_cntl          ( std__pe37__lane10_strm0_cntl       ),      
               .std__pe37__lane10_strm0_data          ( std__pe37__lane10_strm0_data       ),      
               .std__pe37__lane10_strm0_data_valid    ( std__pe37__lane10_strm0_data_valid ),      
               .std__pe37__lane10_strm0_data_mask     ( std__pe37__lane10_strm0_data_mask  ),      

               .pe37__std__lane10_strm1_ready         ( pe37__std__lane10_strm1_ready      ),      
               .std__pe37__lane10_strm1_cntl          ( std__pe37__lane10_strm1_cntl       ),      
               .std__pe37__lane10_strm1_data          ( std__pe37__lane10_strm1_data       ),      
               .std__pe37__lane10_strm1_data_valid    ( std__pe37__lane10_strm1_data_valid ),      
               .std__pe37__lane10_strm1_data_mask     ( std__pe37__lane10_strm1_data_mask  ),      

               // PE 37, Lane 11                 
               .pe37__std__lane11_strm0_ready         ( pe37__std__lane11_strm0_ready      ),      
               .std__pe37__lane11_strm0_cntl          ( std__pe37__lane11_strm0_cntl       ),      
               .std__pe37__lane11_strm0_data          ( std__pe37__lane11_strm0_data       ),      
               .std__pe37__lane11_strm0_data_valid    ( std__pe37__lane11_strm0_data_valid ),      
               .std__pe37__lane11_strm0_data_mask     ( std__pe37__lane11_strm0_data_mask  ),      

               .pe37__std__lane11_strm1_ready         ( pe37__std__lane11_strm1_ready      ),      
               .std__pe37__lane11_strm1_cntl          ( std__pe37__lane11_strm1_cntl       ),      
               .std__pe37__lane11_strm1_data          ( std__pe37__lane11_strm1_data       ),      
               .std__pe37__lane11_strm1_data_valid    ( std__pe37__lane11_strm1_data_valid ),      
               .std__pe37__lane11_strm1_data_mask     ( std__pe37__lane11_strm1_data_mask  ),      

               // PE 37, Lane 12                 
               .pe37__std__lane12_strm0_ready         ( pe37__std__lane12_strm0_ready      ),      
               .std__pe37__lane12_strm0_cntl          ( std__pe37__lane12_strm0_cntl       ),      
               .std__pe37__lane12_strm0_data          ( std__pe37__lane12_strm0_data       ),      
               .std__pe37__lane12_strm0_data_valid    ( std__pe37__lane12_strm0_data_valid ),      
               .std__pe37__lane12_strm0_data_mask     ( std__pe37__lane12_strm0_data_mask  ),      

               .pe37__std__lane12_strm1_ready         ( pe37__std__lane12_strm1_ready      ),      
               .std__pe37__lane12_strm1_cntl          ( std__pe37__lane12_strm1_cntl       ),      
               .std__pe37__lane12_strm1_data          ( std__pe37__lane12_strm1_data       ),      
               .std__pe37__lane12_strm1_data_valid    ( std__pe37__lane12_strm1_data_valid ),      
               .std__pe37__lane12_strm1_data_mask     ( std__pe37__lane12_strm1_data_mask  ),      

               // PE 37, Lane 13                 
               .pe37__std__lane13_strm0_ready         ( pe37__std__lane13_strm0_ready      ),      
               .std__pe37__lane13_strm0_cntl          ( std__pe37__lane13_strm0_cntl       ),      
               .std__pe37__lane13_strm0_data          ( std__pe37__lane13_strm0_data       ),      
               .std__pe37__lane13_strm0_data_valid    ( std__pe37__lane13_strm0_data_valid ),      
               .std__pe37__lane13_strm0_data_mask     ( std__pe37__lane13_strm0_data_mask  ),      

               .pe37__std__lane13_strm1_ready         ( pe37__std__lane13_strm1_ready      ),      
               .std__pe37__lane13_strm1_cntl          ( std__pe37__lane13_strm1_cntl       ),      
               .std__pe37__lane13_strm1_data          ( std__pe37__lane13_strm1_data       ),      
               .std__pe37__lane13_strm1_data_valid    ( std__pe37__lane13_strm1_data_valid ),      
               .std__pe37__lane13_strm1_data_mask     ( std__pe37__lane13_strm1_data_mask  ),      

               // PE 37, Lane 14                 
               .pe37__std__lane14_strm0_ready         ( pe37__std__lane14_strm0_ready      ),      
               .std__pe37__lane14_strm0_cntl          ( std__pe37__lane14_strm0_cntl       ),      
               .std__pe37__lane14_strm0_data          ( std__pe37__lane14_strm0_data       ),      
               .std__pe37__lane14_strm0_data_valid    ( std__pe37__lane14_strm0_data_valid ),      
               .std__pe37__lane14_strm0_data_mask     ( std__pe37__lane14_strm0_data_mask  ),      

               .pe37__std__lane14_strm1_ready         ( pe37__std__lane14_strm1_ready      ),      
               .std__pe37__lane14_strm1_cntl          ( std__pe37__lane14_strm1_cntl       ),      
               .std__pe37__lane14_strm1_data          ( std__pe37__lane14_strm1_data       ),      
               .std__pe37__lane14_strm1_data_valid    ( std__pe37__lane14_strm1_data_valid ),      
               .std__pe37__lane14_strm1_data_mask     ( std__pe37__lane14_strm1_data_mask  ),      

               // PE 37, Lane 15                 
               .pe37__std__lane15_strm0_ready         ( pe37__std__lane15_strm0_ready      ),      
               .std__pe37__lane15_strm0_cntl          ( std__pe37__lane15_strm0_cntl       ),      
               .std__pe37__lane15_strm0_data          ( std__pe37__lane15_strm0_data       ),      
               .std__pe37__lane15_strm0_data_valid    ( std__pe37__lane15_strm0_data_valid ),      
               .std__pe37__lane15_strm0_data_mask     ( std__pe37__lane15_strm0_data_mask  ),      

               .pe37__std__lane15_strm1_ready         ( pe37__std__lane15_strm1_ready      ),      
               .std__pe37__lane15_strm1_cntl          ( std__pe37__lane15_strm1_cntl       ),      
               .std__pe37__lane15_strm1_data          ( std__pe37__lane15_strm1_data       ),      
               .std__pe37__lane15_strm1_data_valid    ( std__pe37__lane15_strm1_data_valid ),      
               .std__pe37__lane15_strm1_data_mask     ( std__pe37__lane15_strm1_data_mask  ),      

               // PE 37, Lane 16                 
               .pe37__std__lane16_strm0_ready         ( pe37__std__lane16_strm0_ready      ),      
               .std__pe37__lane16_strm0_cntl          ( std__pe37__lane16_strm0_cntl       ),      
               .std__pe37__lane16_strm0_data          ( std__pe37__lane16_strm0_data       ),      
               .std__pe37__lane16_strm0_data_valid    ( std__pe37__lane16_strm0_data_valid ),      
               .std__pe37__lane16_strm0_data_mask     ( std__pe37__lane16_strm0_data_mask  ),      

               .pe37__std__lane16_strm1_ready         ( pe37__std__lane16_strm1_ready      ),      
               .std__pe37__lane16_strm1_cntl          ( std__pe37__lane16_strm1_cntl       ),      
               .std__pe37__lane16_strm1_data          ( std__pe37__lane16_strm1_data       ),      
               .std__pe37__lane16_strm1_data_valid    ( std__pe37__lane16_strm1_data_valid ),      
               .std__pe37__lane16_strm1_data_mask     ( std__pe37__lane16_strm1_data_mask  ),      

               // PE 37, Lane 17                 
               .pe37__std__lane17_strm0_ready         ( pe37__std__lane17_strm0_ready      ),      
               .std__pe37__lane17_strm0_cntl          ( std__pe37__lane17_strm0_cntl       ),      
               .std__pe37__lane17_strm0_data          ( std__pe37__lane17_strm0_data       ),      
               .std__pe37__lane17_strm0_data_valid    ( std__pe37__lane17_strm0_data_valid ),      
               .std__pe37__lane17_strm0_data_mask     ( std__pe37__lane17_strm0_data_mask  ),      

               .pe37__std__lane17_strm1_ready         ( pe37__std__lane17_strm1_ready      ),      
               .std__pe37__lane17_strm1_cntl          ( std__pe37__lane17_strm1_cntl       ),      
               .std__pe37__lane17_strm1_data          ( std__pe37__lane17_strm1_data       ),      
               .std__pe37__lane17_strm1_data_valid    ( std__pe37__lane17_strm1_data_valid ),      
               .std__pe37__lane17_strm1_data_mask     ( std__pe37__lane17_strm1_data_mask  ),      

               // PE 37, Lane 18                 
               .pe37__std__lane18_strm0_ready         ( pe37__std__lane18_strm0_ready      ),      
               .std__pe37__lane18_strm0_cntl          ( std__pe37__lane18_strm0_cntl       ),      
               .std__pe37__lane18_strm0_data          ( std__pe37__lane18_strm0_data       ),      
               .std__pe37__lane18_strm0_data_valid    ( std__pe37__lane18_strm0_data_valid ),      
               .std__pe37__lane18_strm0_data_mask     ( std__pe37__lane18_strm0_data_mask  ),      

               .pe37__std__lane18_strm1_ready         ( pe37__std__lane18_strm1_ready      ),      
               .std__pe37__lane18_strm1_cntl          ( std__pe37__lane18_strm1_cntl       ),      
               .std__pe37__lane18_strm1_data          ( std__pe37__lane18_strm1_data       ),      
               .std__pe37__lane18_strm1_data_valid    ( std__pe37__lane18_strm1_data_valid ),      
               .std__pe37__lane18_strm1_data_mask     ( std__pe37__lane18_strm1_data_mask  ),      

               // PE 37, Lane 19                 
               .pe37__std__lane19_strm0_ready         ( pe37__std__lane19_strm0_ready      ),      
               .std__pe37__lane19_strm0_cntl          ( std__pe37__lane19_strm0_cntl       ),      
               .std__pe37__lane19_strm0_data          ( std__pe37__lane19_strm0_data       ),      
               .std__pe37__lane19_strm0_data_valid    ( std__pe37__lane19_strm0_data_valid ),      
               .std__pe37__lane19_strm0_data_mask     ( std__pe37__lane19_strm0_data_mask  ),      

               .pe37__std__lane19_strm1_ready         ( pe37__std__lane19_strm1_ready      ),      
               .std__pe37__lane19_strm1_cntl          ( std__pe37__lane19_strm1_cntl       ),      
               .std__pe37__lane19_strm1_data          ( std__pe37__lane19_strm1_data       ),      
               .std__pe37__lane19_strm1_data_valid    ( std__pe37__lane19_strm1_data_valid ),      
               .std__pe37__lane19_strm1_data_mask     ( std__pe37__lane19_strm1_data_mask  ),      

               // PE 37, Lane 20                 
               .pe37__std__lane20_strm0_ready         ( pe37__std__lane20_strm0_ready      ),      
               .std__pe37__lane20_strm0_cntl          ( std__pe37__lane20_strm0_cntl       ),      
               .std__pe37__lane20_strm0_data          ( std__pe37__lane20_strm0_data       ),      
               .std__pe37__lane20_strm0_data_valid    ( std__pe37__lane20_strm0_data_valid ),      
               .std__pe37__lane20_strm0_data_mask     ( std__pe37__lane20_strm0_data_mask  ),      

               .pe37__std__lane20_strm1_ready         ( pe37__std__lane20_strm1_ready      ),      
               .std__pe37__lane20_strm1_cntl          ( std__pe37__lane20_strm1_cntl       ),      
               .std__pe37__lane20_strm1_data          ( std__pe37__lane20_strm1_data       ),      
               .std__pe37__lane20_strm1_data_valid    ( std__pe37__lane20_strm1_data_valid ),      
               .std__pe37__lane20_strm1_data_mask     ( std__pe37__lane20_strm1_data_mask  ),      

               // PE 37, Lane 21                 
               .pe37__std__lane21_strm0_ready         ( pe37__std__lane21_strm0_ready      ),      
               .std__pe37__lane21_strm0_cntl          ( std__pe37__lane21_strm0_cntl       ),      
               .std__pe37__lane21_strm0_data          ( std__pe37__lane21_strm0_data       ),      
               .std__pe37__lane21_strm0_data_valid    ( std__pe37__lane21_strm0_data_valid ),      
               .std__pe37__lane21_strm0_data_mask     ( std__pe37__lane21_strm0_data_mask  ),      

               .pe37__std__lane21_strm1_ready         ( pe37__std__lane21_strm1_ready      ),      
               .std__pe37__lane21_strm1_cntl          ( std__pe37__lane21_strm1_cntl       ),      
               .std__pe37__lane21_strm1_data          ( std__pe37__lane21_strm1_data       ),      
               .std__pe37__lane21_strm1_data_valid    ( std__pe37__lane21_strm1_data_valid ),      
               .std__pe37__lane21_strm1_data_mask     ( std__pe37__lane21_strm1_data_mask  ),      

               // PE 37, Lane 22                 
               .pe37__std__lane22_strm0_ready         ( pe37__std__lane22_strm0_ready      ),      
               .std__pe37__lane22_strm0_cntl          ( std__pe37__lane22_strm0_cntl       ),      
               .std__pe37__lane22_strm0_data          ( std__pe37__lane22_strm0_data       ),      
               .std__pe37__lane22_strm0_data_valid    ( std__pe37__lane22_strm0_data_valid ),      
               .std__pe37__lane22_strm0_data_mask     ( std__pe37__lane22_strm0_data_mask  ),      

               .pe37__std__lane22_strm1_ready         ( pe37__std__lane22_strm1_ready      ),      
               .std__pe37__lane22_strm1_cntl          ( std__pe37__lane22_strm1_cntl       ),      
               .std__pe37__lane22_strm1_data          ( std__pe37__lane22_strm1_data       ),      
               .std__pe37__lane22_strm1_data_valid    ( std__pe37__lane22_strm1_data_valid ),      
               .std__pe37__lane22_strm1_data_mask     ( std__pe37__lane22_strm1_data_mask  ),      

               // PE 37, Lane 23                 
               .pe37__std__lane23_strm0_ready         ( pe37__std__lane23_strm0_ready      ),      
               .std__pe37__lane23_strm0_cntl          ( std__pe37__lane23_strm0_cntl       ),      
               .std__pe37__lane23_strm0_data          ( std__pe37__lane23_strm0_data       ),      
               .std__pe37__lane23_strm0_data_valid    ( std__pe37__lane23_strm0_data_valid ),      
               .std__pe37__lane23_strm0_data_mask     ( std__pe37__lane23_strm0_data_mask  ),      

               .pe37__std__lane23_strm1_ready         ( pe37__std__lane23_strm1_ready      ),      
               .std__pe37__lane23_strm1_cntl          ( std__pe37__lane23_strm1_cntl       ),      
               .std__pe37__lane23_strm1_data          ( std__pe37__lane23_strm1_data       ),      
               .std__pe37__lane23_strm1_data_valid    ( std__pe37__lane23_strm1_data_valid ),      
               .std__pe37__lane23_strm1_data_mask     ( std__pe37__lane23_strm1_data_mask  ),      

               // PE 37, Lane 24                 
               .pe37__std__lane24_strm0_ready         ( pe37__std__lane24_strm0_ready      ),      
               .std__pe37__lane24_strm0_cntl          ( std__pe37__lane24_strm0_cntl       ),      
               .std__pe37__lane24_strm0_data          ( std__pe37__lane24_strm0_data       ),      
               .std__pe37__lane24_strm0_data_valid    ( std__pe37__lane24_strm0_data_valid ),      
               .std__pe37__lane24_strm0_data_mask     ( std__pe37__lane24_strm0_data_mask  ),      

               .pe37__std__lane24_strm1_ready         ( pe37__std__lane24_strm1_ready      ),      
               .std__pe37__lane24_strm1_cntl          ( std__pe37__lane24_strm1_cntl       ),      
               .std__pe37__lane24_strm1_data          ( std__pe37__lane24_strm1_data       ),      
               .std__pe37__lane24_strm1_data_valid    ( std__pe37__lane24_strm1_data_valid ),      
               .std__pe37__lane24_strm1_data_mask     ( std__pe37__lane24_strm1_data_mask  ),      

               // PE 37, Lane 25                 
               .pe37__std__lane25_strm0_ready         ( pe37__std__lane25_strm0_ready      ),      
               .std__pe37__lane25_strm0_cntl          ( std__pe37__lane25_strm0_cntl       ),      
               .std__pe37__lane25_strm0_data          ( std__pe37__lane25_strm0_data       ),      
               .std__pe37__lane25_strm0_data_valid    ( std__pe37__lane25_strm0_data_valid ),      
               .std__pe37__lane25_strm0_data_mask     ( std__pe37__lane25_strm0_data_mask  ),      

               .pe37__std__lane25_strm1_ready         ( pe37__std__lane25_strm1_ready      ),      
               .std__pe37__lane25_strm1_cntl          ( std__pe37__lane25_strm1_cntl       ),      
               .std__pe37__lane25_strm1_data          ( std__pe37__lane25_strm1_data       ),      
               .std__pe37__lane25_strm1_data_valid    ( std__pe37__lane25_strm1_data_valid ),      
               .std__pe37__lane25_strm1_data_mask     ( std__pe37__lane25_strm1_data_mask  ),      

               // PE 37, Lane 26                 
               .pe37__std__lane26_strm0_ready         ( pe37__std__lane26_strm0_ready      ),      
               .std__pe37__lane26_strm0_cntl          ( std__pe37__lane26_strm0_cntl       ),      
               .std__pe37__lane26_strm0_data          ( std__pe37__lane26_strm0_data       ),      
               .std__pe37__lane26_strm0_data_valid    ( std__pe37__lane26_strm0_data_valid ),      
               .std__pe37__lane26_strm0_data_mask     ( std__pe37__lane26_strm0_data_mask  ),      

               .pe37__std__lane26_strm1_ready         ( pe37__std__lane26_strm1_ready      ),      
               .std__pe37__lane26_strm1_cntl          ( std__pe37__lane26_strm1_cntl       ),      
               .std__pe37__lane26_strm1_data          ( std__pe37__lane26_strm1_data       ),      
               .std__pe37__lane26_strm1_data_valid    ( std__pe37__lane26_strm1_data_valid ),      
               .std__pe37__lane26_strm1_data_mask     ( std__pe37__lane26_strm1_data_mask  ),      

               // PE 37, Lane 27                 
               .pe37__std__lane27_strm0_ready         ( pe37__std__lane27_strm0_ready      ),      
               .std__pe37__lane27_strm0_cntl          ( std__pe37__lane27_strm0_cntl       ),      
               .std__pe37__lane27_strm0_data          ( std__pe37__lane27_strm0_data       ),      
               .std__pe37__lane27_strm0_data_valid    ( std__pe37__lane27_strm0_data_valid ),      
               .std__pe37__lane27_strm0_data_mask     ( std__pe37__lane27_strm0_data_mask  ),      

               .pe37__std__lane27_strm1_ready         ( pe37__std__lane27_strm1_ready      ),      
               .std__pe37__lane27_strm1_cntl          ( std__pe37__lane27_strm1_cntl       ),      
               .std__pe37__lane27_strm1_data          ( std__pe37__lane27_strm1_data       ),      
               .std__pe37__lane27_strm1_data_valid    ( std__pe37__lane27_strm1_data_valid ),      
               .std__pe37__lane27_strm1_data_mask     ( std__pe37__lane27_strm1_data_mask  ),      

               // PE 37, Lane 28                 
               .pe37__std__lane28_strm0_ready         ( pe37__std__lane28_strm0_ready      ),      
               .std__pe37__lane28_strm0_cntl          ( std__pe37__lane28_strm0_cntl       ),      
               .std__pe37__lane28_strm0_data          ( std__pe37__lane28_strm0_data       ),      
               .std__pe37__lane28_strm0_data_valid    ( std__pe37__lane28_strm0_data_valid ),      
               .std__pe37__lane28_strm0_data_mask     ( std__pe37__lane28_strm0_data_mask  ),      

               .pe37__std__lane28_strm1_ready         ( pe37__std__lane28_strm1_ready      ),      
               .std__pe37__lane28_strm1_cntl          ( std__pe37__lane28_strm1_cntl       ),      
               .std__pe37__lane28_strm1_data          ( std__pe37__lane28_strm1_data       ),      
               .std__pe37__lane28_strm1_data_valid    ( std__pe37__lane28_strm1_data_valid ),      
               .std__pe37__lane28_strm1_data_mask     ( std__pe37__lane28_strm1_data_mask  ),      

               // PE 37, Lane 29                 
               .pe37__std__lane29_strm0_ready         ( pe37__std__lane29_strm0_ready      ),      
               .std__pe37__lane29_strm0_cntl          ( std__pe37__lane29_strm0_cntl       ),      
               .std__pe37__lane29_strm0_data          ( std__pe37__lane29_strm0_data       ),      
               .std__pe37__lane29_strm0_data_valid    ( std__pe37__lane29_strm0_data_valid ),      
               .std__pe37__lane29_strm0_data_mask     ( std__pe37__lane29_strm0_data_mask  ),      

               .pe37__std__lane29_strm1_ready         ( pe37__std__lane29_strm1_ready      ),      
               .std__pe37__lane29_strm1_cntl          ( std__pe37__lane29_strm1_cntl       ),      
               .std__pe37__lane29_strm1_data          ( std__pe37__lane29_strm1_data       ),      
               .std__pe37__lane29_strm1_data_valid    ( std__pe37__lane29_strm1_data_valid ),      
               .std__pe37__lane29_strm1_data_mask     ( std__pe37__lane29_strm1_data_mask  ),      

               // PE 37, Lane 30                 
               .pe37__std__lane30_strm0_ready         ( pe37__std__lane30_strm0_ready      ),      
               .std__pe37__lane30_strm0_cntl          ( std__pe37__lane30_strm0_cntl       ),      
               .std__pe37__lane30_strm0_data          ( std__pe37__lane30_strm0_data       ),      
               .std__pe37__lane30_strm0_data_valid    ( std__pe37__lane30_strm0_data_valid ),      
               .std__pe37__lane30_strm0_data_mask     ( std__pe37__lane30_strm0_data_mask  ),      

               .pe37__std__lane30_strm1_ready         ( pe37__std__lane30_strm1_ready      ),      
               .std__pe37__lane30_strm1_cntl          ( std__pe37__lane30_strm1_cntl       ),      
               .std__pe37__lane30_strm1_data          ( std__pe37__lane30_strm1_data       ),      
               .std__pe37__lane30_strm1_data_valid    ( std__pe37__lane30_strm1_data_valid ),      
               .std__pe37__lane30_strm1_data_mask     ( std__pe37__lane30_strm1_data_mask  ),      

               // PE 37, Lane 31                 
               .pe37__std__lane31_strm0_ready         ( pe37__std__lane31_strm0_ready      ),      
               .std__pe37__lane31_strm0_cntl          ( std__pe37__lane31_strm0_cntl       ),      
               .std__pe37__lane31_strm0_data          ( std__pe37__lane31_strm0_data       ),      
               .std__pe37__lane31_strm0_data_valid    ( std__pe37__lane31_strm0_data_valid ),      
               .std__pe37__lane31_strm0_data_mask     ( std__pe37__lane31_strm0_data_mask  ),      

               .pe37__std__lane31_strm1_ready         ( pe37__std__lane31_strm1_ready      ),      
               .std__pe37__lane31_strm1_cntl          ( std__pe37__lane31_strm1_cntl       ),      
               .std__pe37__lane31_strm1_data          ( std__pe37__lane31_strm1_data       ),      
               .std__pe37__lane31_strm1_data_valid    ( std__pe37__lane31_strm1_data_valid ),      
               .std__pe37__lane31_strm1_data_mask     ( std__pe37__lane31_strm1_data_mask  ),      

               // PE 38, Lane 0                 
               .pe38__std__lane0_strm0_ready         ( pe38__std__lane0_strm0_ready      ),      
               .std__pe38__lane0_strm0_cntl          ( std__pe38__lane0_strm0_cntl       ),      
               .std__pe38__lane0_strm0_data          ( std__pe38__lane0_strm0_data       ),      
               .std__pe38__lane0_strm0_data_valid    ( std__pe38__lane0_strm0_data_valid ),      
               .std__pe38__lane0_strm0_data_mask     ( std__pe38__lane0_strm0_data_mask  ),      

               .pe38__std__lane0_strm1_ready         ( pe38__std__lane0_strm1_ready      ),      
               .std__pe38__lane0_strm1_cntl          ( std__pe38__lane0_strm1_cntl       ),      
               .std__pe38__lane0_strm1_data          ( std__pe38__lane0_strm1_data       ),      
               .std__pe38__lane0_strm1_data_valid    ( std__pe38__lane0_strm1_data_valid ),      
               .std__pe38__lane0_strm1_data_mask     ( std__pe38__lane0_strm1_data_mask  ),      

               // PE 38, Lane 1                 
               .pe38__std__lane1_strm0_ready         ( pe38__std__lane1_strm0_ready      ),      
               .std__pe38__lane1_strm0_cntl          ( std__pe38__lane1_strm0_cntl       ),      
               .std__pe38__lane1_strm0_data          ( std__pe38__lane1_strm0_data       ),      
               .std__pe38__lane1_strm0_data_valid    ( std__pe38__lane1_strm0_data_valid ),      
               .std__pe38__lane1_strm0_data_mask     ( std__pe38__lane1_strm0_data_mask  ),      

               .pe38__std__lane1_strm1_ready         ( pe38__std__lane1_strm1_ready      ),      
               .std__pe38__lane1_strm1_cntl          ( std__pe38__lane1_strm1_cntl       ),      
               .std__pe38__lane1_strm1_data          ( std__pe38__lane1_strm1_data       ),      
               .std__pe38__lane1_strm1_data_valid    ( std__pe38__lane1_strm1_data_valid ),      
               .std__pe38__lane1_strm1_data_mask     ( std__pe38__lane1_strm1_data_mask  ),      

               // PE 38, Lane 2                 
               .pe38__std__lane2_strm0_ready         ( pe38__std__lane2_strm0_ready      ),      
               .std__pe38__lane2_strm0_cntl          ( std__pe38__lane2_strm0_cntl       ),      
               .std__pe38__lane2_strm0_data          ( std__pe38__lane2_strm0_data       ),      
               .std__pe38__lane2_strm0_data_valid    ( std__pe38__lane2_strm0_data_valid ),      
               .std__pe38__lane2_strm0_data_mask     ( std__pe38__lane2_strm0_data_mask  ),      

               .pe38__std__lane2_strm1_ready         ( pe38__std__lane2_strm1_ready      ),      
               .std__pe38__lane2_strm1_cntl          ( std__pe38__lane2_strm1_cntl       ),      
               .std__pe38__lane2_strm1_data          ( std__pe38__lane2_strm1_data       ),      
               .std__pe38__lane2_strm1_data_valid    ( std__pe38__lane2_strm1_data_valid ),      
               .std__pe38__lane2_strm1_data_mask     ( std__pe38__lane2_strm1_data_mask  ),      

               // PE 38, Lane 3                 
               .pe38__std__lane3_strm0_ready         ( pe38__std__lane3_strm0_ready      ),      
               .std__pe38__lane3_strm0_cntl          ( std__pe38__lane3_strm0_cntl       ),      
               .std__pe38__lane3_strm0_data          ( std__pe38__lane3_strm0_data       ),      
               .std__pe38__lane3_strm0_data_valid    ( std__pe38__lane3_strm0_data_valid ),      
               .std__pe38__lane3_strm0_data_mask     ( std__pe38__lane3_strm0_data_mask  ),      

               .pe38__std__lane3_strm1_ready         ( pe38__std__lane3_strm1_ready      ),      
               .std__pe38__lane3_strm1_cntl          ( std__pe38__lane3_strm1_cntl       ),      
               .std__pe38__lane3_strm1_data          ( std__pe38__lane3_strm1_data       ),      
               .std__pe38__lane3_strm1_data_valid    ( std__pe38__lane3_strm1_data_valid ),      
               .std__pe38__lane3_strm1_data_mask     ( std__pe38__lane3_strm1_data_mask  ),      

               // PE 38, Lane 4                 
               .pe38__std__lane4_strm0_ready         ( pe38__std__lane4_strm0_ready      ),      
               .std__pe38__lane4_strm0_cntl          ( std__pe38__lane4_strm0_cntl       ),      
               .std__pe38__lane4_strm0_data          ( std__pe38__lane4_strm0_data       ),      
               .std__pe38__lane4_strm0_data_valid    ( std__pe38__lane4_strm0_data_valid ),      
               .std__pe38__lane4_strm0_data_mask     ( std__pe38__lane4_strm0_data_mask  ),      

               .pe38__std__lane4_strm1_ready         ( pe38__std__lane4_strm1_ready      ),      
               .std__pe38__lane4_strm1_cntl          ( std__pe38__lane4_strm1_cntl       ),      
               .std__pe38__lane4_strm1_data          ( std__pe38__lane4_strm1_data       ),      
               .std__pe38__lane4_strm1_data_valid    ( std__pe38__lane4_strm1_data_valid ),      
               .std__pe38__lane4_strm1_data_mask     ( std__pe38__lane4_strm1_data_mask  ),      

               // PE 38, Lane 5                 
               .pe38__std__lane5_strm0_ready         ( pe38__std__lane5_strm0_ready      ),      
               .std__pe38__lane5_strm0_cntl          ( std__pe38__lane5_strm0_cntl       ),      
               .std__pe38__lane5_strm0_data          ( std__pe38__lane5_strm0_data       ),      
               .std__pe38__lane5_strm0_data_valid    ( std__pe38__lane5_strm0_data_valid ),      
               .std__pe38__lane5_strm0_data_mask     ( std__pe38__lane5_strm0_data_mask  ),      

               .pe38__std__lane5_strm1_ready         ( pe38__std__lane5_strm1_ready      ),      
               .std__pe38__lane5_strm1_cntl          ( std__pe38__lane5_strm1_cntl       ),      
               .std__pe38__lane5_strm1_data          ( std__pe38__lane5_strm1_data       ),      
               .std__pe38__lane5_strm1_data_valid    ( std__pe38__lane5_strm1_data_valid ),      
               .std__pe38__lane5_strm1_data_mask     ( std__pe38__lane5_strm1_data_mask  ),      

               // PE 38, Lane 6                 
               .pe38__std__lane6_strm0_ready         ( pe38__std__lane6_strm0_ready      ),      
               .std__pe38__lane6_strm0_cntl          ( std__pe38__lane6_strm0_cntl       ),      
               .std__pe38__lane6_strm0_data          ( std__pe38__lane6_strm0_data       ),      
               .std__pe38__lane6_strm0_data_valid    ( std__pe38__lane6_strm0_data_valid ),      
               .std__pe38__lane6_strm0_data_mask     ( std__pe38__lane6_strm0_data_mask  ),      

               .pe38__std__lane6_strm1_ready         ( pe38__std__lane6_strm1_ready      ),      
               .std__pe38__lane6_strm1_cntl          ( std__pe38__lane6_strm1_cntl       ),      
               .std__pe38__lane6_strm1_data          ( std__pe38__lane6_strm1_data       ),      
               .std__pe38__lane6_strm1_data_valid    ( std__pe38__lane6_strm1_data_valid ),      
               .std__pe38__lane6_strm1_data_mask     ( std__pe38__lane6_strm1_data_mask  ),      

               // PE 38, Lane 7                 
               .pe38__std__lane7_strm0_ready         ( pe38__std__lane7_strm0_ready      ),      
               .std__pe38__lane7_strm0_cntl          ( std__pe38__lane7_strm0_cntl       ),      
               .std__pe38__lane7_strm0_data          ( std__pe38__lane7_strm0_data       ),      
               .std__pe38__lane7_strm0_data_valid    ( std__pe38__lane7_strm0_data_valid ),      
               .std__pe38__lane7_strm0_data_mask     ( std__pe38__lane7_strm0_data_mask  ),      

               .pe38__std__lane7_strm1_ready         ( pe38__std__lane7_strm1_ready      ),      
               .std__pe38__lane7_strm1_cntl          ( std__pe38__lane7_strm1_cntl       ),      
               .std__pe38__lane7_strm1_data          ( std__pe38__lane7_strm1_data       ),      
               .std__pe38__lane7_strm1_data_valid    ( std__pe38__lane7_strm1_data_valid ),      
               .std__pe38__lane7_strm1_data_mask     ( std__pe38__lane7_strm1_data_mask  ),      

               // PE 38, Lane 8                 
               .pe38__std__lane8_strm0_ready         ( pe38__std__lane8_strm0_ready      ),      
               .std__pe38__lane8_strm0_cntl          ( std__pe38__lane8_strm0_cntl       ),      
               .std__pe38__lane8_strm0_data          ( std__pe38__lane8_strm0_data       ),      
               .std__pe38__lane8_strm0_data_valid    ( std__pe38__lane8_strm0_data_valid ),      
               .std__pe38__lane8_strm0_data_mask     ( std__pe38__lane8_strm0_data_mask  ),      

               .pe38__std__lane8_strm1_ready         ( pe38__std__lane8_strm1_ready      ),      
               .std__pe38__lane8_strm1_cntl          ( std__pe38__lane8_strm1_cntl       ),      
               .std__pe38__lane8_strm1_data          ( std__pe38__lane8_strm1_data       ),      
               .std__pe38__lane8_strm1_data_valid    ( std__pe38__lane8_strm1_data_valid ),      
               .std__pe38__lane8_strm1_data_mask     ( std__pe38__lane8_strm1_data_mask  ),      

               // PE 38, Lane 9                 
               .pe38__std__lane9_strm0_ready         ( pe38__std__lane9_strm0_ready      ),      
               .std__pe38__lane9_strm0_cntl          ( std__pe38__lane9_strm0_cntl       ),      
               .std__pe38__lane9_strm0_data          ( std__pe38__lane9_strm0_data       ),      
               .std__pe38__lane9_strm0_data_valid    ( std__pe38__lane9_strm0_data_valid ),      
               .std__pe38__lane9_strm0_data_mask     ( std__pe38__lane9_strm0_data_mask  ),      

               .pe38__std__lane9_strm1_ready         ( pe38__std__lane9_strm1_ready      ),      
               .std__pe38__lane9_strm1_cntl          ( std__pe38__lane9_strm1_cntl       ),      
               .std__pe38__lane9_strm1_data          ( std__pe38__lane9_strm1_data       ),      
               .std__pe38__lane9_strm1_data_valid    ( std__pe38__lane9_strm1_data_valid ),      
               .std__pe38__lane9_strm1_data_mask     ( std__pe38__lane9_strm1_data_mask  ),      

               // PE 38, Lane 10                 
               .pe38__std__lane10_strm0_ready         ( pe38__std__lane10_strm0_ready      ),      
               .std__pe38__lane10_strm0_cntl          ( std__pe38__lane10_strm0_cntl       ),      
               .std__pe38__lane10_strm0_data          ( std__pe38__lane10_strm0_data       ),      
               .std__pe38__lane10_strm0_data_valid    ( std__pe38__lane10_strm0_data_valid ),      
               .std__pe38__lane10_strm0_data_mask     ( std__pe38__lane10_strm0_data_mask  ),      

               .pe38__std__lane10_strm1_ready         ( pe38__std__lane10_strm1_ready      ),      
               .std__pe38__lane10_strm1_cntl          ( std__pe38__lane10_strm1_cntl       ),      
               .std__pe38__lane10_strm1_data          ( std__pe38__lane10_strm1_data       ),      
               .std__pe38__lane10_strm1_data_valid    ( std__pe38__lane10_strm1_data_valid ),      
               .std__pe38__lane10_strm1_data_mask     ( std__pe38__lane10_strm1_data_mask  ),      

               // PE 38, Lane 11                 
               .pe38__std__lane11_strm0_ready         ( pe38__std__lane11_strm0_ready      ),      
               .std__pe38__lane11_strm0_cntl          ( std__pe38__lane11_strm0_cntl       ),      
               .std__pe38__lane11_strm0_data          ( std__pe38__lane11_strm0_data       ),      
               .std__pe38__lane11_strm0_data_valid    ( std__pe38__lane11_strm0_data_valid ),      
               .std__pe38__lane11_strm0_data_mask     ( std__pe38__lane11_strm0_data_mask  ),      

               .pe38__std__lane11_strm1_ready         ( pe38__std__lane11_strm1_ready      ),      
               .std__pe38__lane11_strm1_cntl          ( std__pe38__lane11_strm1_cntl       ),      
               .std__pe38__lane11_strm1_data          ( std__pe38__lane11_strm1_data       ),      
               .std__pe38__lane11_strm1_data_valid    ( std__pe38__lane11_strm1_data_valid ),      
               .std__pe38__lane11_strm1_data_mask     ( std__pe38__lane11_strm1_data_mask  ),      

               // PE 38, Lane 12                 
               .pe38__std__lane12_strm0_ready         ( pe38__std__lane12_strm0_ready      ),      
               .std__pe38__lane12_strm0_cntl          ( std__pe38__lane12_strm0_cntl       ),      
               .std__pe38__lane12_strm0_data          ( std__pe38__lane12_strm0_data       ),      
               .std__pe38__lane12_strm0_data_valid    ( std__pe38__lane12_strm0_data_valid ),      
               .std__pe38__lane12_strm0_data_mask     ( std__pe38__lane12_strm0_data_mask  ),      

               .pe38__std__lane12_strm1_ready         ( pe38__std__lane12_strm1_ready      ),      
               .std__pe38__lane12_strm1_cntl          ( std__pe38__lane12_strm1_cntl       ),      
               .std__pe38__lane12_strm1_data          ( std__pe38__lane12_strm1_data       ),      
               .std__pe38__lane12_strm1_data_valid    ( std__pe38__lane12_strm1_data_valid ),      
               .std__pe38__lane12_strm1_data_mask     ( std__pe38__lane12_strm1_data_mask  ),      

               // PE 38, Lane 13                 
               .pe38__std__lane13_strm0_ready         ( pe38__std__lane13_strm0_ready      ),      
               .std__pe38__lane13_strm0_cntl          ( std__pe38__lane13_strm0_cntl       ),      
               .std__pe38__lane13_strm0_data          ( std__pe38__lane13_strm0_data       ),      
               .std__pe38__lane13_strm0_data_valid    ( std__pe38__lane13_strm0_data_valid ),      
               .std__pe38__lane13_strm0_data_mask     ( std__pe38__lane13_strm0_data_mask  ),      

               .pe38__std__lane13_strm1_ready         ( pe38__std__lane13_strm1_ready      ),      
               .std__pe38__lane13_strm1_cntl          ( std__pe38__lane13_strm1_cntl       ),      
               .std__pe38__lane13_strm1_data          ( std__pe38__lane13_strm1_data       ),      
               .std__pe38__lane13_strm1_data_valid    ( std__pe38__lane13_strm1_data_valid ),      
               .std__pe38__lane13_strm1_data_mask     ( std__pe38__lane13_strm1_data_mask  ),      

               // PE 38, Lane 14                 
               .pe38__std__lane14_strm0_ready         ( pe38__std__lane14_strm0_ready      ),      
               .std__pe38__lane14_strm0_cntl          ( std__pe38__lane14_strm0_cntl       ),      
               .std__pe38__lane14_strm0_data          ( std__pe38__lane14_strm0_data       ),      
               .std__pe38__lane14_strm0_data_valid    ( std__pe38__lane14_strm0_data_valid ),      
               .std__pe38__lane14_strm0_data_mask     ( std__pe38__lane14_strm0_data_mask  ),      

               .pe38__std__lane14_strm1_ready         ( pe38__std__lane14_strm1_ready      ),      
               .std__pe38__lane14_strm1_cntl          ( std__pe38__lane14_strm1_cntl       ),      
               .std__pe38__lane14_strm1_data          ( std__pe38__lane14_strm1_data       ),      
               .std__pe38__lane14_strm1_data_valid    ( std__pe38__lane14_strm1_data_valid ),      
               .std__pe38__lane14_strm1_data_mask     ( std__pe38__lane14_strm1_data_mask  ),      

               // PE 38, Lane 15                 
               .pe38__std__lane15_strm0_ready         ( pe38__std__lane15_strm0_ready      ),      
               .std__pe38__lane15_strm0_cntl          ( std__pe38__lane15_strm0_cntl       ),      
               .std__pe38__lane15_strm0_data          ( std__pe38__lane15_strm0_data       ),      
               .std__pe38__lane15_strm0_data_valid    ( std__pe38__lane15_strm0_data_valid ),      
               .std__pe38__lane15_strm0_data_mask     ( std__pe38__lane15_strm0_data_mask  ),      

               .pe38__std__lane15_strm1_ready         ( pe38__std__lane15_strm1_ready      ),      
               .std__pe38__lane15_strm1_cntl          ( std__pe38__lane15_strm1_cntl       ),      
               .std__pe38__lane15_strm1_data          ( std__pe38__lane15_strm1_data       ),      
               .std__pe38__lane15_strm1_data_valid    ( std__pe38__lane15_strm1_data_valid ),      
               .std__pe38__lane15_strm1_data_mask     ( std__pe38__lane15_strm1_data_mask  ),      

               // PE 38, Lane 16                 
               .pe38__std__lane16_strm0_ready         ( pe38__std__lane16_strm0_ready      ),      
               .std__pe38__lane16_strm0_cntl          ( std__pe38__lane16_strm0_cntl       ),      
               .std__pe38__lane16_strm0_data          ( std__pe38__lane16_strm0_data       ),      
               .std__pe38__lane16_strm0_data_valid    ( std__pe38__lane16_strm0_data_valid ),      
               .std__pe38__lane16_strm0_data_mask     ( std__pe38__lane16_strm0_data_mask  ),      

               .pe38__std__lane16_strm1_ready         ( pe38__std__lane16_strm1_ready      ),      
               .std__pe38__lane16_strm1_cntl          ( std__pe38__lane16_strm1_cntl       ),      
               .std__pe38__lane16_strm1_data          ( std__pe38__lane16_strm1_data       ),      
               .std__pe38__lane16_strm1_data_valid    ( std__pe38__lane16_strm1_data_valid ),      
               .std__pe38__lane16_strm1_data_mask     ( std__pe38__lane16_strm1_data_mask  ),      

               // PE 38, Lane 17                 
               .pe38__std__lane17_strm0_ready         ( pe38__std__lane17_strm0_ready      ),      
               .std__pe38__lane17_strm0_cntl          ( std__pe38__lane17_strm0_cntl       ),      
               .std__pe38__lane17_strm0_data          ( std__pe38__lane17_strm0_data       ),      
               .std__pe38__lane17_strm0_data_valid    ( std__pe38__lane17_strm0_data_valid ),      
               .std__pe38__lane17_strm0_data_mask     ( std__pe38__lane17_strm0_data_mask  ),      

               .pe38__std__lane17_strm1_ready         ( pe38__std__lane17_strm1_ready      ),      
               .std__pe38__lane17_strm1_cntl          ( std__pe38__lane17_strm1_cntl       ),      
               .std__pe38__lane17_strm1_data          ( std__pe38__lane17_strm1_data       ),      
               .std__pe38__lane17_strm1_data_valid    ( std__pe38__lane17_strm1_data_valid ),      
               .std__pe38__lane17_strm1_data_mask     ( std__pe38__lane17_strm1_data_mask  ),      

               // PE 38, Lane 18                 
               .pe38__std__lane18_strm0_ready         ( pe38__std__lane18_strm0_ready      ),      
               .std__pe38__lane18_strm0_cntl          ( std__pe38__lane18_strm0_cntl       ),      
               .std__pe38__lane18_strm0_data          ( std__pe38__lane18_strm0_data       ),      
               .std__pe38__lane18_strm0_data_valid    ( std__pe38__lane18_strm0_data_valid ),      
               .std__pe38__lane18_strm0_data_mask     ( std__pe38__lane18_strm0_data_mask  ),      

               .pe38__std__lane18_strm1_ready         ( pe38__std__lane18_strm1_ready      ),      
               .std__pe38__lane18_strm1_cntl          ( std__pe38__lane18_strm1_cntl       ),      
               .std__pe38__lane18_strm1_data          ( std__pe38__lane18_strm1_data       ),      
               .std__pe38__lane18_strm1_data_valid    ( std__pe38__lane18_strm1_data_valid ),      
               .std__pe38__lane18_strm1_data_mask     ( std__pe38__lane18_strm1_data_mask  ),      

               // PE 38, Lane 19                 
               .pe38__std__lane19_strm0_ready         ( pe38__std__lane19_strm0_ready      ),      
               .std__pe38__lane19_strm0_cntl          ( std__pe38__lane19_strm0_cntl       ),      
               .std__pe38__lane19_strm0_data          ( std__pe38__lane19_strm0_data       ),      
               .std__pe38__lane19_strm0_data_valid    ( std__pe38__lane19_strm0_data_valid ),      
               .std__pe38__lane19_strm0_data_mask     ( std__pe38__lane19_strm0_data_mask  ),      

               .pe38__std__lane19_strm1_ready         ( pe38__std__lane19_strm1_ready      ),      
               .std__pe38__lane19_strm1_cntl          ( std__pe38__lane19_strm1_cntl       ),      
               .std__pe38__lane19_strm1_data          ( std__pe38__lane19_strm1_data       ),      
               .std__pe38__lane19_strm1_data_valid    ( std__pe38__lane19_strm1_data_valid ),      
               .std__pe38__lane19_strm1_data_mask     ( std__pe38__lane19_strm1_data_mask  ),      

               // PE 38, Lane 20                 
               .pe38__std__lane20_strm0_ready         ( pe38__std__lane20_strm0_ready      ),      
               .std__pe38__lane20_strm0_cntl          ( std__pe38__lane20_strm0_cntl       ),      
               .std__pe38__lane20_strm0_data          ( std__pe38__lane20_strm0_data       ),      
               .std__pe38__lane20_strm0_data_valid    ( std__pe38__lane20_strm0_data_valid ),      
               .std__pe38__lane20_strm0_data_mask     ( std__pe38__lane20_strm0_data_mask  ),      

               .pe38__std__lane20_strm1_ready         ( pe38__std__lane20_strm1_ready      ),      
               .std__pe38__lane20_strm1_cntl          ( std__pe38__lane20_strm1_cntl       ),      
               .std__pe38__lane20_strm1_data          ( std__pe38__lane20_strm1_data       ),      
               .std__pe38__lane20_strm1_data_valid    ( std__pe38__lane20_strm1_data_valid ),      
               .std__pe38__lane20_strm1_data_mask     ( std__pe38__lane20_strm1_data_mask  ),      

               // PE 38, Lane 21                 
               .pe38__std__lane21_strm0_ready         ( pe38__std__lane21_strm0_ready      ),      
               .std__pe38__lane21_strm0_cntl          ( std__pe38__lane21_strm0_cntl       ),      
               .std__pe38__lane21_strm0_data          ( std__pe38__lane21_strm0_data       ),      
               .std__pe38__lane21_strm0_data_valid    ( std__pe38__lane21_strm0_data_valid ),      
               .std__pe38__lane21_strm0_data_mask     ( std__pe38__lane21_strm0_data_mask  ),      

               .pe38__std__lane21_strm1_ready         ( pe38__std__lane21_strm1_ready      ),      
               .std__pe38__lane21_strm1_cntl          ( std__pe38__lane21_strm1_cntl       ),      
               .std__pe38__lane21_strm1_data          ( std__pe38__lane21_strm1_data       ),      
               .std__pe38__lane21_strm1_data_valid    ( std__pe38__lane21_strm1_data_valid ),      
               .std__pe38__lane21_strm1_data_mask     ( std__pe38__lane21_strm1_data_mask  ),      

               // PE 38, Lane 22                 
               .pe38__std__lane22_strm0_ready         ( pe38__std__lane22_strm0_ready      ),      
               .std__pe38__lane22_strm0_cntl          ( std__pe38__lane22_strm0_cntl       ),      
               .std__pe38__lane22_strm0_data          ( std__pe38__lane22_strm0_data       ),      
               .std__pe38__lane22_strm0_data_valid    ( std__pe38__lane22_strm0_data_valid ),      
               .std__pe38__lane22_strm0_data_mask     ( std__pe38__lane22_strm0_data_mask  ),      

               .pe38__std__lane22_strm1_ready         ( pe38__std__lane22_strm1_ready      ),      
               .std__pe38__lane22_strm1_cntl          ( std__pe38__lane22_strm1_cntl       ),      
               .std__pe38__lane22_strm1_data          ( std__pe38__lane22_strm1_data       ),      
               .std__pe38__lane22_strm1_data_valid    ( std__pe38__lane22_strm1_data_valid ),      
               .std__pe38__lane22_strm1_data_mask     ( std__pe38__lane22_strm1_data_mask  ),      

               // PE 38, Lane 23                 
               .pe38__std__lane23_strm0_ready         ( pe38__std__lane23_strm0_ready      ),      
               .std__pe38__lane23_strm0_cntl          ( std__pe38__lane23_strm0_cntl       ),      
               .std__pe38__lane23_strm0_data          ( std__pe38__lane23_strm0_data       ),      
               .std__pe38__lane23_strm0_data_valid    ( std__pe38__lane23_strm0_data_valid ),      
               .std__pe38__lane23_strm0_data_mask     ( std__pe38__lane23_strm0_data_mask  ),      

               .pe38__std__lane23_strm1_ready         ( pe38__std__lane23_strm1_ready      ),      
               .std__pe38__lane23_strm1_cntl          ( std__pe38__lane23_strm1_cntl       ),      
               .std__pe38__lane23_strm1_data          ( std__pe38__lane23_strm1_data       ),      
               .std__pe38__lane23_strm1_data_valid    ( std__pe38__lane23_strm1_data_valid ),      
               .std__pe38__lane23_strm1_data_mask     ( std__pe38__lane23_strm1_data_mask  ),      

               // PE 38, Lane 24                 
               .pe38__std__lane24_strm0_ready         ( pe38__std__lane24_strm0_ready      ),      
               .std__pe38__lane24_strm0_cntl          ( std__pe38__lane24_strm0_cntl       ),      
               .std__pe38__lane24_strm0_data          ( std__pe38__lane24_strm0_data       ),      
               .std__pe38__lane24_strm0_data_valid    ( std__pe38__lane24_strm0_data_valid ),      
               .std__pe38__lane24_strm0_data_mask     ( std__pe38__lane24_strm0_data_mask  ),      

               .pe38__std__lane24_strm1_ready         ( pe38__std__lane24_strm1_ready      ),      
               .std__pe38__lane24_strm1_cntl          ( std__pe38__lane24_strm1_cntl       ),      
               .std__pe38__lane24_strm1_data          ( std__pe38__lane24_strm1_data       ),      
               .std__pe38__lane24_strm1_data_valid    ( std__pe38__lane24_strm1_data_valid ),      
               .std__pe38__lane24_strm1_data_mask     ( std__pe38__lane24_strm1_data_mask  ),      

               // PE 38, Lane 25                 
               .pe38__std__lane25_strm0_ready         ( pe38__std__lane25_strm0_ready      ),      
               .std__pe38__lane25_strm0_cntl          ( std__pe38__lane25_strm0_cntl       ),      
               .std__pe38__lane25_strm0_data          ( std__pe38__lane25_strm0_data       ),      
               .std__pe38__lane25_strm0_data_valid    ( std__pe38__lane25_strm0_data_valid ),      
               .std__pe38__lane25_strm0_data_mask     ( std__pe38__lane25_strm0_data_mask  ),      

               .pe38__std__lane25_strm1_ready         ( pe38__std__lane25_strm1_ready      ),      
               .std__pe38__lane25_strm1_cntl          ( std__pe38__lane25_strm1_cntl       ),      
               .std__pe38__lane25_strm1_data          ( std__pe38__lane25_strm1_data       ),      
               .std__pe38__lane25_strm1_data_valid    ( std__pe38__lane25_strm1_data_valid ),      
               .std__pe38__lane25_strm1_data_mask     ( std__pe38__lane25_strm1_data_mask  ),      

               // PE 38, Lane 26                 
               .pe38__std__lane26_strm0_ready         ( pe38__std__lane26_strm0_ready      ),      
               .std__pe38__lane26_strm0_cntl          ( std__pe38__lane26_strm0_cntl       ),      
               .std__pe38__lane26_strm0_data          ( std__pe38__lane26_strm0_data       ),      
               .std__pe38__lane26_strm0_data_valid    ( std__pe38__lane26_strm0_data_valid ),      
               .std__pe38__lane26_strm0_data_mask     ( std__pe38__lane26_strm0_data_mask  ),      

               .pe38__std__lane26_strm1_ready         ( pe38__std__lane26_strm1_ready      ),      
               .std__pe38__lane26_strm1_cntl          ( std__pe38__lane26_strm1_cntl       ),      
               .std__pe38__lane26_strm1_data          ( std__pe38__lane26_strm1_data       ),      
               .std__pe38__lane26_strm1_data_valid    ( std__pe38__lane26_strm1_data_valid ),      
               .std__pe38__lane26_strm1_data_mask     ( std__pe38__lane26_strm1_data_mask  ),      

               // PE 38, Lane 27                 
               .pe38__std__lane27_strm0_ready         ( pe38__std__lane27_strm0_ready      ),      
               .std__pe38__lane27_strm0_cntl          ( std__pe38__lane27_strm0_cntl       ),      
               .std__pe38__lane27_strm0_data          ( std__pe38__lane27_strm0_data       ),      
               .std__pe38__lane27_strm0_data_valid    ( std__pe38__lane27_strm0_data_valid ),      
               .std__pe38__lane27_strm0_data_mask     ( std__pe38__lane27_strm0_data_mask  ),      

               .pe38__std__lane27_strm1_ready         ( pe38__std__lane27_strm1_ready      ),      
               .std__pe38__lane27_strm1_cntl          ( std__pe38__lane27_strm1_cntl       ),      
               .std__pe38__lane27_strm1_data          ( std__pe38__lane27_strm1_data       ),      
               .std__pe38__lane27_strm1_data_valid    ( std__pe38__lane27_strm1_data_valid ),      
               .std__pe38__lane27_strm1_data_mask     ( std__pe38__lane27_strm1_data_mask  ),      

               // PE 38, Lane 28                 
               .pe38__std__lane28_strm0_ready         ( pe38__std__lane28_strm0_ready      ),      
               .std__pe38__lane28_strm0_cntl          ( std__pe38__lane28_strm0_cntl       ),      
               .std__pe38__lane28_strm0_data          ( std__pe38__lane28_strm0_data       ),      
               .std__pe38__lane28_strm0_data_valid    ( std__pe38__lane28_strm0_data_valid ),      
               .std__pe38__lane28_strm0_data_mask     ( std__pe38__lane28_strm0_data_mask  ),      

               .pe38__std__lane28_strm1_ready         ( pe38__std__lane28_strm1_ready      ),      
               .std__pe38__lane28_strm1_cntl          ( std__pe38__lane28_strm1_cntl       ),      
               .std__pe38__lane28_strm1_data          ( std__pe38__lane28_strm1_data       ),      
               .std__pe38__lane28_strm1_data_valid    ( std__pe38__lane28_strm1_data_valid ),      
               .std__pe38__lane28_strm1_data_mask     ( std__pe38__lane28_strm1_data_mask  ),      

               // PE 38, Lane 29                 
               .pe38__std__lane29_strm0_ready         ( pe38__std__lane29_strm0_ready      ),      
               .std__pe38__lane29_strm0_cntl          ( std__pe38__lane29_strm0_cntl       ),      
               .std__pe38__lane29_strm0_data          ( std__pe38__lane29_strm0_data       ),      
               .std__pe38__lane29_strm0_data_valid    ( std__pe38__lane29_strm0_data_valid ),      
               .std__pe38__lane29_strm0_data_mask     ( std__pe38__lane29_strm0_data_mask  ),      

               .pe38__std__lane29_strm1_ready         ( pe38__std__lane29_strm1_ready      ),      
               .std__pe38__lane29_strm1_cntl          ( std__pe38__lane29_strm1_cntl       ),      
               .std__pe38__lane29_strm1_data          ( std__pe38__lane29_strm1_data       ),      
               .std__pe38__lane29_strm1_data_valid    ( std__pe38__lane29_strm1_data_valid ),      
               .std__pe38__lane29_strm1_data_mask     ( std__pe38__lane29_strm1_data_mask  ),      

               // PE 38, Lane 30                 
               .pe38__std__lane30_strm0_ready         ( pe38__std__lane30_strm0_ready      ),      
               .std__pe38__lane30_strm0_cntl          ( std__pe38__lane30_strm0_cntl       ),      
               .std__pe38__lane30_strm0_data          ( std__pe38__lane30_strm0_data       ),      
               .std__pe38__lane30_strm0_data_valid    ( std__pe38__lane30_strm0_data_valid ),      
               .std__pe38__lane30_strm0_data_mask     ( std__pe38__lane30_strm0_data_mask  ),      

               .pe38__std__lane30_strm1_ready         ( pe38__std__lane30_strm1_ready      ),      
               .std__pe38__lane30_strm1_cntl          ( std__pe38__lane30_strm1_cntl       ),      
               .std__pe38__lane30_strm1_data          ( std__pe38__lane30_strm1_data       ),      
               .std__pe38__lane30_strm1_data_valid    ( std__pe38__lane30_strm1_data_valid ),      
               .std__pe38__lane30_strm1_data_mask     ( std__pe38__lane30_strm1_data_mask  ),      

               // PE 38, Lane 31                 
               .pe38__std__lane31_strm0_ready         ( pe38__std__lane31_strm0_ready      ),      
               .std__pe38__lane31_strm0_cntl          ( std__pe38__lane31_strm0_cntl       ),      
               .std__pe38__lane31_strm0_data          ( std__pe38__lane31_strm0_data       ),      
               .std__pe38__lane31_strm0_data_valid    ( std__pe38__lane31_strm0_data_valid ),      
               .std__pe38__lane31_strm0_data_mask     ( std__pe38__lane31_strm0_data_mask  ),      

               .pe38__std__lane31_strm1_ready         ( pe38__std__lane31_strm1_ready      ),      
               .std__pe38__lane31_strm1_cntl          ( std__pe38__lane31_strm1_cntl       ),      
               .std__pe38__lane31_strm1_data          ( std__pe38__lane31_strm1_data       ),      
               .std__pe38__lane31_strm1_data_valid    ( std__pe38__lane31_strm1_data_valid ),      
               .std__pe38__lane31_strm1_data_mask     ( std__pe38__lane31_strm1_data_mask  ),      

               // PE 39, Lane 0                 
               .pe39__std__lane0_strm0_ready         ( pe39__std__lane0_strm0_ready      ),      
               .std__pe39__lane0_strm0_cntl          ( std__pe39__lane0_strm0_cntl       ),      
               .std__pe39__lane0_strm0_data          ( std__pe39__lane0_strm0_data       ),      
               .std__pe39__lane0_strm0_data_valid    ( std__pe39__lane0_strm0_data_valid ),      
               .std__pe39__lane0_strm0_data_mask     ( std__pe39__lane0_strm0_data_mask  ),      

               .pe39__std__lane0_strm1_ready         ( pe39__std__lane0_strm1_ready      ),      
               .std__pe39__lane0_strm1_cntl          ( std__pe39__lane0_strm1_cntl       ),      
               .std__pe39__lane0_strm1_data          ( std__pe39__lane0_strm1_data       ),      
               .std__pe39__lane0_strm1_data_valid    ( std__pe39__lane0_strm1_data_valid ),      
               .std__pe39__lane0_strm1_data_mask     ( std__pe39__lane0_strm1_data_mask  ),      

               // PE 39, Lane 1                 
               .pe39__std__lane1_strm0_ready         ( pe39__std__lane1_strm0_ready      ),      
               .std__pe39__lane1_strm0_cntl          ( std__pe39__lane1_strm0_cntl       ),      
               .std__pe39__lane1_strm0_data          ( std__pe39__lane1_strm0_data       ),      
               .std__pe39__lane1_strm0_data_valid    ( std__pe39__lane1_strm0_data_valid ),      
               .std__pe39__lane1_strm0_data_mask     ( std__pe39__lane1_strm0_data_mask  ),      

               .pe39__std__lane1_strm1_ready         ( pe39__std__lane1_strm1_ready      ),      
               .std__pe39__lane1_strm1_cntl          ( std__pe39__lane1_strm1_cntl       ),      
               .std__pe39__lane1_strm1_data          ( std__pe39__lane1_strm1_data       ),      
               .std__pe39__lane1_strm1_data_valid    ( std__pe39__lane1_strm1_data_valid ),      
               .std__pe39__lane1_strm1_data_mask     ( std__pe39__lane1_strm1_data_mask  ),      

               // PE 39, Lane 2                 
               .pe39__std__lane2_strm0_ready         ( pe39__std__lane2_strm0_ready      ),      
               .std__pe39__lane2_strm0_cntl          ( std__pe39__lane2_strm0_cntl       ),      
               .std__pe39__lane2_strm0_data          ( std__pe39__lane2_strm0_data       ),      
               .std__pe39__lane2_strm0_data_valid    ( std__pe39__lane2_strm0_data_valid ),      
               .std__pe39__lane2_strm0_data_mask     ( std__pe39__lane2_strm0_data_mask  ),      

               .pe39__std__lane2_strm1_ready         ( pe39__std__lane2_strm1_ready      ),      
               .std__pe39__lane2_strm1_cntl          ( std__pe39__lane2_strm1_cntl       ),      
               .std__pe39__lane2_strm1_data          ( std__pe39__lane2_strm1_data       ),      
               .std__pe39__lane2_strm1_data_valid    ( std__pe39__lane2_strm1_data_valid ),      
               .std__pe39__lane2_strm1_data_mask     ( std__pe39__lane2_strm1_data_mask  ),      

               // PE 39, Lane 3                 
               .pe39__std__lane3_strm0_ready         ( pe39__std__lane3_strm0_ready      ),      
               .std__pe39__lane3_strm0_cntl          ( std__pe39__lane3_strm0_cntl       ),      
               .std__pe39__lane3_strm0_data          ( std__pe39__lane3_strm0_data       ),      
               .std__pe39__lane3_strm0_data_valid    ( std__pe39__lane3_strm0_data_valid ),      
               .std__pe39__lane3_strm0_data_mask     ( std__pe39__lane3_strm0_data_mask  ),      

               .pe39__std__lane3_strm1_ready         ( pe39__std__lane3_strm1_ready      ),      
               .std__pe39__lane3_strm1_cntl          ( std__pe39__lane3_strm1_cntl       ),      
               .std__pe39__lane3_strm1_data          ( std__pe39__lane3_strm1_data       ),      
               .std__pe39__lane3_strm1_data_valid    ( std__pe39__lane3_strm1_data_valid ),      
               .std__pe39__lane3_strm1_data_mask     ( std__pe39__lane3_strm1_data_mask  ),      

               // PE 39, Lane 4                 
               .pe39__std__lane4_strm0_ready         ( pe39__std__lane4_strm0_ready      ),      
               .std__pe39__lane4_strm0_cntl          ( std__pe39__lane4_strm0_cntl       ),      
               .std__pe39__lane4_strm0_data          ( std__pe39__lane4_strm0_data       ),      
               .std__pe39__lane4_strm0_data_valid    ( std__pe39__lane4_strm0_data_valid ),      
               .std__pe39__lane4_strm0_data_mask     ( std__pe39__lane4_strm0_data_mask  ),      

               .pe39__std__lane4_strm1_ready         ( pe39__std__lane4_strm1_ready      ),      
               .std__pe39__lane4_strm1_cntl          ( std__pe39__lane4_strm1_cntl       ),      
               .std__pe39__lane4_strm1_data          ( std__pe39__lane4_strm1_data       ),      
               .std__pe39__lane4_strm1_data_valid    ( std__pe39__lane4_strm1_data_valid ),      
               .std__pe39__lane4_strm1_data_mask     ( std__pe39__lane4_strm1_data_mask  ),      

               // PE 39, Lane 5                 
               .pe39__std__lane5_strm0_ready         ( pe39__std__lane5_strm0_ready      ),      
               .std__pe39__lane5_strm0_cntl          ( std__pe39__lane5_strm0_cntl       ),      
               .std__pe39__lane5_strm0_data          ( std__pe39__lane5_strm0_data       ),      
               .std__pe39__lane5_strm0_data_valid    ( std__pe39__lane5_strm0_data_valid ),      
               .std__pe39__lane5_strm0_data_mask     ( std__pe39__lane5_strm0_data_mask  ),      

               .pe39__std__lane5_strm1_ready         ( pe39__std__lane5_strm1_ready      ),      
               .std__pe39__lane5_strm1_cntl          ( std__pe39__lane5_strm1_cntl       ),      
               .std__pe39__lane5_strm1_data          ( std__pe39__lane5_strm1_data       ),      
               .std__pe39__lane5_strm1_data_valid    ( std__pe39__lane5_strm1_data_valid ),      
               .std__pe39__lane5_strm1_data_mask     ( std__pe39__lane5_strm1_data_mask  ),      

               // PE 39, Lane 6                 
               .pe39__std__lane6_strm0_ready         ( pe39__std__lane6_strm0_ready      ),      
               .std__pe39__lane6_strm0_cntl          ( std__pe39__lane6_strm0_cntl       ),      
               .std__pe39__lane6_strm0_data          ( std__pe39__lane6_strm0_data       ),      
               .std__pe39__lane6_strm0_data_valid    ( std__pe39__lane6_strm0_data_valid ),      
               .std__pe39__lane6_strm0_data_mask     ( std__pe39__lane6_strm0_data_mask  ),      

               .pe39__std__lane6_strm1_ready         ( pe39__std__lane6_strm1_ready      ),      
               .std__pe39__lane6_strm1_cntl          ( std__pe39__lane6_strm1_cntl       ),      
               .std__pe39__lane6_strm1_data          ( std__pe39__lane6_strm1_data       ),      
               .std__pe39__lane6_strm1_data_valid    ( std__pe39__lane6_strm1_data_valid ),      
               .std__pe39__lane6_strm1_data_mask     ( std__pe39__lane6_strm1_data_mask  ),      

               // PE 39, Lane 7                 
               .pe39__std__lane7_strm0_ready         ( pe39__std__lane7_strm0_ready      ),      
               .std__pe39__lane7_strm0_cntl          ( std__pe39__lane7_strm0_cntl       ),      
               .std__pe39__lane7_strm0_data          ( std__pe39__lane7_strm0_data       ),      
               .std__pe39__lane7_strm0_data_valid    ( std__pe39__lane7_strm0_data_valid ),      
               .std__pe39__lane7_strm0_data_mask     ( std__pe39__lane7_strm0_data_mask  ),      

               .pe39__std__lane7_strm1_ready         ( pe39__std__lane7_strm1_ready      ),      
               .std__pe39__lane7_strm1_cntl          ( std__pe39__lane7_strm1_cntl       ),      
               .std__pe39__lane7_strm1_data          ( std__pe39__lane7_strm1_data       ),      
               .std__pe39__lane7_strm1_data_valid    ( std__pe39__lane7_strm1_data_valid ),      
               .std__pe39__lane7_strm1_data_mask     ( std__pe39__lane7_strm1_data_mask  ),      

               // PE 39, Lane 8                 
               .pe39__std__lane8_strm0_ready         ( pe39__std__lane8_strm0_ready      ),      
               .std__pe39__lane8_strm0_cntl          ( std__pe39__lane8_strm0_cntl       ),      
               .std__pe39__lane8_strm0_data          ( std__pe39__lane8_strm0_data       ),      
               .std__pe39__lane8_strm0_data_valid    ( std__pe39__lane8_strm0_data_valid ),      
               .std__pe39__lane8_strm0_data_mask     ( std__pe39__lane8_strm0_data_mask  ),      

               .pe39__std__lane8_strm1_ready         ( pe39__std__lane8_strm1_ready      ),      
               .std__pe39__lane8_strm1_cntl          ( std__pe39__lane8_strm1_cntl       ),      
               .std__pe39__lane8_strm1_data          ( std__pe39__lane8_strm1_data       ),      
               .std__pe39__lane8_strm1_data_valid    ( std__pe39__lane8_strm1_data_valid ),      
               .std__pe39__lane8_strm1_data_mask     ( std__pe39__lane8_strm1_data_mask  ),      

               // PE 39, Lane 9                 
               .pe39__std__lane9_strm0_ready         ( pe39__std__lane9_strm0_ready      ),      
               .std__pe39__lane9_strm0_cntl          ( std__pe39__lane9_strm0_cntl       ),      
               .std__pe39__lane9_strm0_data          ( std__pe39__lane9_strm0_data       ),      
               .std__pe39__lane9_strm0_data_valid    ( std__pe39__lane9_strm0_data_valid ),      
               .std__pe39__lane9_strm0_data_mask     ( std__pe39__lane9_strm0_data_mask  ),      

               .pe39__std__lane9_strm1_ready         ( pe39__std__lane9_strm1_ready      ),      
               .std__pe39__lane9_strm1_cntl          ( std__pe39__lane9_strm1_cntl       ),      
               .std__pe39__lane9_strm1_data          ( std__pe39__lane9_strm1_data       ),      
               .std__pe39__lane9_strm1_data_valid    ( std__pe39__lane9_strm1_data_valid ),      
               .std__pe39__lane9_strm1_data_mask     ( std__pe39__lane9_strm1_data_mask  ),      

               // PE 39, Lane 10                 
               .pe39__std__lane10_strm0_ready         ( pe39__std__lane10_strm0_ready      ),      
               .std__pe39__lane10_strm0_cntl          ( std__pe39__lane10_strm0_cntl       ),      
               .std__pe39__lane10_strm0_data          ( std__pe39__lane10_strm0_data       ),      
               .std__pe39__lane10_strm0_data_valid    ( std__pe39__lane10_strm0_data_valid ),      
               .std__pe39__lane10_strm0_data_mask     ( std__pe39__lane10_strm0_data_mask  ),      

               .pe39__std__lane10_strm1_ready         ( pe39__std__lane10_strm1_ready      ),      
               .std__pe39__lane10_strm1_cntl          ( std__pe39__lane10_strm1_cntl       ),      
               .std__pe39__lane10_strm1_data          ( std__pe39__lane10_strm1_data       ),      
               .std__pe39__lane10_strm1_data_valid    ( std__pe39__lane10_strm1_data_valid ),      
               .std__pe39__lane10_strm1_data_mask     ( std__pe39__lane10_strm1_data_mask  ),      

               // PE 39, Lane 11                 
               .pe39__std__lane11_strm0_ready         ( pe39__std__lane11_strm0_ready      ),      
               .std__pe39__lane11_strm0_cntl          ( std__pe39__lane11_strm0_cntl       ),      
               .std__pe39__lane11_strm0_data          ( std__pe39__lane11_strm0_data       ),      
               .std__pe39__lane11_strm0_data_valid    ( std__pe39__lane11_strm0_data_valid ),      
               .std__pe39__lane11_strm0_data_mask     ( std__pe39__lane11_strm0_data_mask  ),      

               .pe39__std__lane11_strm1_ready         ( pe39__std__lane11_strm1_ready      ),      
               .std__pe39__lane11_strm1_cntl          ( std__pe39__lane11_strm1_cntl       ),      
               .std__pe39__lane11_strm1_data          ( std__pe39__lane11_strm1_data       ),      
               .std__pe39__lane11_strm1_data_valid    ( std__pe39__lane11_strm1_data_valid ),      
               .std__pe39__lane11_strm1_data_mask     ( std__pe39__lane11_strm1_data_mask  ),      

               // PE 39, Lane 12                 
               .pe39__std__lane12_strm0_ready         ( pe39__std__lane12_strm0_ready      ),      
               .std__pe39__lane12_strm0_cntl          ( std__pe39__lane12_strm0_cntl       ),      
               .std__pe39__lane12_strm0_data          ( std__pe39__lane12_strm0_data       ),      
               .std__pe39__lane12_strm0_data_valid    ( std__pe39__lane12_strm0_data_valid ),      
               .std__pe39__lane12_strm0_data_mask     ( std__pe39__lane12_strm0_data_mask  ),      

               .pe39__std__lane12_strm1_ready         ( pe39__std__lane12_strm1_ready      ),      
               .std__pe39__lane12_strm1_cntl          ( std__pe39__lane12_strm1_cntl       ),      
               .std__pe39__lane12_strm1_data          ( std__pe39__lane12_strm1_data       ),      
               .std__pe39__lane12_strm1_data_valid    ( std__pe39__lane12_strm1_data_valid ),      
               .std__pe39__lane12_strm1_data_mask     ( std__pe39__lane12_strm1_data_mask  ),      

               // PE 39, Lane 13                 
               .pe39__std__lane13_strm0_ready         ( pe39__std__lane13_strm0_ready      ),      
               .std__pe39__lane13_strm0_cntl          ( std__pe39__lane13_strm0_cntl       ),      
               .std__pe39__lane13_strm0_data          ( std__pe39__lane13_strm0_data       ),      
               .std__pe39__lane13_strm0_data_valid    ( std__pe39__lane13_strm0_data_valid ),      
               .std__pe39__lane13_strm0_data_mask     ( std__pe39__lane13_strm0_data_mask  ),      

               .pe39__std__lane13_strm1_ready         ( pe39__std__lane13_strm1_ready      ),      
               .std__pe39__lane13_strm1_cntl          ( std__pe39__lane13_strm1_cntl       ),      
               .std__pe39__lane13_strm1_data          ( std__pe39__lane13_strm1_data       ),      
               .std__pe39__lane13_strm1_data_valid    ( std__pe39__lane13_strm1_data_valid ),      
               .std__pe39__lane13_strm1_data_mask     ( std__pe39__lane13_strm1_data_mask  ),      

               // PE 39, Lane 14                 
               .pe39__std__lane14_strm0_ready         ( pe39__std__lane14_strm0_ready      ),      
               .std__pe39__lane14_strm0_cntl          ( std__pe39__lane14_strm0_cntl       ),      
               .std__pe39__lane14_strm0_data          ( std__pe39__lane14_strm0_data       ),      
               .std__pe39__lane14_strm0_data_valid    ( std__pe39__lane14_strm0_data_valid ),      
               .std__pe39__lane14_strm0_data_mask     ( std__pe39__lane14_strm0_data_mask  ),      

               .pe39__std__lane14_strm1_ready         ( pe39__std__lane14_strm1_ready      ),      
               .std__pe39__lane14_strm1_cntl          ( std__pe39__lane14_strm1_cntl       ),      
               .std__pe39__lane14_strm1_data          ( std__pe39__lane14_strm1_data       ),      
               .std__pe39__lane14_strm1_data_valid    ( std__pe39__lane14_strm1_data_valid ),      
               .std__pe39__lane14_strm1_data_mask     ( std__pe39__lane14_strm1_data_mask  ),      

               // PE 39, Lane 15                 
               .pe39__std__lane15_strm0_ready         ( pe39__std__lane15_strm0_ready      ),      
               .std__pe39__lane15_strm0_cntl          ( std__pe39__lane15_strm0_cntl       ),      
               .std__pe39__lane15_strm0_data          ( std__pe39__lane15_strm0_data       ),      
               .std__pe39__lane15_strm0_data_valid    ( std__pe39__lane15_strm0_data_valid ),      
               .std__pe39__lane15_strm0_data_mask     ( std__pe39__lane15_strm0_data_mask  ),      

               .pe39__std__lane15_strm1_ready         ( pe39__std__lane15_strm1_ready      ),      
               .std__pe39__lane15_strm1_cntl          ( std__pe39__lane15_strm1_cntl       ),      
               .std__pe39__lane15_strm1_data          ( std__pe39__lane15_strm1_data       ),      
               .std__pe39__lane15_strm1_data_valid    ( std__pe39__lane15_strm1_data_valid ),      
               .std__pe39__lane15_strm1_data_mask     ( std__pe39__lane15_strm1_data_mask  ),      

               // PE 39, Lane 16                 
               .pe39__std__lane16_strm0_ready         ( pe39__std__lane16_strm0_ready      ),      
               .std__pe39__lane16_strm0_cntl          ( std__pe39__lane16_strm0_cntl       ),      
               .std__pe39__lane16_strm0_data          ( std__pe39__lane16_strm0_data       ),      
               .std__pe39__lane16_strm0_data_valid    ( std__pe39__lane16_strm0_data_valid ),      
               .std__pe39__lane16_strm0_data_mask     ( std__pe39__lane16_strm0_data_mask  ),      

               .pe39__std__lane16_strm1_ready         ( pe39__std__lane16_strm1_ready      ),      
               .std__pe39__lane16_strm1_cntl          ( std__pe39__lane16_strm1_cntl       ),      
               .std__pe39__lane16_strm1_data          ( std__pe39__lane16_strm1_data       ),      
               .std__pe39__lane16_strm1_data_valid    ( std__pe39__lane16_strm1_data_valid ),      
               .std__pe39__lane16_strm1_data_mask     ( std__pe39__lane16_strm1_data_mask  ),      

               // PE 39, Lane 17                 
               .pe39__std__lane17_strm0_ready         ( pe39__std__lane17_strm0_ready      ),      
               .std__pe39__lane17_strm0_cntl          ( std__pe39__lane17_strm0_cntl       ),      
               .std__pe39__lane17_strm0_data          ( std__pe39__lane17_strm0_data       ),      
               .std__pe39__lane17_strm0_data_valid    ( std__pe39__lane17_strm0_data_valid ),      
               .std__pe39__lane17_strm0_data_mask     ( std__pe39__lane17_strm0_data_mask  ),      

               .pe39__std__lane17_strm1_ready         ( pe39__std__lane17_strm1_ready      ),      
               .std__pe39__lane17_strm1_cntl          ( std__pe39__lane17_strm1_cntl       ),      
               .std__pe39__lane17_strm1_data          ( std__pe39__lane17_strm1_data       ),      
               .std__pe39__lane17_strm1_data_valid    ( std__pe39__lane17_strm1_data_valid ),      
               .std__pe39__lane17_strm1_data_mask     ( std__pe39__lane17_strm1_data_mask  ),      

               // PE 39, Lane 18                 
               .pe39__std__lane18_strm0_ready         ( pe39__std__lane18_strm0_ready      ),      
               .std__pe39__lane18_strm0_cntl          ( std__pe39__lane18_strm0_cntl       ),      
               .std__pe39__lane18_strm0_data          ( std__pe39__lane18_strm0_data       ),      
               .std__pe39__lane18_strm0_data_valid    ( std__pe39__lane18_strm0_data_valid ),      
               .std__pe39__lane18_strm0_data_mask     ( std__pe39__lane18_strm0_data_mask  ),      

               .pe39__std__lane18_strm1_ready         ( pe39__std__lane18_strm1_ready      ),      
               .std__pe39__lane18_strm1_cntl          ( std__pe39__lane18_strm1_cntl       ),      
               .std__pe39__lane18_strm1_data          ( std__pe39__lane18_strm1_data       ),      
               .std__pe39__lane18_strm1_data_valid    ( std__pe39__lane18_strm1_data_valid ),      
               .std__pe39__lane18_strm1_data_mask     ( std__pe39__lane18_strm1_data_mask  ),      

               // PE 39, Lane 19                 
               .pe39__std__lane19_strm0_ready         ( pe39__std__lane19_strm0_ready      ),      
               .std__pe39__lane19_strm0_cntl          ( std__pe39__lane19_strm0_cntl       ),      
               .std__pe39__lane19_strm0_data          ( std__pe39__lane19_strm0_data       ),      
               .std__pe39__lane19_strm0_data_valid    ( std__pe39__lane19_strm0_data_valid ),      
               .std__pe39__lane19_strm0_data_mask     ( std__pe39__lane19_strm0_data_mask  ),      

               .pe39__std__lane19_strm1_ready         ( pe39__std__lane19_strm1_ready      ),      
               .std__pe39__lane19_strm1_cntl          ( std__pe39__lane19_strm1_cntl       ),      
               .std__pe39__lane19_strm1_data          ( std__pe39__lane19_strm1_data       ),      
               .std__pe39__lane19_strm1_data_valid    ( std__pe39__lane19_strm1_data_valid ),      
               .std__pe39__lane19_strm1_data_mask     ( std__pe39__lane19_strm1_data_mask  ),      

               // PE 39, Lane 20                 
               .pe39__std__lane20_strm0_ready         ( pe39__std__lane20_strm0_ready      ),      
               .std__pe39__lane20_strm0_cntl          ( std__pe39__lane20_strm0_cntl       ),      
               .std__pe39__lane20_strm0_data          ( std__pe39__lane20_strm0_data       ),      
               .std__pe39__lane20_strm0_data_valid    ( std__pe39__lane20_strm0_data_valid ),      
               .std__pe39__lane20_strm0_data_mask     ( std__pe39__lane20_strm0_data_mask  ),      

               .pe39__std__lane20_strm1_ready         ( pe39__std__lane20_strm1_ready      ),      
               .std__pe39__lane20_strm1_cntl          ( std__pe39__lane20_strm1_cntl       ),      
               .std__pe39__lane20_strm1_data          ( std__pe39__lane20_strm1_data       ),      
               .std__pe39__lane20_strm1_data_valid    ( std__pe39__lane20_strm1_data_valid ),      
               .std__pe39__lane20_strm1_data_mask     ( std__pe39__lane20_strm1_data_mask  ),      

               // PE 39, Lane 21                 
               .pe39__std__lane21_strm0_ready         ( pe39__std__lane21_strm0_ready      ),      
               .std__pe39__lane21_strm0_cntl          ( std__pe39__lane21_strm0_cntl       ),      
               .std__pe39__lane21_strm0_data          ( std__pe39__lane21_strm0_data       ),      
               .std__pe39__lane21_strm0_data_valid    ( std__pe39__lane21_strm0_data_valid ),      
               .std__pe39__lane21_strm0_data_mask     ( std__pe39__lane21_strm0_data_mask  ),      

               .pe39__std__lane21_strm1_ready         ( pe39__std__lane21_strm1_ready      ),      
               .std__pe39__lane21_strm1_cntl          ( std__pe39__lane21_strm1_cntl       ),      
               .std__pe39__lane21_strm1_data          ( std__pe39__lane21_strm1_data       ),      
               .std__pe39__lane21_strm1_data_valid    ( std__pe39__lane21_strm1_data_valid ),      
               .std__pe39__lane21_strm1_data_mask     ( std__pe39__lane21_strm1_data_mask  ),      

               // PE 39, Lane 22                 
               .pe39__std__lane22_strm0_ready         ( pe39__std__lane22_strm0_ready      ),      
               .std__pe39__lane22_strm0_cntl          ( std__pe39__lane22_strm0_cntl       ),      
               .std__pe39__lane22_strm0_data          ( std__pe39__lane22_strm0_data       ),      
               .std__pe39__lane22_strm0_data_valid    ( std__pe39__lane22_strm0_data_valid ),      
               .std__pe39__lane22_strm0_data_mask     ( std__pe39__lane22_strm0_data_mask  ),      

               .pe39__std__lane22_strm1_ready         ( pe39__std__lane22_strm1_ready      ),      
               .std__pe39__lane22_strm1_cntl          ( std__pe39__lane22_strm1_cntl       ),      
               .std__pe39__lane22_strm1_data          ( std__pe39__lane22_strm1_data       ),      
               .std__pe39__lane22_strm1_data_valid    ( std__pe39__lane22_strm1_data_valid ),      
               .std__pe39__lane22_strm1_data_mask     ( std__pe39__lane22_strm1_data_mask  ),      

               // PE 39, Lane 23                 
               .pe39__std__lane23_strm0_ready         ( pe39__std__lane23_strm0_ready      ),      
               .std__pe39__lane23_strm0_cntl          ( std__pe39__lane23_strm0_cntl       ),      
               .std__pe39__lane23_strm0_data          ( std__pe39__lane23_strm0_data       ),      
               .std__pe39__lane23_strm0_data_valid    ( std__pe39__lane23_strm0_data_valid ),      
               .std__pe39__lane23_strm0_data_mask     ( std__pe39__lane23_strm0_data_mask  ),      

               .pe39__std__lane23_strm1_ready         ( pe39__std__lane23_strm1_ready      ),      
               .std__pe39__lane23_strm1_cntl          ( std__pe39__lane23_strm1_cntl       ),      
               .std__pe39__lane23_strm1_data          ( std__pe39__lane23_strm1_data       ),      
               .std__pe39__lane23_strm1_data_valid    ( std__pe39__lane23_strm1_data_valid ),      
               .std__pe39__lane23_strm1_data_mask     ( std__pe39__lane23_strm1_data_mask  ),      

               // PE 39, Lane 24                 
               .pe39__std__lane24_strm0_ready         ( pe39__std__lane24_strm0_ready      ),      
               .std__pe39__lane24_strm0_cntl          ( std__pe39__lane24_strm0_cntl       ),      
               .std__pe39__lane24_strm0_data          ( std__pe39__lane24_strm0_data       ),      
               .std__pe39__lane24_strm0_data_valid    ( std__pe39__lane24_strm0_data_valid ),      
               .std__pe39__lane24_strm0_data_mask     ( std__pe39__lane24_strm0_data_mask  ),      

               .pe39__std__lane24_strm1_ready         ( pe39__std__lane24_strm1_ready      ),      
               .std__pe39__lane24_strm1_cntl          ( std__pe39__lane24_strm1_cntl       ),      
               .std__pe39__lane24_strm1_data          ( std__pe39__lane24_strm1_data       ),      
               .std__pe39__lane24_strm1_data_valid    ( std__pe39__lane24_strm1_data_valid ),      
               .std__pe39__lane24_strm1_data_mask     ( std__pe39__lane24_strm1_data_mask  ),      

               // PE 39, Lane 25                 
               .pe39__std__lane25_strm0_ready         ( pe39__std__lane25_strm0_ready      ),      
               .std__pe39__lane25_strm0_cntl          ( std__pe39__lane25_strm0_cntl       ),      
               .std__pe39__lane25_strm0_data          ( std__pe39__lane25_strm0_data       ),      
               .std__pe39__lane25_strm0_data_valid    ( std__pe39__lane25_strm0_data_valid ),      
               .std__pe39__lane25_strm0_data_mask     ( std__pe39__lane25_strm0_data_mask  ),      

               .pe39__std__lane25_strm1_ready         ( pe39__std__lane25_strm1_ready      ),      
               .std__pe39__lane25_strm1_cntl          ( std__pe39__lane25_strm1_cntl       ),      
               .std__pe39__lane25_strm1_data          ( std__pe39__lane25_strm1_data       ),      
               .std__pe39__lane25_strm1_data_valid    ( std__pe39__lane25_strm1_data_valid ),      
               .std__pe39__lane25_strm1_data_mask     ( std__pe39__lane25_strm1_data_mask  ),      

               // PE 39, Lane 26                 
               .pe39__std__lane26_strm0_ready         ( pe39__std__lane26_strm0_ready      ),      
               .std__pe39__lane26_strm0_cntl          ( std__pe39__lane26_strm0_cntl       ),      
               .std__pe39__lane26_strm0_data          ( std__pe39__lane26_strm0_data       ),      
               .std__pe39__lane26_strm0_data_valid    ( std__pe39__lane26_strm0_data_valid ),      
               .std__pe39__lane26_strm0_data_mask     ( std__pe39__lane26_strm0_data_mask  ),      

               .pe39__std__lane26_strm1_ready         ( pe39__std__lane26_strm1_ready      ),      
               .std__pe39__lane26_strm1_cntl          ( std__pe39__lane26_strm1_cntl       ),      
               .std__pe39__lane26_strm1_data          ( std__pe39__lane26_strm1_data       ),      
               .std__pe39__lane26_strm1_data_valid    ( std__pe39__lane26_strm1_data_valid ),      
               .std__pe39__lane26_strm1_data_mask     ( std__pe39__lane26_strm1_data_mask  ),      

               // PE 39, Lane 27                 
               .pe39__std__lane27_strm0_ready         ( pe39__std__lane27_strm0_ready      ),      
               .std__pe39__lane27_strm0_cntl          ( std__pe39__lane27_strm0_cntl       ),      
               .std__pe39__lane27_strm0_data          ( std__pe39__lane27_strm0_data       ),      
               .std__pe39__lane27_strm0_data_valid    ( std__pe39__lane27_strm0_data_valid ),      
               .std__pe39__lane27_strm0_data_mask     ( std__pe39__lane27_strm0_data_mask  ),      

               .pe39__std__lane27_strm1_ready         ( pe39__std__lane27_strm1_ready      ),      
               .std__pe39__lane27_strm1_cntl          ( std__pe39__lane27_strm1_cntl       ),      
               .std__pe39__lane27_strm1_data          ( std__pe39__lane27_strm1_data       ),      
               .std__pe39__lane27_strm1_data_valid    ( std__pe39__lane27_strm1_data_valid ),      
               .std__pe39__lane27_strm1_data_mask     ( std__pe39__lane27_strm1_data_mask  ),      

               // PE 39, Lane 28                 
               .pe39__std__lane28_strm0_ready         ( pe39__std__lane28_strm0_ready      ),      
               .std__pe39__lane28_strm0_cntl          ( std__pe39__lane28_strm0_cntl       ),      
               .std__pe39__lane28_strm0_data          ( std__pe39__lane28_strm0_data       ),      
               .std__pe39__lane28_strm0_data_valid    ( std__pe39__lane28_strm0_data_valid ),      
               .std__pe39__lane28_strm0_data_mask     ( std__pe39__lane28_strm0_data_mask  ),      

               .pe39__std__lane28_strm1_ready         ( pe39__std__lane28_strm1_ready      ),      
               .std__pe39__lane28_strm1_cntl          ( std__pe39__lane28_strm1_cntl       ),      
               .std__pe39__lane28_strm1_data          ( std__pe39__lane28_strm1_data       ),      
               .std__pe39__lane28_strm1_data_valid    ( std__pe39__lane28_strm1_data_valid ),      
               .std__pe39__lane28_strm1_data_mask     ( std__pe39__lane28_strm1_data_mask  ),      

               // PE 39, Lane 29                 
               .pe39__std__lane29_strm0_ready         ( pe39__std__lane29_strm0_ready      ),      
               .std__pe39__lane29_strm0_cntl          ( std__pe39__lane29_strm0_cntl       ),      
               .std__pe39__lane29_strm0_data          ( std__pe39__lane29_strm0_data       ),      
               .std__pe39__lane29_strm0_data_valid    ( std__pe39__lane29_strm0_data_valid ),      
               .std__pe39__lane29_strm0_data_mask     ( std__pe39__lane29_strm0_data_mask  ),      

               .pe39__std__lane29_strm1_ready         ( pe39__std__lane29_strm1_ready      ),      
               .std__pe39__lane29_strm1_cntl          ( std__pe39__lane29_strm1_cntl       ),      
               .std__pe39__lane29_strm1_data          ( std__pe39__lane29_strm1_data       ),      
               .std__pe39__lane29_strm1_data_valid    ( std__pe39__lane29_strm1_data_valid ),      
               .std__pe39__lane29_strm1_data_mask     ( std__pe39__lane29_strm1_data_mask  ),      

               // PE 39, Lane 30                 
               .pe39__std__lane30_strm0_ready         ( pe39__std__lane30_strm0_ready      ),      
               .std__pe39__lane30_strm0_cntl          ( std__pe39__lane30_strm0_cntl       ),      
               .std__pe39__lane30_strm0_data          ( std__pe39__lane30_strm0_data       ),      
               .std__pe39__lane30_strm0_data_valid    ( std__pe39__lane30_strm0_data_valid ),      
               .std__pe39__lane30_strm0_data_mask     ( std__pe39__lane30_strm0_data_mask  ),      

               .pe39__std__lane30_strm1_ready         ( pe39__std__lane30_strm1_ready      ),      
               .std__pe39__lane30_strm1_cntl          ( std__pe39__lane30_strm1_cntl       ),      
               .std__pe39__lane30_strm1_data          ( std__pe39__lane30_strm1_data       ),      
               .std__pe39__lane30_strm1_data_valid    ( std__pe39__lane30_strm1_data_valid ),      
               .std__pe39__lane30_strm1_data_mask     ( std__pe39__lane30_strm1_data_mask  ),      

               // PE 39, Lane 31                 
               .pe39__std__lane31_strm0_ready         ( pe39__std__lane31_strm0_ready      ),      
               .std__pe39__lane31_strm0_cntl          ( std__pe39__lane31_strm0_cntl       ),      
               .std__pe39__lane31_strm0_data          ( std__pe39__lane31_strm0_data       ),      
               .std__pe39__lane31_strm0_data_valid    ( std__pe39__lane31_strm0_data_valid ),      
               .std__pe39__lane31_strm0_data_mask     ( std__pe39__lane31_strm0_data_mask  ),      

               .pe39__std__lane31_strm1_ready         ( pe39__std__lane31_strm1_ready      ),      
               .std__pe39__lane31_strm1_cntl          ( std__pe39__lane31_strm1_cntl       ),      
               .std__pe39__lane31_strm1_data          ( std__pe39__lane31_strm1_data       ),      
               .std__pe39__lane31_strm1_data_valid    ( std__pe39__lane31_strm1_data_valid ),      
               .std__pe39__lane31_strm1_data_mask     ( std__pe39__lane31_strm1_data_mask  ),      

               // PE 40, Lane 0                 
               .pe40__std__lane0_strm0_ready         ( pe40__std__lane0_strm0_ready      ),      
               .std__pe40__lane0_strm0_cntl          ( std__pe40__lane0_strm0_cntl       ),      
               .std__pe40__lane0_strm0_data          ( std__pe40__lane0_strm0_data       ),      
               .std__pe40__lane0_strm0_data_valid    ( std__pe40__lane0_strm0_data_valid ),      
               .std__pe40__lane0_strm0_data_mask     ( std__pe40__lane0_strm0_data_mask  ),      

               .pe40__std__lane0_strm1_ready         ( pe40__std__lane0_strm1_ready      ),      
               .std__pe40__lane0_strm1_cntl          ( std__pe40__lane0_strm1_cntl       ),      
               .std__pe40__lane0_strm1_data          ( std__pe40__lane0_strm1_data       ),      
               .std__pe40__lane0_strm1_data_valid    ( std__pe40__lane0_strm1_data_valid ),      
               .std__pe40__lane0_strm1_data_mask     ( std__pe40__lane0_strm1_data_mask  ),      

               // PE 40, Lane 1                 
               .pe40__std__lane1_strm0_ready         ( pe40__std__lane1_strm0_ready      ),      
               .std__pe40__lane1_strm0_cntl          ( std__pe40__lane1_strm0_cntl       ),      
               .std__pe40__lane1_strm0_data          ( std__pe40__lane1_strm0_data       ),      
               .std__pe40__lane1_strm0_data_valid    ( std__pe40__lane1_strm0_data_valid ),      
               .std__pe40__lane1_strm0_data_mask     ( std__pe40__lane1_strm0_data_mask  ),      

               .pe40__std__lane1_strm1_ready         ( pe40__std__lane1_strm1_ready      ),      
               .std__pe40__lane1_strm1_cntl          ( std__pe40__lane1_strm1_cntl       ),      
               .std__pe40__lane1_strm1_data          ( std__pe40__lane1_strm1_data       ),      
               .std__pe40__lane1_strm1_data_valid    ( std__pe40__lane1_strm1_data_valid ),      
               .std__pe40__lane1_strm1_data_mask     ( std__pe40__lane1_strm1_data_mask  ),      

               // PE 40, Lane 2                 
               .pe40__std__lane2_strm0_ready         ( pe40__std__lane2_strm0_ready      ),      
               .std__pe40__lane2_strm0_cntl          ( std__pe40__lane2_strm0_cntl       ),      
               .std__pe40__lane2_strm0_data          ( std__pe40__lane2_strm0_data       ),      
               .std__pe40__lane2_strm0_data_valid    ( std__pe40__lane2_strm0_data_valid ),      
               .std__pe40__lane2_strm0_data_mask     ( std__pe40__lane2_strm0_data_mask  ),      

               .pe40__std__lane2_strm1_ready         ( pe40__std__lane2_strm1_ready      ),      
               .std__pe40__lane2_strm1_cntl          ( std__pe40__lane2_strm1_cntl       ),      
               .std__pe40__lane2_strm1_data          ( std__pe40__lane2_strm1_data       ),      
               .std__pe40__lane2_strm1_data_valid    ( std__pe40__lane2_strm1_data_valid ),      
               .std__pe40__lane2_strm1_data_mask     ( std__pe40__lane2_strm1_data_mask  ),      

               // PE 40, Lane 3                 
               .pe40__std__lane3_strm0_ready         ( pe40__std__lane3_strm0_ready      ),      
               .std__pe40__lane3_strm0_cntl          ( std__pe40__lane3_strm0_cntl       ),      
               .std__pe40__lane3_strm0_data          ( std__pe40__lane3_strm0_data       ),      
               .std__pe40__lane3_strm0_data_valid    ( std__pe40__lane3_strm0_data_valid ),      
               .std__pe40__lane3_strm0_data_mask     ( std__pe40__lane3_strm0_data_mask  ),      

               .pe40__std__lane3_strm1_ready         ( pe40__std__lane3_strm1_ready      ),      
               .std__pe40__lane3_strm1_cntl          ( std__pe40__lane3_strm1_cntl       ),      
               .std__pe40__lane3_strm1_data          ( std__pe40__lane3_strm1_data       ),      
               .std__pe40__lane3_strm1_data_valid    ( std__pe40__lane3_strm1_data_valid ),      
               .std__pe40__lane3_strm1_data_mask     ( std__pe40__lane3_strm1_data_mask  ),      

               // PE 40, Lane 4                 
               .pe40__std__lane4_strm0_ready         ( pe40__std__lane4_strm0_ready      ),      
               .std__pe40__lane4_strm0_cntl          ( std__pe40__lane4_strm0_cntl       ),      
               .std__pe40__lane4_strm0_data          ( std__pe40__lane4_strm0_data       ),      
               .std__pe40__lane4_strm0_data_valid    ( std__pe40__lane4_strm0_data_valid ),      
               .std__pe40__lane4_strm0_data_mask     ( std__pe40__lane4_strm0_data_mask  ),      

               .pe40__std__lane4_strm1_ready         ( pe40__std__lane4_strm1_ready      ),      
               .std__pe40__lane4_strm1_cntl          ( std__pe40__lane4_strm1_cntl       ),      
               .std__pe40__lane4_strm1_data          ( std__pe40__lane4_strm1_data       ),      
               .std__pe40__lane4_strm1_data_valid    ( std__pe40__lane4_strm1_data_valid ),      
               .std__pe40__lane4_strm1_data_mask     ( std__pe40__lane4_strm1_data_mask  ),      

               // PE 40, Lane 5                 
               .pe40__std__lane5_strm0_ready         ( pe40__std__lane5_strm0_ready      ),      
               .std__pe40__lane5_strm0_cntl          ( std__pe40__lane5_strm0_cntl       ),      
               .std__pe40__lane5_strm0_data          ( std__pe40__lane5_strm0_data       ),      
               .std__pe40__lane5_strm0_data_valid    ( std__pe40__lane5_strm0_data_valid ),      
               .std__pe40__lane5_strm0_data_mask     ( std__pe40__lane5_strm0_data_mask  ),      

               .pe40__std__lane5_strm1_ready         ( pe40__std__lane5_strm1_ready      ),      
               .std__pe40__lane5_strm1_cntl          ( std__pe40__lane5_strm1_cntl       ),      
               .std__pe40__lane5_strm1_data          ( std__pe40__lane5_strm1_data       ),      
               .std__pe40__lane5_strm1_data_valid    ( std__pe40__lane5_strm1_data_valid ),      
               .std__pe40__lane5_strm1_data_mask     ( std__pe40__lane5_strm1_data_mask  ),      

               // PE 40, Lane 6                 
               .pe40__std__lane6_strm0_ready         ( pe40__std__lane6_strm0_ready      ),      
               .std__pe40__lane6_strm0_cntl          ( std__pe40__lane6_strm0_cntl       ),      
               .std__pe40__lane6_strm0_data          ( std__pe40__lane6_strm0_data       ),      
               .std__pe40__lane6_strm0_data_valid    ( std__pe40__lane6_strm0_data_valid ),      
               .std__pe40__lane6_strm0_data_mask     ( std__pe40__lane6_strm0_data_mask  ),      

               .pe40__std__lane6_strm1_ready         ( pe40__std__lane6_strm1_ready      ),      
               .std__pe40__lane6_strm1_cntl          ( std__pe40__lane6_strm1_cntl       ),      
               .std__pe40__lane6_strm1_data          ( std__pe40__lane6_strm1_data       ),      
               .std__pe40__lane6_strm1_data_valid    ( std__pe40__lane6_strm1_data_valid ),      
               .std__pe40__lane6_strm1_data_mask     ( std__pe40__lane6_strm1_data_mask  ),      

               // PE 40, Lane 7                 
               .pe40__std__lane7_strm0_ready         ( pe40__std__lane7_strm0_ready      ),      
               .std__pe40__lane7_strm0_cntl          ( std__pe40__lane7_strm0_cntl       ),      
               .std__pe40__lane7_strm0_data          ( std__pe40__lane7_strm0_data       ),      
               .std__pe40__lane7_strm0_data_valid    ( std__pe40__lane7_strm0_data_valid ),      
               .std__pe40__lane7_strm0_data_mask     ( std__pe40__lane7_strm0_data_mask  ),      

               .pe40__std__lane7_strm1_ready         ( pe40__std__lane7_strm1_ready      ),      
               .std__pe40__lane7_strm1_cntl          ( std__pe40__lane7_strm1_cntl       ),      
               .std__pe40__lane7_strm1_data          ( std__pe40__lane7_strm1_data       ),      
               .std__pe40__lane7_strm1_data_valid    ( std__pe40__lane7_strm1_data_valid ),      
               .std__pe40__lane7_strm1_data_mask     ( std__pe40__lane7_strm1_data_mask  ),      

               // PE 40, Lane 8                 
               .pe40__std__lane8_strm0_ready         ( pe40__std__lane8_strm0_ready      ),      
               .std__pe40__lane8_strm0_cntl          ( std__pe40__lane8_strm0_cntl       ),      
               .std__pe40__lane8_strm0_data          ( std__pe40__lane8_strm0_data       ),      
               .std__pe40__lane8_strm0_data_valid    ( std__pe40__lane8_strm0_data_valid ),      
               .std__pe40__lane8_strm0_data_mask     ( std__pe40__lane8_strm0_data_mask  ),      

               .pe40__std__lane8_strm1_ready         ( pe40__std__lane8_strm1_ready      ),      
               .std__pe40__lane8_strm1_cntl          ( std__pe40__lane8_strm1_cntl       ),      
               .std__pe40__lane8_strm1_data          ( std__pe40__lane8_strm1_data       ),      
               .std__pe40__lane8_strm1_data_valid    ( std__pe40__lane8_strm1_data_valid ),      
               .std__pe40__lane8_strm1_data_mask     ( std__pe40__lane8_strm1_data_mask  ),      

               // PE 40, Lane 9                 
               .pe40__std__lane9_strm0_ready         ( pe40__std__lane9_strm0_ready      ),      
               .std__pe40__lane9_strm0_cntl          ( std__pe40__lane9_strm0_cntl       ),      
               .std__pe40__lane9_strm0_data          ( std__pe40__lane9_strm0_data       ),      
               .std__pe40__lane9_strm0_data_valid    ( std__pe40__lane9_strm0_data_valid ),      
               .std__pe40__lane9_strm0_data_mask     ( std__pe40__lane9_strm0_data_mask  ),      

               .pe40__std__lane9_strm1_ready         ( pe40__std__lane9_strm1_ready      ),      
               .std__pe40__lane9_strm1_cntl          ( std__pe40__lane9_strm1_cntl       ),      
               .std__pe40__lane9_strm1_data          ( std__pe40__lane9_strm1_data       ),      
               .std__pe40__lane9_strm1_data_valid    ( std__pe40__lane9_strm1_data_valid ),      
               .std__pe40__lane9_strm1_data_mask     ( std__pe40__lane9_strm1_data_mask  ),      

               // PE 40, Lane 10                 
               .pe40__std__lane10_strm0_ready         ( pe40__std__lane10_strm0_ready      ),      
               .std__pe40__lane10_strm0_cntl          ( std__pe40__lane10_strm0_cntl       ),      
               .std__pe40__lane10_strm0_data          ( std__pe40__lane10_strm0_data       ),      
               .std__pe40__lane10_strm0_data_valid    ( std__pe40__lane10_strm0_data_valid ),      
               .std__pe40__lane10_strm0_data_mask     ( std__pe40__lane10_strm0_data_mask  ),      

               .pe40__std__lane10_strm1_ready         ( pe40__std__lane10_strm1_ready      ),      
               .std__pe40__lane10_strm1_cntl          ( std__pe40__lane10_strm1_cntl       ),      
               .std__pe40__lane10_strm1_data          ( std__pe40__lane10_strm1_data       ),      
               .std__pe40__lane10_strm1_data_valid    ( std__pe40__lane10_strm1_data_valid ),      
               .std__pe40__lane10_strm1_data_mask     ( std__pe40__lane10_strm1_data_mask  ),      

               // PE 40, Lane 11                 
               .pe40__std__lane11_strm0_ready         ( pe40__std__lane11_strm0_ready      ),      
               .std__pe40__lane11_strm0_cntl          ( std__pe40__lane11_strm0_cntl       ),      
               .std__pe40__lane11_strm0_data          ( std__pe40__lane11_strm0_data       ),      
               .std__pe40__lane11_strm0_data_valid    ( std__pe40__lane11_strm0_data_valid ),      
               .std__pe40__lane11_strm0_data_mask     ( std__pe40__lane11_strm0_data_mask  ),      

               .pe40__std__lane11_strm1_ready         ( pe40__std__lane11_strm1_ready      ),      
               .std__pe40__lane11_strm1_cntl          ( std__pe40__lane11_strm1_cntl       ),      
               .std__pe40__lane11_strm1_data          ( std__pe40__lane11_strm1_data       ),      
               .std__pe40__lane11_strm1_data_valid    ( std__pe40__lane11_strm1_data_valid ),      
               .std__pe40__lane11_strm1_data_mask     ( std__pe40__lane11_strm1_data_mask  ),      

               // PE 40, Lane 12                 
               .pe40__std__lane12_strm0_ready         ( pe40__std__lane12_strm0_ready      ),      
               .std__pe40__lane12_strm0_cntl          ( std__pe40__lane12_strm0_cntl       ),      
               .std__pe40__lane12_strm0_data          ( std__pe40__lane12_strm0_data       ),      
               .std__pe40__lane12_strm0_data_valid    ( std__pe40__lane12_strm0_data_valid ),      
               .std__pe40__lane12_strm0_data_mask     ( std__pe40__lane12_strm0_data_mask  ),      

               .pe40__std__lane12_strm1_ready         ( pe40__std__lane12_strm1_ready      ),      
               .std__pe40__lane12_strm1_cntl          ( std__pe40__lane12_strm1_cntl       ),      
               .std__pe40__lane12_strm1_data          ( std__pe40__lane12_strm1_data       ),      
               .std__pe40__lane12_strm1_data_valid    ( std__pe40__lane12_strm1_data_valid ),      
               .std__pe40__lane12_strm1_data_mask     ( std__pe40__lane12_strm1_data_mask  ),      

               // PE 40, Lane 13                 
               .pe40__std__lane13_strm0_ready         ( pe40__std__lane13_strm0_ready      ),      
               .std__pe40__lane13_strm0_cntl          ( std__pe40__lane13_strm0_cntl       ),      
               .std__pe40__lane13_strm0_data          ( std__pe40__lane13_strm0_data       ),      
               .std__pe40__lane13_strm0_data_valid    ( std__pe40__lane13_strm0_data_valid ),      
               .std__pe40__lane13_strm0_data_mask     ( std__pe40__lane13_strm0_data_mask  ),      

               .pe40__std__lane13_strm1_ready         ( pe40__std__lane13_strm1_ready      ),      
               .std__pe40__lane13_strm1_cntl          ( std__pe40__lane13_strm1_cntl       ),      
               .std__pe40__lane13_strm1_data          ( std__pe40__lane13_strm1_data       ),      
               .std__pe40__lane13_strm1_data_valid    ( std__pe40__lane13_strm1_data_valid ),      
               .std__pe40__lane13_strm1_data_mask     ( std__pe40__lane13_strm1_data_mask  ),      

               // PE 40, Lane 14                 
               .pe40__std__lane14_strm0_ready         ( pe40__std__lane14_strm0_ready      ),      
               .std__pe40__lane14_strm0_cntl          ( std__pe40__lane14_strm0_cntl       ),      
               .std__pe40__lane14_strm0_data          ( std__pe40__lane14_strm0_data       ),      
               .std__pe40__lane14_strm0_data_valid    ( std__pe40__lane14_strm0_data_valid ),      
               .std__pe40__lane14_strm0_data_mask     ( std__pe40__lane14_strm0_data_mask  ),      

               .pe40__std__lane14_strm1_ready         ( pe40__std__lane14_strm1_ready      ),      
               .std__pe40__lane14_strm1_cntl          ( std__pe40__lane14_strm1_cntl       ),      
               .std__pe40__lane14_strm1_data          ( std__pe40__lane14_strm1_data       ),      
               .std__pe40__lane14_strm1_data_valid    ( std__pe40__lane14_strm1_data_valid ),      
               .std__pe40__lane14_strm1_data_mask     ( std__pe40__lane14_strm1_data_mask  ),      

               // PE 40, Lane 15                 
               .pe40__std__lane15_strm0_ready         ( pe40__std__lane15_strm0_ready      ),      
               .std__pe40__lane15_strm0_cntl          ( std__pe40__lane15_strm0_cntl       ),      
               .std__pe40__lane15_strm0_data          ( std__pe40__lane15_strm0_data       ),      
               .std__pe40__lane15_strm0_data_valid    ( std__pe40__lane15_strm0_data_valid ),      
               .std__pe40__lane15_strm0_data_mask     ( std__pe40__lane15_strm0_data_mask  ),      

               .pe40__std__lane15_strm1_ready         ( pe40__std__lane15_strm1_ready      ),      
               .std__pe40__lane15_strm1_cntl          ( std__pe40__lane15_strm1_cntl       ),      
               .std__pe40__lane15_strm1_data          ( std__pe40__lane15_strm1_data       ),      
               .std__pe40__lane15_strm1_data_valid    ( std__pe40__lane15_strm1_data_valid ),      
               .std__pe40__lane15_strm1_data_mask     ( std__pe40__lane15_strm1_data_mask  ),      

               // PE 40, Lane 16                 
               .pe40__std__lane16_strm0_ready         ( pe40__std__lane16_strm0_ready      ),      
               .std__pe40__lane16_strm0_cntl          ( std__pe40__lane16_strm0_cntl       ),      
               .std__pe40__lane16_strm0_data          ( std__pe40__lane16_strm0_data       ),      
               .std__pe40__lane16_strm0_data_valid    ( std__pe40__lane16_strm0_data_valid ),      
               .std__pe40__lane16_strm0_data_mask     ( std__pe40__lane16_strm0_data_mask  ),      

               .pe40__std__lane16_strm1_ready         ( pe40__std__lane16_strm1_ready      ),      
               .std__pe40__lane16_strm1_cntl          ( std__pe40__lane16_strm1_cntl       ),      
               .std__pe40__lane16_strm1_data          ( std__pe40__lane16_strm1_data       ),      
               .std__pe40__lane16_strm1_data_valid    ( std__pe40__lane16_strm1_data_valid ),      
               .std__pe40__lane16_strm1_data_mask     ( std__pe40__lane16_strm1_data_mask  ),      

               // PE 40, Lane 17                 
               .pe40__std__lane17_strm0_ready         ( pe40__std__lane17_strm0_ready      ),      
               .std__pe40__lane17_strm0_cntl          ( std__pe40__lane17_strm0_cntl       ),      
               .std__pe40__lane17_strm0_data          ( std__pe40__lane17_strm0_data       ),      
               .std__pe40__lane17_strm0_data_valid    ( std__pe40__lane17_strm0_data_valid ),      
               .std__pe40__lane17_strm0_data_mask     ( std__pe40__lane17_strm0_data_mask  ),      

               .pe40__std__lane17_strm1_ready         ( pe40__std__lane17_strm1_ready      ),      
               .std__pe40__lane17_strm1_cntl          ( std__pe40__lane17_strm1_cntl       ),      
               .std__pe40__lane17_strm1_data          ( std__pe40__lane17_strm1_data       ),      
               .std__pe40__lane17_strm1_data_valid    ( std__pe40__lane17_strm1_data_valid ),      
               .std__pe40__lane17_strm1_data_mask     ( std__pe40__lane17_strm1_data_mask  ),      

               // PE 40, Lane 18                 
               .pe40__std__lane18_strm0_ready         ( pe40__std__lane18_strm0_ready      ),      
               .std__pe40__lane18_strm0_cntl          ( std__pe40__lane18_strm0_cntl       ),      
               .std__pe40__lane18_strm0_data          ( std__pe40__lane18_strm0_data       ),      
               .std__pe40__lane18_strm0_data_valid    ( std__pe40__lane18_strm0_data_valid ),      
               .std__pe40__lane18_strm0_data_mask     ( std__pe40__lane18_strm0_data_mask  ),      

               .pe40__std__lane18_strm1_ready         ( pe40__std__lane18_strm1_ready      ),      
               .std__pe40__lane18_strm1_cntl          ( std__pe40__lane18_strm1_cntl       ),      
               .std__pe40__lane18_strm1_data          ( std__pe40__lane18_strm1_data       ),      
               .std__pe40__lane18_strm1_data_valid    ( std__pe40__lane18_strm1_data_valid ),      
               .std__pe40__lane18_strm1_data_mask     ( std__pe40__lane18_strm1_data_mask  ),      

               // PE 40, Lane 19                 
               .pe40__std__lane19_strm0_ready         ( pe40__std__lane19_strm0_ready      ),      
               .std__pe40__lane19_strm0_cntl          ( std__pe40__lane19_strm0_cntl       ),      
               .std__pe40__lane19_strm0_data          ( std__pe40__lane19_strm0_data       ),      
               .std__pe40__lane19_strm0_data_valid    ( std__pe40__lane19_strm0_data_valid ),      
               .std__pe40__lane19_strm0_data_mask     ( std__pe40__lane19_strm0_data_mask  ),      

               .pe40__std__lane19_strm1_ready         ( pe40__std__lane19_strm1_ready      ),      
               .std__pe40__lane19_strm1_cntl          ( std__pe40__lane19_strm1_cntl       ),      
               .std__pe40__lane19_strm1_data          ( std__pe40__lane19_strm1_data       ),      
               .std__pe40__lane19_strm1_data_valid    ( std__pe40__lane19_strm1_data_valid ),      
               .std__pe40__lane19_strm1_data_mask     ( std__pe40__lane19_strm1_data_mask  ),      

               // PE 40, Lane 20                 
               .pe40__std__lane20_strm0_ready         ( pe40__std__lane20_strm0_ready      ),      
               .std__pe40__lane20_strm0_cntl          ( std__pe40__lane20_strm0_cntl       ),      
               .std__pe40__lane20_strm0_data          ( std__pe40__lane20_strm0_data       ),      
               .std__pe40__lane20_strm0_data_valid    ( std__pe40__lane20_strm0_data_valid ),      
               .std__pe40__lane20_strm0_data_mask     ( std__pe40__lane20_strm0_data_mask  ),      

               .pe40__std__lane20_strm1_ready         ( pe40__std__lane20_strm1_ready      ),      
               .std__pe40__lane20_strm1_cntl          ( std__pe40__lane20_strm1_cntl       ),      
               .std__pe40__lane20_strm1_data          ( std__pe40__lane20_strm1_data       ),      
               .std__pe40__lane20_strm1_data_valid    ( std__pe40__lane20_strm1_data_valid ),      
               .std__pe40__lane20_strm1_data_mask     ( std__pe40__lane20_strm1_data_mask  ),      

               // PE 40, Lane 21                 
               .pe40__std__lane21_strm0_ready         ( pe40__std__lane21_strm0_ready      ),      
               .std__pe40__lane21_strm0_cntl          ( std__pe40__lane21_strm0_cntl       ),      
               .std__pe40__lane21_strm0_data          ( std__pe40__lane21_strm0_data       ),      
               .std__pe40__lane21_strm0_data_valid    ( std__pe40__lane21_strm0_data_valid ),      
               .std__pe40__lane21_strm0_data_mask     ( std__pe40__lane21_strm0_data_mask  ),      

               .pe40__std__lane21_strm1_ready         ( pe40__std__lane21_strm1_ready      ),      
               .std__pe40__lane21_strm1_cntl          ( std__pe40__lane21_strm1_cntl       ),      
               .std__pe40__lane21_strm1_data          ( std__pe40__lane21_strm1_data       ),      
               .std__pe40__lane21_strm1_data_valid    ( std__pe40__lane21_strm1_data_valid ),      
               .std__pe40__lane21_strm1_data_mask     ( std__pe40__lane21_strm1_data_mask  ),      

               // PE 40, Lane 22                 
               .pe40__std__lane22_strm0_ready         ( pe40__std__lane22_strm0_ready      ),      
               .std__pe40__lane22_strm0_cntl          ( std__pe40__lane22_strm0_cntl       ),      
               .std__pe40__lane22_strm0_data          ( std__pe40__lane22_strm0_data       ),      
               .std__pe40__lane22_strm0_data_valid    ( std__pe40__lane22_strm0_data_valid ),      
               .std__pe40__lane22_strm0_data_mask     ( std__pe40__lane22_strm0_data_mask  ),      

               .pe40__std__lane22_strm1_ready         ( pe40__std__lane22_strm1_ready      ),      
               .std__pe40__lane22_strm1_cntl          ( std__pe40__lane22_strm1_cntl       ),      
               .std__pe40__lane22_strm1_data          ( std__pe40__lane22_strm1_data       ),      
               .std__pe40__lane22_strm1_data_valid    ( std__pe40__lane22_strm1_data_valid ),      
               .std__pe40__lane22_strm1_data_mask     ( std__pe40__lane22_strm1_data_mask  ),      

               // PE 40, Lane 23                 
               .pe40__std__lane23_strm0_ready         ( pe40__std__lane23_strm0_ready      ),      
               .std__pe40__lane23_strm0_cntl          ( std__pe40__lane23_strm0_cntl       ),      
               .std__pe40__lane23_strm0_data          ( std__pe40__lane23_strm0_data       ),      
               .std__pe40__lane23_strm0_data_valid    ( std__pe40__lane23_strm0_data_valid ),      
               .std__pe40__lane23_strm0_data_mask     ( std__pe40__lane23_strm0_data_mask  ),      

               .pe40__std__lane23_strm1_ready         ( pe40__std__lane23_strm1_ready      ),      
               .std__pe40__lane23_strm1_cntl          ( std__pe40__lane23_strm1_cntl       ),      
               .std__pe40__lane23_strm1_data          ( std__pe40__lane23_strm1_data       ),      
               .std__pe40__lane23_strm1_data_valid    ( std__pe40__lane23_strm1_data_valid ),      
               .std__pe40__lane23_strm1_data_mask     ( std__pe40__lane23_strm1_data_mask  ),      

               // PE 40, Lane 24                 
               .pe40__std__lane24_strm0_ready         ( pe40__std__lane24_strm0_ready      ),      
               .std__pe40__lane24_strm0_cntl          ( std__pe40__lane24_strm0_cntl       ),      
               .std__pe40__lane24_strm0_data          ( std__pe40__lane24_strm0_data       ),      
               .std__pe40__lane24_strm0_data_valid    ( std__pe40__lane24_strm0_data_valid ),      
               .std__pe40__lane24_strm0_data_mask     ( std__pe40__lane24_strm0_data_mask  ),      

               .pe40__std__lane24_strm1_ready         ( pe40__std__lane24_strm1_ready      ),      
               .std__pe40__lane24_strm1_cntl          ( std__pe40__lane24_strm1_cntl       ),      
               .std__pe40__lane24_strm1_data          ( std__pe40__lane24_strm1_data       ),      
               .std__pe40__lane24_strm1_data_valid    ( std__pe40__lane24_strm1_data_valid ),      
               .std__pe40__lane24_strm1_data_mask     ( std__pe40__lane24_strm1_data_mask  ),      

               // PE 40, Lane 25                 
               .pe40__std__lane25_strm0_ready         ( pe40__std__lane25_strm0_ready      ),      
               .std__pe40__lane25_strm0_cntl          ( std__pe40__lane25_strm0_cntl       ),      
               .std__pe40__lane25_strm0_data          ( std__pe40__lane25_strm0_data       ),      
               .std__pe40__lane25_strm0_data_valid    ( std__pe40__lane25_strm0_data_valid ),      
               .std__pe40__lane25_strm0_data_mask     ( std__pe40__lane25_strm0_data_mask  ),      

               .pe40__std__lane25_strm1_ready         ( pe40__std__lane25_strm1_ready      ),      
               .std__pe40__lane25_strm1_cntl          ( std__pe40__lane25_strm1_cntl       ),      
               .std__pe40__lane25_strm1_data          ( std__pe40__lane25_strm1_data       ),      
               .std__pe40__lane25_strm1_data_valid    ( std__pe40__lane25_strm1_data_valid ),      
               .std__pe40__lane25_strm1_data_mask     ( std__pe40__lane25_strm1_data_mask  ),      

               // PE 40, Lane 26                 
               .pe40__std__lane26_strm0_ready         ( pe40__std__lane26_strm0_ready      ),      
               .std__pe40__lane26_strm0_cntl          ( std__pe40__lane26_strm0_cntl       ),      
               .std__pe40__lane26_strm0_data          ( std__pe40__lane26_strm0_data       ),      
               .std__pe40__lane26_strm0_data_valid    ( std__pe40__lane26_strm0_data_valid ),      
               .std__pe40__lane26_strm0_data_mask     ( std__pe40__lane26_strm0_data_mask  ),      

               .pe40__std__lane26_strm1_ready         ( pe40__std__lane26_strm1_ready      ),      
               .std__pe40__lane26_strm1_cntl          ( std__pe40__lane26_strm1_cntl       ),      
               .std__pe40__lane26_strm1_data          ( std__pe40__lane26_strm1_data       ),      
               .std__pe40__lane26_strm1_data_valid    ( std__pe40__lane26_strm1_data_valid ),      
               .std__pe40__lane26_strm1_data_mask     ( std__pe40__lane26_strm1_data_mask  ),      

               // PE 40, Lane 27                 
               .pe40__std__lane27_strm0_ready         ( pe40__std__lane27_strm0_ready      ),      
               .std__pe40__lane27_strm0_cntl          ( std__pe40__lane27_strm0_cntl       ),      
               .std__pe40__lane27_strm0_data          ( std__pe40__lane27_strm0_data       ),      
               .std__pe40__lane27_strm0_data_valid    ( std__pe40__lane27_strm0_data_valid ),      
               .std__pe40__lane27_strm0_data_mask     ( std__pe40__lane27_strm0_data_mask  ),      

               .pe40__std__lane27_strm1_ready         ( pe40__std__lane27_strm1_ready      ),      
               .std__pe40__lane27_strm1_cntl          ( std__pe40__lane27_strm1_cntl       ),      
               .std__pe40__lane27_strm1_data          ( std__pe40__lane27_strm1_data       ),      
               .std__pe40__lane27_strm1_data_valid    ( std__pe40__lane27_strm1_data_valid ),      
               .std__pe40__lane27_strm1_data_mask     ( std__pe40__lane27_strm1_data_mask  ),      

               // PE 40, Lane 28                 
               .pe40__std__lane28_strm0_ready         ( pe40__std__lane28_strm0_ready      ),      
               .std__pe40__lane28_strm0_cntl          ( std__pe40__lane28_strm0_cntl       ),      
               .std__pe40__lane28_strm0_data          ( std__pe40__lane28_strm0_data       ),      
               .std__pe40__lane28_strm0_data_valid    ( std__pe40__lane28_strm0_data_valid ),      
               .std__pe40__lane28_strm0_data_mask     ( std__pe40__lane28_strm0_data_mask  ),      

               .pe40__std__lane28_strm1_ready         ( pe40__std__lane28_strm1_ready      ),      
               .std__pe40__lane28_strm1_cntl          ( std__pe40__lane28_strm1_cntl       ),      
               .std__pe40__lane28_strm1_data          ( std__pe40__lane28_strm1_data       ),      
               .std__pe40__lane28_strm1_data_valid    ( std__pe40__lane28_strm1_data_valid ),      
               .std__pe40__lane28_strm1_data_mask     ( std__pe40__lane28_strm1_data_mask  ),      

               // PE 40, Lane 29                 
               .pe40__std__lane29_strm0_ready         ( pe40__std__lane29_strm0_ready      ),      
               .std__pe40__lane29_strm0_cntl          ( std__pe40__lane29_strm0_cntl       ),      
               .std__pe40__lane29_strm0_data          ( std__pe40__lane29_strm0_data       ),      
               .std__pe40__lane29_strm0_data_valid    ( std__pe40__lane29_strm0_data_valid ),      
               .std__pe40__lane29_strm0_data_mask     ( std__pe40__lane29_strm0_data_mask  ),      

               .pe40__std__lane29_strm1_ready         ( pe40__std__lane29_strm1_ready      ),      
               .std__pe40__lane29_strm1_cntl          ( std__pe40__lane29_strm1_cntl       ),      
               .std__pe40__lane29_strm1_data          ( std__pe40__lane29_strm1_data       ),      
               .std__pe40__lane29_strm1_data_valid    ( std__pe40__lane29_strm1_data_valid ),      
               .std__pe40__lane29_strm1_data_mask     ( std__pe40__lane29_strm1_data_mask  ),      

               // PE 40, Lane 30                 
               .pe40__std__lane30_strm0_ready         ( pe40__std__lane30_strm0_ready      ),      
               .std__pe40__lane30_strm0_cntl          ( std__pe40__lane30_strm0_cntl       ),      
               .std__pe40__lane30_strm0_data          ( std__pe40__lane30_strm0_data       ),      
               .std__pe40__lane30_strm0_data_valid    ( std__pe40__lane30_strm0_data_valid ),      
               .std__pe40__lane30_strm0_data_mask     ( std__pe40__lane30_strm0_data_mask  ),      

               .pe40__std__lane30_strm1_ready         ( pe40__std__lane30_strm1_ready      ),      
               .std__pe40__lane30_strm1_cntl          ( std__pe40__lane30_strm1_cntl       ),      
               .std__pe40__lane30_strm1_data          ( std__pe40__lane30_strm1_data       ),      
               .std__pe40__lane30_strm1_data_valid    ( std__pe40__lane30_strm1_data_valid ),      
               .std__pe40__lane30_strm1_data_mask     ( std__pe40__lane30_strm1_data_mask  ),      

               // PE 40, Lane 31                 
               .pe40__std__lane31_strm0_ready         ( pe40__std__lane31_strm0_ready      ),      
               .std__pe40__lane31_strm0_cntl          ( std__pe40__lane31_strm0_cntl       ),      
               .std__pe40__lane31_strm0_data          ( std__pe40__lane31_strm0_data       ),      
               .std__pe40__lane31_strm0_data_valid    ( std__pe40__lane31_strm0_data_valid ),      
               .std__pe40__lane31_strm0_data_mask     ( std__pe40__lane31_strm0_data_mask  ),      

               .pe40__std__lane31_strm1_ready         ( pe40__std__lane31_strm1_ready      ),      
               .std__pe40__lane31_strm1_cntl          ( std__pe40__lane31_strm1_cntl       ),      
               .std__pe40__lane31_strm1_data          ( std__pe40__lane31_strm1_data       ),      
               .std__pe40__lane31_strm1_data_valid    ( std__pe40__lane31_strm1_data_valid ),      
               .std__pe40__lane31_strm1_data_mask     ( std__pe40__lane31_strm1_data_mask  ),      

               // PE 41, Lane 0                 
               .pe41__std__lane0_strm0_ready         ( pe41__std__lane0_strm0_ready      ),      
               .std__pe41__lane0_strm0_cntl          ( std__pe41__lane0_strm0_cntl       ),      
               .std__pe41__lane0_strm0_data          ( std__pe41__lane0_strm0_data       ),      
               .std__pe41__lane0_strm0_data_valid    ( std__pe41__lane0_strm0_data_valid ),      
               .std__pe41__lane0_strm0_data_mask     ( std__pe41__lane0_strm0_data_mask  ),      

               .pe41__std__lane0_strm1_ready         ( pe41__std__lane0_strm1_ready      ),      
               .std__pe41__lane0_strm1_cntl          ( std__pe41__lane0_strm1_cntl       ),      
               .std__pe41__lane0_strm1_data          ( std__pe41__lane0_strm1_data       ),      
               .std__pe41__lane0_strm1_data_valid    ( std__pe41__lane0_strm1_data_valid ),      
               .std__pe41__lane0_strm1_data_mask     ( std__pe41__lane0_strm1_data_mask  ),      

               // PE 41, Lane 1                 
               .pe41__std__lane1_strm0_ready         ( pe41__std__lane1_strm0_ready      ),      
               .std__pe41__lane1_strm0_cntl          ( std__pe41__lane1_strm0_cntl       ),      
               .std__pe41__lane1_strm0_data          ( std__pe41__lane1_strm0_data       ),      
               .std__pe41__lane1_strm0_data_valid    ( std__pe41__lane1_strm0_data_valid ),      
               .std__pe41__lane1_strm0_data_mask     ( std__pe41__lane1_strm0_data_mask  ),      

               .pe41__std__lane1_strm1_ready         ( pe41__std__lane1_strm1_ready      ),      
               .std__pe41__lane1_strm1_cntl          ( std__pe41__lane1_strm1_cntl       ),      
               .std__pe41__lane1_strm1_data          ( std__pe41__lane1_strm1_data       ),      
               .std__pe41__lane1_strm1_data_valid    ( std__pe41__lane1_strm1_data_valid ),      
               .std__pe41__lane1_strm1_data_mask     ( std__pe41__lane1_strm1_data_mask  ),      

               // PE 41, Lane 2                 
               .pe41__std__lane2_strm0_ready         ( pe41__std__lane2_strm0_ready      ),      
               .std__pe41__lane2_strm0_cntl          ( std__pe41__lane2_strm0_cntl       ),      
               .std__pe41__lane2_strm0_data          ( std__pe41__lane2_strm0_data       ),      
               .std__pe41__lane2_strm0_data_valid    ( std__pe41__lane2_strm0_data_valid ),      
               .std__pe41__lane2_strm0_data_mask     ( std__pe41__lane2_strm0_data_mask  ),      

               .pe41__std__lane2_strm1_ready         ( pe41__std__lane2_strm1_ready      ),      
               .std__pe41__lane2_strm1_cntl          ( std__pe41__lane2_strm1_cntl       ),      
               .std__pe41__lane2_strm1_data          ( std__pe41__lane2_strm1_data       ),      
               .std__pe41__lane2_strm1_data_valid    ( std__pe41__lane2_strm1_data_valid ),      
               .std__pe41__lane2_strm1_data_mask     ( std__pe41__lane2_strm1_data_mask  ),      

               // PE 41, Lane 3                 
               .pe41__std__lane3_strm0_ready         ( pe41__std__lane3_strm0_ready      ),      
               .std__pe41__lane3_strm0_cntl          ( std__pe41__lane3_strm0_cntl       ),      
               .std__pe41__lane3_strm0_data          ( std__pe41__lane3_strm0_data       ),      
               .std__pe41__lane3_strm0_data_valid    ( std__pe41__lane3_strm0_data_valid ),      
               .std__pe41__lane3_strm0_data_mask     ( std__pe41__lane3_strm0_data_mask  ),      

               .pe41__std__lane3_strm1_ready         ( pe41__std__lane3_strm1_ready      ),      
               .std__pe41__lane3_strm1_cntl          ( std__pe41__lane3_strm1_cntl       ),      
               .std__pe41__lane3_strm1_data          ( std__pe41__lane3_strm1_data       ),      
               .std__pe41__lane3_strm1_data_valid    ( std__pe41__lane3_strm1_data_valid ),      
               .std__pe41__lane3_strm1_data_mask     ( std__pe41__lane3_strm1_data_mask  ),      

               // PE 41, Lane 4                 
               .pe41__std__lane4_strm0_ready         ( pe41__std__lane4_strm0_ready      ),      
               .std__pe41__lane4_strm0_cntl          ( std__pe41__lane4_strm0_cntl       ),      
               .std__pe41__lane4_strm0_data          ( std__pe41__lane4_strm0_data       ),      
               .std__pe41__lane4_strm0_data_valid    ( std__pe41__lane4_strm0_data_valid ),      
               .std__pe41__lane4_strm0_data_mask     ( std__pe41__lane4_strm0_data_mask  ),      

               .pe41__std__lane4_strm1_ready         ( pe41__std__lane4_strm1_ready      ),      
               .std__pe41__lane4_strm1_cntl          ( std__pe41__lane4_strm1_cntl       ),      
               .std__pe41__lane4_strm1_data          ( std__pe41__lane4_strm1_data       ),      
               .std__pe41__lane4_strm1_data_valid    ( std__pe41__lane4_strm1_data_valid ),      
               .std__pe41__lane4_strm1_data_mask     ( std__pe41__lane4_strm1_data_mask  ),      

               // PE 41, Lane 5                 
               .pe41__std__lane5_strm0_ready         ( pe41__std__lane5_strm0_ready      ),      
               .std__pe41__lane5_strm0_cntl          ( std__pe41__lane5_strm0_cntl       ),      
               .std__pe41__lane5_strm0_data          ( std__pe41__lane5_strm0_data       ),      
               .std__pe41__lane5_strm0_data_valid    ( std__pe41__lane5_strm0_data_valid ),      
               .std__pe41__lane5_strm0_data_mask     ( std__pe41__lane5_strm0_data_mask  ),      

               .pe41__std__lane5_strm1_ready         ( pe41__std__lane5_strm1_ready      ),      
               .std__pe41__lane5_strm1_cntl          ( std__pe41__lane5_strm1_cntl       ),      
               .std__pe41__lane5_strm1_data          ( std__pe41__lane5_strm1_data       ),      
               .std__pe41__lane5_strm1_data_valid    ( std__pe41__lane5_strm1_data_valid ),      
               .std__pe41__lane5_strm1_data_mask     ( std__pe41__lane5_strm1_data_mask  ),      

               // PE 41, Lane 6                 
               .pe41__std__lane6_strm0_ready         ( pe41__std__lane6_strm0_ready      ),      
               .std__pe41__lane6_strm0_cntl          ( std__pe41__lane6_strm0_cntl       ),      
               .std__pe41__lane6_strm0_data          ( std__pe41__lane6_strm0_data       ),      
               .std__pe41__lane6_strm0_data_valid    ( std__pe41__lane6_strm0_data_valid ),      
               .std__pe41__lane6_strm0_data_mask     ( std__pe41__lane6_strm0_data_mask  ),      

               .pe41__std__lane6_strm1_ready         ( pe41__std__lane6_strm1_ready      ),      
               .std__pe41__lane6_strm1_cntl          ( std__pe41__lane6_strm1_cntl       ),      
               .std__pe41__lane6_strm1_data          ( std__pe41__lane6_strm1_data       ),      
               .std__pe41__lane6_strm1_data_valid    ( std__pe41__lane6_strm1_data_valid ),      
               .std__pe41__lane6_strm1_data_mask     ( std__pe41__lane6_strm1_data_mask  ),      

               // PE 41, Lane 7                 
               .pe41__std__lane7_strm0_ready         ( pe41__std__lane7_strm0_ready      ),      
               .std__pe41__lane7_strm0_cntl          ( std__pe41__lane7_strm0_cntl       ),      
               .std__pe41__lane7_strm0_data          ( std__pe41__lane7_strm0_data       ),      
               .std__pe41__lane7_strm0_data_valid    ( std__pe41__lane7_strm0_data_valid ),      
               .std__pe41__lane7_strm0_data_mask     ( std__pe41__lane7_strm0_data_mask  ),      

               .pe41__std__lane7_strm1_ready         ( pe41__std__lane7_strm1_ready      ),      
               .std__pe41__lane7_strm1_cntl          ( std__pe41__lane7_strm1_cntl       ),      
               .std__pe41__lane7_strm1_data          ( std__pe41__lane7_strm1_data       ),      
               .std__pe41__lane7_strm1_data_valid    ( std__pe41__lane7_strm1_data_valid ),      
               .std__pe41__lane7_strm1_data_mask     ( std__pe41__lane7_strm1_data_mask  ),      

               // PE 41, Lane 8                 
               .pe41__std__lane8_strm0_ready         ( pe41__std__lane8_strm0_ready      ),      
               .std__pe41__lane8_strm0_cntl          ( std__pe41__lane8_strm0_cntl       ),      
               .std__pe41__lane8_strm0_data          ( std__pe41__lane8_strm0_data       ),      
               .std__pe41__lane8_strm0_data_valid    ( std__pe41__lane8_strm0_data_valid ),      
               .std__pe41__lane8_strm0_data_mask     ( std__pe41__lane8_strm0_data_mask  ),      

               .pe41__std__lane8_strm1_ready         ( pe41__std__lane8_strm1_ready      ),      
               .std__pe41__lane8_strm1_cntl          ( std__pe41__lane8_strm1_cntl       ),      
               .std__pe41__lane8_strm1_data          ( std__pe41__lane8_strm1_data       ),      
               .std__pe41__lane8_strm1_data_valid    ( std__pe41__lane8_strm1_data_valid ),      
               .std__pe41__lane8_strm1_data_mask     ( std__pe41__lane8_strm1_data_mask  ),      

               // PE 41, Lane 9                 
               .pe41__std__lane9_strm0_ready         ( pe41__std__lane9_strm0_ready      ),      
               .std__pe41__lane9_strm0_cntl          ( std__pe41__lane9_strm0_cntl       ),      
               .std__pe41__lane9_strm0_data          ( std__pe41__lane9_strm0_data       ),      
               .std__pe41__lane9_strm0_data_valid    ( std__pe41__lane9_strm0_data_valid ),      
               .std__pe41__lane9_strm0_data_mask     ( std__pe41__lane9_strm0_data_mask  ),      

               .pe41__std__lane9_strm1_ready         ( pe41__std__lane9_strm1_ready      ),      
               .std__pe41__lane9_strm1_cntl          ( std__pe41__lane9_strm1_cntl       ),      
               .std__pe41__lane9_strm1_data          ( std__pe41__lane9_strm1_data       ),      
               .std__pe41__lane9_strm1_data_valid    ( std__pe41__lane9_strm1_data_valid ),      
               .std__pe41__lane9_strm1_data_mask     ( std__pe41__lane9_strm1_data_mask  ),      

               // PE 41, Lane 10                 
               .pe41__std__lane10_strm0_ready         ( pe41__std__lane10_strm0_ready      ),      
               .std__pe41__lane10_strm0_cntl          ( std__pe41__lane10_strm0_cntl       ),      
               .std__pe41__lane10_strm0_data          ( std__pe41__lane10_strm0_data       ),      
               .std__pe41__lane10_strm0_data_valid    ( std__pe41__lane10_strm0_data_valid ),      
               .std__pe41__lane10_strm0_data_mask     ( std__pe41__lane10_strm0_data_mask  ),      

               .pe41__std__lane10_strm1_ready         ( pe41__std__lane10_strm1_ready      ),      
               .std__pe41__lane10_strm1_cntl          ( std__pe41__lane10_strm1_cntl       ),      
               .std__pe41__lane10_strm1_data          ( std__pe41__lane10_strm1_data       ),      
               .std__pe41__lane10_strm1_data_valid    ( std__pe41__lane10_strm1_data_valid ),      
               .std__pe41__lane10_strm1_data_mask     ( std__pe41__lane10_strm1_data_mask  ),      

               // PE 41, Lane 11                 
               .pe41__std__lane11_strm0_ready         ( pe41__std__lane11_strm0_ready      ),      
               .std__pe41__lane11_strm0_cntl          ( std__pe41__lane11_strm0_cntl       ),      
               .std__pe41__lane11_strm0_data          ( std__pe41__lane11_strm0_data       ),      
               .std__pe41__lane11_strm0_data_valid    ( std__pe41__lane11_strm0_data_valid ),      
               .std__pe41__lane11_strm0_data_mask     ( std__pe41__lane11_strm0_data_mask  ),      

               .pe41__std__lane11_strm1_ready         ( pe41__std__lane11_strm1_ready      ),      
               .std__pe41__lane11_strm1_cntl          ( std__pe41__lane11_strm1_cntl       ),      
               .std__pe41__lane11_strm1_data          ( std__pe41__lane11_strm1_data       ),      
               .std__pe41__lane11_strm1_data_valid    ( std__pe41__lane11_strm1_data_valid ),      
               .std__pe41__lane11_strm1_data_mask     ( std__pe41__lane11_strm1_data_mask  ),      

               // PE 41, Lane 12                 
               .pe41__std__lane12_strm0_ready         ( pe41__std__lane12_strm0_ready      ),      
               .std__pe41__lane12_strm0_cntl          ( std__pe41__lane12_strm0_cntl       ),      
               .std__pe41__lane12_strm0_data          ( std__pe41__lane12_strm0_data       ),      
               .std__pe41__lane12_strm0_data_valid    ( std__pe41__lane12_strm0_data_valid ),      
               .std__pe41__lane12_strm0_data_mask     ( std__pe41__lane12_strm0_data_mask  ),      

               .pe41__std__lane12_strm1_ready         ( pe41__std__lane12_strm1_ready      ),      
               .std__pe41__lane12_strm1_cntl          ( std__pe41__lane12_strm1_cntl       ),      
               .std__pe41__lane12_strm1_data          ( std__pe41__lane12_strm1_data       ),      
               .std__pe41__lane12_strm1_data_valid    ( std__pe41__lane12_strm1_data_valid ),      
               .std__pe41__lane12_strm1_data_mask     ( std__pe41__lane12_strm1_data_mask  ),      

               // PE 41, Lane 13                 
               .pe41__std__lane13_strm0_ready         ( pe41__std__lane13_strm0_ready      ),      
               .std__pe41__lane13_strm0_cntl          ( std__pe41__lane13_strm0_cntl       ),      
               .std__pe41__lane13_strm0_data          ( std__pe41__lane13_strm0_data       ),      
               .std__pe41__lane13_strm0_data_valid    ( std__pe41__lane13_strm0_data_valid ),      
               .std__pe41__lane13_strm0_data_mask     ( std__pe41__lane13_strm0_data_mask  ),      

               .pe41__std__lane13_strm1_ready         ( pe41__std__lane13_strm1_ready      ),      
               .std__pe41__lane13_strm1_cntl          ( std__pe41__lane13_strm1_cntl       ),      
               .std__pe41__lane13_strm1_data          ( std__pe41__lane13_strm1_data       ),      
               .std__pe41__lane13_strm1_data_valid    ( std__pe41__lane13_strm1_data_valid ),      
               .std__pe41__lane13_strm1_data_mask     ( std__pe41__lane13_strm1_data_mask  ),      

               // PE 41, Lane 14                 
               .pe41__std__lane14_strm0_ready         ( pe41__std__lane14_strm0_ready      ),      
               .std__pe41__lane14_strm0_cntl          ( std__pe41__lane14_strm0_cntl       ),      
               .std__pe41__lane14_strm0_data          ( std__pe41__lane14_strm0_data       ),      
               .std__pe41__lane14_strm0_data_valid    ( std__pe41__lane14_strm0_data_valid ),      
               .std__pe41__lane14_strm0_data_mask     ( std__pe41__lane14_strm0_data_mask  ),      

               .pe41__std__lane14_strm1_ready         ( pe41__std__lane14_strm1_ready      ),      
               .std__pe41__lane14_strm1_cntl          ( std__pe41__lane14_strm1_cntl       ),      
               .std__pe41__lane14_strm1_data          ( std__pe41__lane14_strm1_data       ),      
               .std__pe41__lane14_strm1_data_valid    ( std__pe41__lane14_strm1_data_valid ),      
               .std__pe41__lane14_strm1_data_mask     ( std__pe41__lane14_strm1_data_mask  ),      

               // PE 41, Lane 15                 
               .pe41__std__lane15_strm0_ready         ( pe41__std__lane15_strm0_ready      ),      
               .std__pe41__lane15_strm0_cntl          ( std__pe41__lane15_strm0_cntl       ),      
               .std__pe41__lane15_strm0_data          ( std__pe41__lane15_strm0_data       ),      
               .std__pe41__lane15_strm0_data_valid    ( std__pe41__lane15_strm0_data_valid ),      
               .std__pe41__lane15_strm0_data_mask     ( std__pe41__lane15_strm0_data_mask  ),      

               .pe41__std__lane15_strm1_ready         ( pe41__std__lane15_strm1_ready      ),      
               .std__pe41__lane15_strm1_cntl          ( std__pe41__lane15_strm1_cntl       ),      
               .std__pe41__lane15_strm1_data          ( std__pe41__lane15_strm1_data       ),      
               .std__pe41__lane15_strm1_data_valid    ( std__pe41__lane15_strm1_data_valid ),      
               .std__pe41__lane15_strm1_data_mask     ( std__pe41__lane15_strm1_data_mask  ),      

               // PE 41, Lane 16                 
               .pe41__std__lane16_strm0_ready         ( pe41__std__lane16_strm0_ready      ),      
               .std__pe41__lane16_strm0_cntl          ( std__pe41__lane16_strm0_cntl       ),      
               .std__pe41__lane16_strm0_data          ( std__pe41__lane16_strm0_data       ),      
               .std__pe41__lane16_strm0_data_valid    ( std__pe41__lane16_strm0_data_valid ),      
               .std__pe41__lane16_strm0_data_mask     ( std__pe41__lane16_strm0_data_mask  ),      

               .pe41__std__lane16_strm1_ready         ( pe41__std__lane16_strm1_ready      ),      
               .std__pe41__lane16_strm1_cntl          ( std__pe41__lane16_strm1_cntl       ),      
               .std__pe41__lane16_strm1_data          ( std__pe41__lane16_strm1_data       ),      
               .std__pe41__lane16_strm1_data_valid    ( std__pe41__lane16_strm1_data_valid ),      
               .std__pe41__lane16_strm1_data_mask     ( std__pe41__lane16_strm1_data_mask  ),      

               // PE 41, Lane 17                 
               .pe41__std__lane17_strm0_ready         ( pe41__std__lane17_strm0_ready      ),      
               .std__pe41__lane17_strm0_cntl          ( std__pe41__lane17_strm0_cntl       ),      
               .std__pe41__lane17_strm0_data          ( std__pe41__lane17_strm0_data       ),      
               .std__pe41__lane17_strm0_data_valid    ( std__pe41__lane17_strm0_data_valid ),      
               .std__pe41__lane17_strm0_data_mask     ( std__pe41__lane17_strm0_data_mask  ),      

               .pe41__std__lane17_strm1_ready         ( pe41__std__lane17_strm1_ready      ),      
               .std__pe41__lane17_strm1_cntl          ( std__pe41__lane17_strm1_cntl       ),      
               .std__pe41__lane17_strm1_data          ( std__pe41__lane17_strm1_data       ),      
               .std__pe41__lane17_strm1_data_valid    ( std__pe41__lane17_strm1_data_valid ),      
               .std__pe41__lane17_strm1_data_mask     ( std__pe41__lane17_strm1_data_mask  ),      

               // PE 41, Lane 18                 
               .pe41__std__lane18_strm0_ready         ( pe41__std__lane18_strm0_ready      ),      
               .std__pe41__lane18_strm0_cntl          ( std__pe41__lane18_strm0_cntl       ),      
               .std__pe41__lane18_strm0_data          ( std__pe41__lane18_strm0_data       ),      
               .std__pe41__lane18_strm0_data_valid    ( std__pe41__lane18_strm0_data_valid ),      
               .std__pe41__lane18_strm0_data_mask     ( std__pe41__lane18_strm0_data_mask  ),      

               .pe41__std__lane18_strm1_ready         ( pe41__std__lane18_strm1_ready      ),      
               .std__pe41__lane18_strm1_cntl          ( std__pe41__lane18_strm1_cntl       ),      
               .std__pe41__lane18_strm1_data          ( std__pe41__lane18_strm1_data       ),      
               .std__pe41__lane18_strm1_data_valid    ( std__pe41__lane18_strm1_data_valid ),      
               .std__pe41__lane18_strm1_data_mask     ( std__pe41__lane18_strm1_data_mask  ),      

               // PE 41, Lane 19                 
               .pe41__std__lane19_strm0_ready         ( pe41__std__lane19_strm0_ready      ),      
               .std__pe41__lane19_strm0_cntl          ( std__pe41__lane19_strm0_cntl       ),      
               .std__pe41__lane19_strm0_data          ( std__pe41__lane19_strm0_data       ),      
               .std__pe41__lane19_strm0_data_valid    ( std__pe41__lane19_strm0_data_valid ),      
               .std__pe41__lane19_strm0_data_mask     ( std__pe41__lane19_strm0_data_mask  ),      

               .pe41__std__lane19_strm1_ready         ( pe41__std__lane19_strm1_ready      ),      
               .std__pe41__lane19_strm1_cntl          ( std__pe41__lane19_strm1_cntl       ),      
               .std__pe41__lane19_strm1_data          ( std__pe41__lane19_strm1_data       ),      
               .std__pe41__lane19_strm1_data_valid    ( std__pe41__lane19_strm1_data_valid ),      
               .std__pe41__lane19_strm1_data_mask     ( std__pe41__lane19_strm1_data_mask  ),      

               // PE 41, Lane 20                 
               .pe41__std__lane20_strm0_ready         ( pe41__std__lane20_strm0_ready      ),      
               .std__pe41__lane20_strm0_cntl          ( std__pe41__lane20_strm0_cntl       ),      
               .std__pe41__lane20_strm0_data          ( std__pe41__lane20_strm0_data       ),      
               .std__pe41__lane20_strm0_data_valid    ( std__pe41__lane20_strm0_data_valid ),      
               .std__pe41__lane20_strm0_data_mask     ( std__pe41__lane20_strm0_data_mask  ),      

               .pe41__std__lane20_strm1_ready         ( pe41__std__lane20_strm1_ready      ),      
               .std__pe41__lane20_strm1_cntl          ( std__pe41__lane20_strm1_cntl       ),      
               .std__pe41__lane20_strm1_data          ( std__pe41__lane20_strm1_data       ),      
               .std__pe41__lane20_strm1_data_valid    ( std__pe41__lane20_strm1_data_valid ),      
               .std__pe41__lane20_strm1_data_mask     ( std__pe41__lane20_strm1_data_mask  ),      

               // PE 41, Lane 21                 
               .pe41__std__lane21_strm0_ready         ( pe41__std__lane21_strm0_ready      ),      
               .std__pe41__lane21_strm0_cntl          ( std__pe41__lane21_strm0_cntl       ),      
               .std__pe41__lane21_strm0_data          ( std__pe41__lane21_strm0_data       ),      
               .std__pe41__lane21_strm0_data_valid    ( std__pe41__lane21_strm0_data_valid ),      
               .std__pe41__lane21_strm0_data_mask     ( std__pe41__lane21_strm0_data_mask  ),      

               .pe41__std__lane21_strm1_ready         ( pe41__std__lane21_strm1_ready      ),      
               .std__pe41__lane21_strm1_cntl          ( std__pe41__lane21_strm1_cntl       ),      
               .std__pe41__lane21_strm1_data          ( std__pe41__lane21_strm1_data       ),      
               .std__pe41__lane21_strm1_data_valid    ( std__pe41__lane21_strm1_data_valid ),      
               .std__pe41__lane21_strm1_data_mask     ( std__pe41__lane21_strm1_data_mask  ),      

               // PE 41, Lane 22                 
               .pe41__std__lane22_strm0_ready         ( pe41__std__lane22_strm0_ready      ),      
               .std__pe41__lane22_strm0_cntl          ( std__pe41__lane22_strm0_cntl       ),      
               .std__pe41__lane22_strm0_data          ( std__pe41__lane22_strm0_data       ),      
               .std__pe41__lane22_strm0_data_valid    ( std__pe41__lane22_strm0_data_valid ),      
               .std__pe41__lane22_strm0_data_mask     ( std__pe41__lane22_strm0_data_mask  ),      

               .pe41__std__lane22_strm1_ready         ( pe41__std__lane22_strm1_ready      ),      
               .std__pe41__lane22_strm1_cntl          ( std__pe41__lane22_strm1_cntl       ),      
               .std__pe41__lane22_strm1_data          ( std__pe41__lane22_strm1_data       ),      
               .std__pe41__lane22_strm1_data_valid    ( std__pe41__lane22_strm1_data_valid ),      
               .std__pe41__lane22_strm1_data_mask     ( std__pe41__lane22_strm1_data_mask  ),      

               // PE 41, Lane 23                 
               .pe41__std__lane23_strm0_ready         ( pe41__std__lane23_strm0_ready      ),      
               .std__pe41__lane23_strm0_cntl          ( std__pe41__lane23_strm0_cntl       ),      
               .std__pe41__lane23_strm0_data          ( std__pe41__lane23_strm0_data       ),      
               .std__pe41__lane23_strm0_data_valid    ( std__pe41__lane23_strm0_data_valid ),      
               .std__pe41__lane23_strm0_data_mask     ( std__pe41__lane23_strm0_data_mask  ),      

               .pe41__std__lane23_strm1_ready         ( pe41__std__lane23_strm1_ready      ),      
               .std__pe41__lane23_strm1_cntl          ( std__pe41__lane23_strm1_cntl       ),      
               .std__pe41__lane23_strm1_data          ( std__pe41__lane23_strm1_data       ),      
               .std__pe41__lane23_strm1_data_valid    ( std__pe41__lane23_strm1_data_valid ),      
               .std__pe41__lane23_strm1_data_mask     ( std__pe41__lane23_strm1_data_mask  ),      

               // PE 41, Lane 24                 
               .pe41__std__lane24_strm0_ready         ( pe41__std__lane24_strm0_ready      ),      
               .std__pe41__lane24_strm0_cntl          ( std__pe41__lane24_strm0_cntl       ),      
               .std__pe41__lane24_strm0_data          ( std__pe41__lane24_strm0_data       ),      
               .std__pe41__lane24_strm0_data_valid    ( std__pe41__lane24_strm0_data_valid ),      
               .std__pe41__lane24_strm0_data_mask     ( std__pe41__lane24_strm0_data_mask  ),      

               .pe41__std__lane24_strm1_ready         ( pe41__std__lane24_strm1_ready      ),      
               .std__pe41__lane24_strm1_cntl          ( std__pe41__lane24_strm1_cntl       ),      
               .std__pe41__lane24_strm1_data          ( std__pe41__lane24_strm1_data       ),      
               .std__pe41__lane24_strm1_data_valid    ( std__pe41__lane24_strm1_data_valid ),      
               .std__pe41__lane24_strm1_data_mask     ( std__pe41__lane24_strm1_data_mask  ),      

               // PE 41, Lane 25                 
               .pe41__std__lane25_strm0_ready         ( pe41__std__lane25_strm0_ready      ),      
               .std__pe41__lane25_strm0_cntl          ( std__pe41__lane25_strm0_cntl       ),      
               .std__pe41__lane25_strm0_data          ( std__pe41__lane25_strm0_data       ),      
               .std__pe41__lane25_strm0_data_valid    ( std__pe41__lane25_strm0_data_valid ),      
               .std__pe41__lane25_strm0_data_mask     ( std__pe41__lane25_strm0_data_mask  ),      

               .pe41__std__lane25_strm1_ready         ( pe41__std__lane25_strm1_ready      ),      
               .std__pe41__lane25_strm1_cntl          ( std__pe41__lane25_strm1_cntl       ),      
               .std__pe41__lane25_strm1_data          ( std__pe41__lane25_strm1_data       ),      
               .std__pe41__lane25_strm1_data_valid    ( std__pe41__lane25_strm1_data_valid ),      
               .std__pe41__lane25_strm1_data_mask     ( std__pe41__lane25_strm1_data_mask  ),      

               // PE 41, Lane 26                 
               .pe41__std__lane26_strm0_ready         ( pe41__std__lane26_strm0_ready      ),      
               .std__pe41__lane26_strm0_cntl          ( std__pe41__lane26_strm0_cntl       ),      
               .std__pe41__lane26_strm0_data          ( std__pe41__lane26_strm0_data       ),      
               .std__pe41__lane26_strm0_data_valid    ( std__pe41__lane26_strm0_data_valid ),      
               .std__pe41__lane26_strm0_data_mask     ( std__pe41__lane26_strm0_data_mask  ),      

               .pe41__std__lane26_strm1_ready         ( pe41__std__lane26_strm1_ready      ),      
               .std__pe41__lane26_strm1_cntl          ( std__pe41__lane26_strm1_cntl       ),      
               .std__pe41__lane26_strm1_data          ( std__pe41__lane26_strm1_data       ),      
               .std__pe41__lane26_strm1_data_valid    ( std__pe41__lane26_strm1_data_valid ),      
               .std__pe41__lane26_strm1_data_mask     ( std__pe41__lane26_strm1_data_mask  ),      

               // PE 41, Lane 27                 
               .pe41__std__lane27_strm0_ready         ( pe41__std__lane27_strm0_ready      ),      
               .std__pe41__lane27_strm0_cntl          ( std__pe41__lane27_strm0_cntl       ),      
               .std__pe41__lane27_strm0_data          ( std__pe41__lane27_strm0_data       ),      
               .std__pe41__lane27_strm0_data_valid    ( std__pe41__lane27_strm0_data_valid ),      
               .std__pe41__lane27_strm0_data_mask     ( std__pe41__lane27_strm0_data_mask  ),      

               .pe41__std__lane27_strm1_ready         ( pe41__std__lane27_strm1_ready      ),      
               .std__pe41__lane27_strm1_cntl          ( std__pe41__lane27_strm1_cntl       ),      
               .std__pe41__lane27_strm1_data          ( std__pe41__lane27_strm1_data       ),      
               .std__pe41__lane27_strm1_data_valid    ( std__pe41__lane27_strm1_data_valid ),      
               .std__pe41__lane27_strm1_data_mask     ( std__pe41__lane27_strm1_data_mask  ),      

               // PE 41, Lane 28                 
               .pe41__std__lane28_strm0_ready         ( pe41__std__lane28_strm0_ready      ),      
               .std__pe41__lane28_strm0_cntl          ( std__pe41__lane28_strm0_cntl       ),      
               .std__pe41__lane28_strm0_data          ( std__pe41__lane28_strm0_data       ),      
               .std__pe41__lane28_strm0_data_valid    ( std__pe41__lane28_strm0_data_valid ),      
               .std__pe41__lane28_strm0_data_mask     ( std__pe41__lane28_strm0_data_mask  ),      

               .pe41__std__lane28_strm1_ready         ( pe41__std__lane28_strm1_ready      ),      
               .std__pe41__lane28_strm1_cntl          ( std__pe41__lane28_strm1_cntl       ),      
               .std__pe41__lane28_strm1_data          ( std__pe41__lane28_strm1_data       ),      
               .std__pe41__lane28_strm1_data_valid    ( std__pe41__lane28_strm1_data_valid ),      
               .std__pe41__lane28_strm1_data_mask     ( std__pe41__lane28_strm1_data_mask  ),      

               // PE 41, Lane 29                 
               .pe41__std__lane29_strm0_ready         ( pe41__std__lane29_strm0_ready      ),      
               .std__pe41__lane29_strm0_cntl          ( std__pe41__lane29_strm0_cntl       ),      
               .std__pe41__lane29_strm0_data          ( std__pe41__lane29_strm0_data       ),      
               .std__pe41__lane29_strm0_data_valid    ( std__pe41__lane29_strm0_data_valid ),      
               .std__pe41__lane29_strm0_data_mask     ( std__pe41__lane29_strm0_data_mask  ),      

               .pe41__std__lane29_strm1_ready         ( pe41__std__lane29_strm1_ready      ),      
               .std__pe41__lane29_strm1_cntl          ( std__pe41__lane29_strm1_cntl       ),      
               .std__pe41__lane29_strm1_data          ( std__pe41__lane29_strm1_data       ),      
               .std__pe41__lane29_strm1_data_valid    ( std__pe41__lane29_strm1_data_valid ),      
               .std__pe41__lane29_strm1_data_mask     ( std__pe41__lane29_strm1_data_mask  ),      

               // PE 41, Lane 30                 
               .pe41__std__lane30_strm0_ready         ( pe41__std__lane30_strm0_ready      ),      
               .std__pe41__lane30_strm0_cntl          ( std__pe41__lane30_strm0_cntl       ),      
               .std__pe41__lane30_strm0_data          ( std__pe41__lane30_strm0_data       ),      
               .std__pe41__lane30_strm0_data_valid    ( std__pe41__lane30_strm0_data_valid ),      
               .std__pe41__lane30_strm0_data_mask     ( std__pe41__lane30_strm0_data_mask  ),      

               .pe41__std__lane30_strm1_ready         ( pe41__std__lane30_strm1_ready      ),      
               .std__pe41__lane30_strm1_cntl          ( std__pe41__lane30_strm1_cntl       ),      
               .std__pe41__lane30_strm1_data          ( std__pe41__lane30_strm1_data       ),      
               .std__pe41__lane30_strm1_data_valid    ( std__pe41__lane30_strm1_data_valid ),      
               .std__pe41__lane30_strm1_data_mask     ( std__pe41__lane30_strm1_data_mask  ),      

               // PE 41, Lane 31                 
               .pe41__std__lane31_strm0_ready         ( pe41__std__lane31_strm0_ready      ),      
               .std__pe41__lane31_strm0_cntl          ( std__pe41__lane31_strm0_cntl       ),      
               .std__pe41__lane31_strm0_data          ( std__pe41__lane31_strm0_data       ),      
               .std__pe41__lane31_strm0_data_valid    ( std__pe41__lane31_strm0_data_valid ),      
               .std__pe41__lane31_strm0_data_mask     ( std__pe41__lane31_strm0_data_mask  ),      

               .pe41__std__lane31_strm1_ready         ( pe41__std__lane31_strm1_ready      ),      
               .std__pe41__lane31_strm1_cntl          ( std__pe41__lane31_strm1_cntl       ),      
               .std__pe41__lane31_strm1_data          ( std__pe41__lane31_strm1_data       ),      
               .std__pe41__lane31_strm1_data_valid    ( std__pe41__lane31_strm1_data_valid ),      
               .std__pe41__lane31_strm1_data_mask     ( std__pe41__lane31_strm1_data_mask  ),      

               // PE 42, Lane 0                 
               .pe42__std__lane0_strm0_ready         ( pe42__std__lane0_strm0_ready      ),      
               .std__pe42__lane0_strm0_cntl          ( std__pe42__lane0_strm0_cntl       ),      
               .std__pe42__lane0_strm0_data          ( std__pe42__lane0_strm0_data       ),      
               .std__pe42__lane0_strm0_data_valid    ( std__pe42__lane0_strm0_data_valid ),      
               .std__pe42__lane0_strm0_data_mask     ( std__pe42__lane0_strm0_data_mask  ),      

               .pe42__std__lane0_strm1_ready         ( pe42__std__lane0_strm1_ready      ),      
               .std__pe42__lane0_strm1_cntl          ( std__pe42__lane0_strm1_cntl       ),      
               .std__pe42__lane0_strm1_data          ( std__pe42__lane0_strm1_data       ),      
               .std__pe42__lane0_strm1_data_valid    ( std__pe42__lane0_strm1_data_valid ),      
               .std__pe42__lane0_strm1_data_mask     ( std__pe42__lane0_strm1_data_mask  ),      

               // PE 42, Lane 1                 
               .pe42__std__lane1_strm0_ready         ( pe42__std__lane1_strm0_ready      ),      
               .std__pe42__lane1_strm0_cntl          ( std__pe42__lane1_strm0_cntl       ),      
               .std__pe42__lane1_strm0_data          ( std__pe42__lane1_strm0_data       ),      
               .std__pe42__lane1_strm0_data_valid    ( std__pe42__lane1_strm0_data_valid ),      
               .std__pe42__lane1_strm0_data_mask     ( std__pe42__lane1_strm0_data_mask  ),      

               .pe42__std__lane1_strm1_ready         ( pe42__std__lane1_strm1_ready      ),      
               .std__pe42__lane1_strm1_cntl          ( std__pe42__lane1_strm1_cntl       ),      
               .std__pe42__lane1_strm1_data          ( std__pe42__lane1_strm1_data       ),      
               .std__pe42__lane1_strm1_data_valid    ( std__pe42__lane1_strm1_data_valid ),      
               .std__pe42__lane1_strm1_data_mask     ( std__pe42__lane1_strm1_data_mask  ),      

               // PE 42, Lane 2                 
               .pe42__std__lane2_strm0_ready         ( pe42__std__lane2_strm0_ready      ),      
               .std__pe42__lane2_strm0_cntl          ( std__pe42__lane2_strm0_cntl       ),      
               .std__pe42__lane2_strm0_data          ( std__pe42__lane2_strm0_data       ),      
               .std__pe42__lane2_strm0_data_valid    ( std__pe42__lane2_strm0_data_valid ),      
               .std__pe42__lane2_strm0_data_mask     ( std__pe42__lane2_strm0_data_mask  ),      

               .pe42__std__lane2_strm1_ready         ( pe42__std__lane2_strm1_ready      ),      
               .std__pe42__lane2_strm1_cntl          ( std__pe42__lane2_strm1_cntl       ),      
               .std__pe42__lane2_strm1_data          ( std__pe42__lane2_strm1_data       ),      
               .std__pe42__lane2_strm1_data_valid    ( std__pe42__lane2_strm1_data_valid ),      
               .std__pe42__lane2_strm1_data_mask     ( std__pe42__lane2_strm1_data_mask  ),      

               // PE 42, Lane 3                 
               .pe42__std__lane3_strm0_ready         ( pe42__std__lane3_strm0_ready      ),      
               .std__pe42__lane3_strm0_cntl          ( std__pe42__lane3_strm0_cntl       ),      
               .std__pe42__lane3_strm0_data          ( std__pe42__lane3_strm0_data       ),      
               .std__pe42__lane3_strm0_data_valid    ( std__pe42__lane3_strm0_data_valid ),      
               .std__pe42__lane3_strm0_data_mask     ( std__pe42__lane3_strm0_data_mask  ),      

               .pe42__std__lane3_strm1_ready         ( pe42__std__lane3_strm1_ready      ),      
               .std__pe42__lane3_strm1_cntl          ( std__pe42__lane3_strm1_cntl       ),      
               .std__pe42__lane3_strm1_data          ( std__pe42__lane3_strm1_data       ),      
               .std__pe42__lane3_strm1_data_valid    ( std__pe42__lane3_strm1_data_valid ),      
               .std__pe42__lane3_strm1_data_mask     ( std__pe42__lane3_strm1_data_mask  ),      

               // PE 42, Lane 4                 
               .pe42__std__lane4_strm0_ready         ( pe42__std__lane4_strm0_ready      ),      
               .std__pe42__lane4_strm0_cntl          ( std__pe42__lane4_strm0_cntl       ),      
               .std__pe42__lane4_strm0_data          ( std__pe42__lane4_strm0_data       ),      
               .std__pe42__lane4_strm0_data_valid    ( std__pe42__lane4_strm0_data_valid ),      
               .std__pe42__lane4_strm0_data_mask     ( std__pe42__lane4_strm0_data_mask  ),      

               .pe42__std__lane4_strm1_ready         ( pe42__std__lane4_strm1_ready      ),      
               .std__pe42__lane4_strm1_cntl          ( std__pe42__lane4_strm1_cntl       ),      
               .std__pe42__lane4_strm1_data          ( std__pe42__lane4_strm1_data       ),      
               .std__pe42__lane4_strm1_data_valid    ( std__pe42__lane4_strm1_data_valid ),      
               .std__pe42__lane4_strm1_data_mask     ( std__pe42__lane4_strm1_data_mask  ),      

               // PE 42, Lane 5                 
               .pe42__std__lane5_strm0_ready         ( pe42__std__lane5_strm0_ready      ),      
               .std__pe42__lane5_strm0_cntl          ( std__pe42__lane5_strm0_cntl       ),      
               .std__pe42__lane5_strm0_data          ( std__pe42__lane5_strm0_data       ),      
               .std__pe42__lane5_strm0_data_valid    ( std__pe42__lane5_strm0_data_valid ),      
               .std__pe42__lane5_strm0_data_mask     ( std__pe42__lane5_strm0_data_mask  ),      

               .pe42__std__lane5_strm1_ready         ( pe42__std__lane5_strm1_ready      ),      
               .std__pe42__lane5_strm1_cntl          ( std__pe42__lane5_strm1_cntl       ),      
               .std__pe42__lane5_strm1_data          ( std__pe42__lane5_strm1_data       ),      
               .std__pe42__lane5_strm1_data_valid    ( std__pe42__lane5_strm1_data_valid ),      
               .std__pe42__lane5_strm1_data_mask     ( std__pe42__lane5_strm1_data_mask  ),      

               // PE 42, Lane 6                 
               .pe42__std__lane6_strm0_ready         ( pe42__std__lane6_strm0_ready      ),      
               .std__pe42__lane6_strm0_cntl          ( std__pe42__lane6_strm0_cntl       ),      
               .std__pe42__lane6_strm0_data          ( std__pe42__lane6_strm0_data       ),      
               .std__pe42__lane6_strm0_data_valid    ( std__pe42__lane6_strm0_data_valid ),      
               .std__pe42__lane6_strm0_data_mask     ( std__pe42__lane6_strm0_data_mask  ),      

               .pe42__std__lane6_strm1_ready         ( pe42__std__lane6_strm1_ready      ),      
               .std__pe42__lane6_strm1_cntl          ( std__pe42__lane6_strm1_cntl       ),      
               .std__pe42__lane6_strm1_data          ( std__pe42__lane6_strm1_data       ),      
               .std__pe42__lane6_strm1_data_valid    ( std__pe42__lane6_strm1_data_valid ),      
               .std__pe42__lane6_strm1_data_mask     ( std__pe42__lane6_strm1_data_mask  ),      

               // PE 42, Lane 7                 
               .pe42__std__lane7_strm0_ready         ( pe42__std__lane7_strm0_ready      ),      
               .std__pe42__lane7_strm0_cntl          ( std__pe42__lane7_strm0_cntl       ),      
               .std__pe42__lane7_strm0_data          ( std__pe42__lane7_strm0_data       ),      
               .std__pe42__lane7_strm0_data_valid    ( std__pe42__lane7_strm0_data_valid ),      
               .std__pe42__lane7_strm0_data_mask     ( std__pe42__lane7_strm0_data_mask  ),      

               .pe42__std__lane7_strm1_ready         ( pe42__std__lane7_strm1_ready      ),      
               .std__pe42__lane7_strm1_cntl          ( std__pe42__lane7_strm1_cntl       ),      
               .std__pe42__lane7_strm1_data          ( std__pe42__lane7_strm1_data       ),      
               .std__pe42__lane7_strm1_data_valid    ( std__pe42__lane7_strm1_data_valid ),      
               .std__pe42__lane7_strm1_data_mask     ( std__pe42__lane7_strm1_data_mask  ),      

               // PE 42, Lane 8                 
               .pe42__std__lane8_strm0_ready         ( pe42__std__lane8_strm0_ready      ),      
               .std__pe42__lane8_strm0_cntl          ( std__pe42__lane8_strm0_cntl       ),      
               .std__pe42__lane8_strm0_data          ( std__pe42__lane8_strm0_data       ),      
               .std__pe42__lane8_strm0_data_valid    ( std__pe42__lane8_strm0_data_valid ),      
               .std__pe42__lane8_strm0_data_mask     ( std__pe42__lane8_strm0_data_mask  ),      

               .pe42__std__lane8_strm1_ready         ( pe42__std__lane8_strm1_ready      ),      
               .std__pe42__lane8_strm1_cntl          ( std__pe42__lane8_strm1_cntl       ),      
               .std__pe42__lane8_strm1_data          ( std__pe42__lane8_strm1_data       ),      
               .std__pe42__lane8_strm1_data_valid    ( std__pe42__lane8_strm1_data_valid ),      
               .std__pe42__lane8_strm1_data_mask     ( std__pe42__lane8_strm1_data_mask  ),      

               // PE 42, Lane 9                 
               .pe42__std__lane9_strm0_ready         ( pe42__std__lane9_strm0_ready      ),      
               .std__pe42__lane9_strm0_cntl          ( std__pe42__lane9_strm0_cntl       ),      
               .std__pe42__lane9_strm0_data          ( std__pe42__lane9_strm0_data       ),      
               .std__pe42__lane9_strm0_data_valid    ( std__pe42__lane9_strm0_data_valid ),      
               .std__pe42__lane9_strm0_data_mask     ( std__pe42__lane9_strm0_data_mask  ),      

               .pe42__std__lane9_strm1_ready         ( pe42__std__lane9_strm1_ready      ),      
               .std__pe42__lane9_strm1_cntl          ( std__pe42__lane9_strm1_cntl       ),      
               .std__pe42__lane9_strm1_data          ( std__pe42__lane9_strm1_data       ),      
               .std__pe42__lane9_strm1_data_valid    ( std__pe42__lane9_strm1_data_valid ),      
               .std__pe42__lane9_strm1_data_mask     ( std__pe42__lane9_strm1_data_mask  ),      

               // PE 42, Lane 10                 
               .pe42__std__lane10_strm0_ready         ( pe42__std__lane10_strm0_ready      ),      
               .std__pe42__lane10_strm0_cntl          ( std__pe42__lane10_strm0_cntl       ),      
               .std__pe42__lane10_strm0_data          ( std__pe42__lane10_strm0_data       ),      
               .std__pe42__lane10_strm0_data_valid    ( std__pe42__lane10_strm0_data_valid ),      
               .std__pe42__lane10_strm0_data_mask     ( std__pe42__lane10_strm0_data_mask  ),      

               .pe42__std__lane10_strm1_ready         ( pe42__std__lane10_strm1_ready      ),      
               .std__pe42__lane10_strm1_cntl          ( std__pe42__lane10_strm1_cntl       ),      
               .std__pe42__lane10_strm1_data          ( std__pe42__lane10_strm1_data       ),      
               .std__pe42__lane10_strm1_data_valid    ( std__pe42__lane10_strm1_data_valid ),      
               .std__pe42__lane10_strm1_data_mask     ( std__pe42__lane10_strm1_data_mask  ),      

               // PE 42, Lane 11                 
               .pe42__std__lane11_strm0_ready         ( pe42__std__lane11_strm0_ready      ),      
               .std__pe42__lane11_strm0_cntl          ( std__pe42__lane11_strm0_cntl       ),      
               .std__pe42__lane11_strm0_data          ( std__pe42__lane11_strm0_data       ),      
               .std__pe42__lane11_strm0_data_valid    ( std__pe42__lane11_strm0_data_valid ),      
               .std__pe42__lane11_strm0_data_mask     ( std__pe42__lane11_strm0_data_mask  ),      

               .pe42__std__lane11_strm1_ready         ( pe42__std__lane11_strm1_ready      ),      
               .std__pe42__lane11_strm1_cntl          ( std__pe42__lane11_strm1_cntl       ),      
               .std__pe42__lane11_strm1_data          ( std__pe42__lane11_strm1_data       ),      
               .std__pe42__lane11_strm1_data_valid    ( std__pe42__lane11_strm1_data_valid ),      
               .std__pe42__lane11_strm1_data_mask     ( std__pe42__lane11_strm1_data_mask  ),      

               // PE 42, Lane 12                 
               .pe42__std__lane12_strm0_ready         ( pe42__std__lane12_strm0_ready      ),      
               .std__pe42__lane12_strm0_cntl          ( std__pe42__lane12_strm0_cntl       ),      
               .std__pe42__lane12_strm0_data          ( std__pe42__lane12_strm0_data       ),      
               .std__pe42__lane12_strm0_data_valid    ( std__pe42__lane12_strm0_data_valid ),      
               .std__pe42__lane12_strm0_data_mask     ( std__pe42__lane12_strm0_data_mask  ),      

               .pe42__std__lane12_strm1_ready         ( pe42__std__lane12_strm1_ready      ),      
               .std__pe42__lane12_strm1_cntl          ( std__pe42__lane12_strm1_cntl       ),      
               .std__pe42__lane12_strm1_data          ( std__pe42__lane12_strm1_data       ),      
               .std__pe42__lane12_strm1_data_valid    ( std__pe42__lane12_strm1_data_valid ),      
               .std__pe42__lane12_strm1_data_mask     ( std__pe42__lane12_strm1_data_mask  ),      

               // PE 42, Lane 13                 
               .pe42__std__lane13_strm0_ready         ( pe42__std__lane13_strm0_ready      ),      
               .std__pe42__lane13_strm0_cntl          ( std__pe42__lane13_strm0_cntl       ),      
               .std__pe42__lane13_strm0_data          ( std__pe42__lane13_strm0_data       ),      
               .std__pe42__lane13_strm0_data_valid    ( std__pe42__lane13_strm0_data_valid ),      
               .std__pe42__lane13_strm0_data_mask     ( std__pe42__lane13_strm0_data_mask  ),      

               .pe42__std__lane13_strm1_ready         ( pe42__std__lane13_strm1_ready      ),      
               .std__pe42__lane13_strm1_cntl          ( std__pe42__lane13_strm1_cntl       ),      
               .std__pe42__lane13_strm1_data          ( std__pe42__lane13_strm1_data       ),      
               .std__pe42__lane13_strm1_data_valid    ( std__pe42__lane13_strm1_data_valid ),      
               .std__pe42__lane13_strm1_data_mask     ( std__pe42__lane13_strm1_data_mask  ),      

               // PE 42, Lane 14                 
               .pe42__std__lane14_strm0_ready         ( pe42__std__lane14_strm0_ready      ),      
               .std__pe42__lane14_strm0_cntl          ( std__pe42__lane14_strm0_cntl       ),      
               .std__pe42__lane14_strm0_data          ( std__pe42__lane14_strm0_data       ),      
               .std__pe42__lane14_strm0_data_valid    ( std__pe42__lane14_strm0_data_valid ),      
               .std__pe42__lane14_strm0_data_mask     ( std__pe42__lane14_strm0_data_mask  ),      

               .pe42__std__lane14_strm1_ready         ( pe42__std__lane14_strm1_ready      ),      
               .std__pe42__lane14_strm1_cntl          ( std__pe42__lane14_strm1_cntl       ),      
               .std__pe42__lane14_strm1_data          ( std__pe42__lane14_strm1_data       ),      
               .std__pe42__lane14_strm1_data_valid    ( std__pe42__lane14_strm1_data_valid ),      
               .std__pe42__lane14_strm1_data_mask     ( std__pe42__lane14_strm1_data_mask  ),      

               // PE 42, Lane 15                 
               .pe42__std__lane15_strm0_ready         ( pe42__std__lane15_strm0_ready      ),      
               .std__pe42__lane15_strm0_cntl          ( std__pe42__lane15_strm0_cntl       ),      
               .std__pe42__lane15_strm0_data          ( std__pe42__lane15_strm0_data       ),      
               .std__pe42__lane15_strm0_data_valid    ( std__pe42__lane15_strm0_data_valid ),      
               .std__pe42__lane15_strm0_data_mask     ( std__pe42__lane15_strm0_data_mask  ),      

               .pe42__std__lane15_strm1_ready         ( pe42__std__lane15_strm1_ready      ),      
               .std__pe42__lane15_strm1_cntl          ( std__pe42__lane15_strm1_cntl       ),      
               .std__pe42__lane15_strm1_data          ( std__pe42__lane15_strm1_data       ),      
               .std__pe42__lane15_strm1_data_valid    ( std__pe42__lane15_strm1_data_valid ),      
               .std__pe42__lane15_strm1_data_mask     ( std__pe42__lane15_strm1_data_mask  ),      

               // PE 42, Lane 16                 
               .pe42__std__lane16_strm0_ready         ( pe42__std__lane16_strm0_ready      ),      
               .std__pe42__lane16_strm0_cntl          ( std__pe42__lane16_strm0_cntl       ),      
               .std__pe42__lane16_strm0_data          ( std__pe42__lane16_strm0_data       ),      
               .std__pe42__lane16_strm0_data_valid    ( std__pe42__lane16_strm0_data_valid ),      
               .std__pe42__lane16_strm0_data_mask     ( std__pe42__lane16_strm0_data_mask  ),      

               .pe42__std__lane16_strm1_ready         ( pe42__std__lane16_strm1_ready      ),      
               .std__pe42__lane16_strm1_cntl          ( std__pe42__lane16_strm1_cntl       ),      
               .std__pe42__lane16_strm1_data          ( std__pe42__lane16_strm1_data       ),      
               .std__pe42__lane16_strm1_data_valid    ( std__pe42__lane16_strm1_data_valid ),      
               .std__pe42__lane16_strm1_data_mask     ( std__pe42__lane16_strm1_data_mask  ),      

               // PE 42, Lane 17                 
               .pe42__std__lane17_strm0_ready         ( pe42__std__lane17_strm0_ready      ),      
               .std__pe42__lane17_strm0_cntl          ( std__pe42__lane17_strm0_cntl       ),      
               .std__pe42__lane17_strm0_data          ( std__pe42__lane17_strm0_data       ),      
               .std__pe42__lane17_strm0_data_valid    ( std__pe42__lane17_strm0_data_valid ),      
               .std__pe42__lane17_strm0_data_mask     ( std__pe42__lane17_strm0_data_mask  ),      

               .pe42__std__lane17_strm1_ready         ( pe42__std__lane17_strm1_ready      ),      
               .std__pe42__lane17_strm1_cntl          ( std__pe42__lane17_strm1_cntl       ),      
               .std__pe42__lane17_strm1_data          ( std__pe42__lane17_strm1_data       ),      
               .std__pe42__lane17_strm1_data_valid    ( std__pe42__lane17_strm1_data_valid ),      
               .std__pe42__lane17_strm1_data_mask     ( std__pe42__lane17_strm1_data_mask  ),      

               // PE 42, Lane 18                 
               .pe42__std__lane18_strm0_ready         ( pe42__std__lane18_strm0_ready      ),      
               .std__pe42__lane18_strm0_cntl          ( std__pe42__lane18_strm0_cntl       ),      
               .std__pe42__lane18_strm0_data          ( std__pe42__lane18_strm0_data       ),      
               .std__pe42__lane18_strm0_data_valid    ( std__pe42__lane18_strm0_data_valid ),      
               .std__pe42__lane18_strm0_data_mask     ( std__pe42__lane18_strm0_data_mask  ),      

               .pe42__std__lane18_strm1_ready         ( pe42__std__lane18_strm1_ready      ),      
               .std__pe42__lane18_strm1_cntl          ( std__pe42__lane18_strm1_cntl       ),      
               .std__pe42__lane18_strm1_data          ( std__pe42__lane18_strm1_data       ),      
               .std__pe42__lane18_strm1_data_valid    ( std__pe42__lane18_strm1_data_valid ),      
               .std__pe42__lane18_strm1_data_mask     ( std__pe42__lane18_strm1_data_mask  ),      

               // PE 42, Lane 19                 
               .pe42__std__lane19_strm0_ready         ( pe42__std__lane19_strm0_ready      ),      
               .std__pe42__lane19_strm0_cntl          ( std__pe42__lane19_strm0_cntl       ),      
               .std__pe42__lane19_strm0_data          ( std__pe42__lane19_strm0_data       ),      
               .std__pe42__lane19_strm0_data_valid    ( std__pe42__lane19_strm0_data_valid ),      
               .std__pe42__lane19_strm0_data_mask     ( std__pe42__lane19_strm0_data_mask  ),      

               .pe42__std__lane19_strm1_ready         ( pe42__std__lane19_strm1_ready      ),      
               .std__pe42__lane19_strm1_cntl          ( std__pe42__lane19_strm1_cntl       ),      
               .std__pe42__lane19_strm1_data          ( std__pe42__lane19_strm1_data       ),      
               .std__pe42__lane19_strm1_data_valid    ( std__pe42__lane19_strm1_data_valid ),      
               .std__pe42__lane19_strm1_data_mask     ( std__pe42__lane19_strm1_data_mask  ),      

               // PE 42, Lane 20                 
               .pe42__std__lane20_strm0_ready         ( pe42__std__lane20_strm0_ready      ),      
               .std__pe42__lane20_strm0_cntl          ( std__pe42__lane20_strm0_cntl       ),      
               .std__pe42__lane20_strm0_data          ( std__pe42__lane20_strm0_data       ),      
               .std__pe42__lane20_strm0_data_valid    ( std__pe42__lane20_strm0_data_valid ),      
               .std__pe42__lane20_strm0_data_mask     ( std__pe42__lane20_strm0_data_mask  ),      

               .pe42__std__lane20_strm1_ready         ( pe42__std__lane20_strm1_ready      ),      
               .std__pe42__lane20_strm1_cntl          ( std__pe42__lane20_strm1_cntl       ),      
               .std__pe42__lane20_strm1_data          ( std__pe42__lane20_strm1_data       ),      
               .std__pe42__lane20_strm1_data_valid    ( std__pe42__lane20_strm1_data_valid ),      
               .std__pe42__lane20_strm1_data_mask     ( std__pe42__lane20_strm1_data_mask  ),      

               // PE 42, Lane 21                 
               .pe42__std__lane21_strm0_ready         ( pe42__std__lane21_strm0_ready      ),      
               .std__pe42__lane21_strm0_cntl          ( std__pe42__lane21_strm0_cntl       ),      
               .std__pe42__lane21_strm0_data          ( std__pe42__lane21_strm0_data       ),      
               .std__pe42__lane21_strm0_data_valid    ( std__pe42__lane21_strm0_data_valid ),      
               .std__pe42__lane21_strm0_data_mask     ( std__pe42__lane21_strm0_data_mask  ),      

               .pe42__std__lane21_strm1_ready         ( pe42__std__lane21_strm1_ready      ),      
               .std__pe42__lane21_strm1_cntl          ( std__pe42__lane21_strm1_cntl       ),      
               .std__pe42__lane21_strm1_data          ( std__pe42__lane21_strm1_data       ),      
               .std__pe42__lane21_strm1_data_valid    ( std__pe42__lane21_strm1_data_valid ),      
               .std__pe42__lane21_strm1_data_mask     ( std__pe42__lane21_strm1_data_mask  ),      

               // PE 42, Lane 22                 
               .pe42__std__lane22_strm0_ready         ( pe42__std__lane22_strm0_ready      ),      
               .std__pe42__lane22_strm0_cntl          ( std__pe42__lane22_strm0_cntl       ),      
               .std__pe42__lane22_strm0_data          ( std__pe42__lane22_strm0_data       ),      
               .std__pe42__lane22_strm0_data_valid    ( std__pe42__lane22_strm0_data_valid ),      
               .std__pe42__lane22_strm0_data_mask     ( std__pe42__lane22_strm0_data_mask  ),      

               .pe42__std__lane22_strm1_ready         ( pe42__std__lane22_strm1_ready      ),      
               .std__pe42__lane22_strm1_cntl          ( std__pe42__lane22_strm1_cntl       ),      
               .std__pe42__lane22_strm1_data          ( std__pe42__lane22_strm1_data       ),      
               .std__pe42__lane22_strm1_data_valid    ( std__pe42__lane22_strm1_data_valid ),      
               .std__pe42__lane22_strm1_data_mask     ( std__pe42__lane22_strm1_data_mask  ),      

               // PE 42, Lane 23                 
               .pe42__std__lane23_strm0_ready         ( pe42__std__lane23_strm0_ready      ),      
               .std__pe42__lane23_strm0_cntl          ( std__pe42__lane23_strm0_cntl       ),      
               .std__pe42__lane23_strm0_data          ( std__pe42__lane23_strm0_data       ),      
               .std__pe42__lane23_strm0_data_valid    ( std__pe42__lane23_strm0_data_valid ),      
               .std__pe42__lane23_strm0_data_mask     ( std__pe42__lane23_strm0_data_mask  ),      

               .pe42__std__lane23_strm1_ready         ( pe42__std__lane23_strm1_ready      ),      
               .std__pe42__lane23_strm1_cntl          ( std__pe42__lane23_strm1_cntl       ),      
               .std__pe42__lane23_strm1_data          ( std__pe42__lane23_strm1_data       ),      
               .std__pe42__lane23_strm1_data_valid    ( std__pe42__lane23_strm1_data_valid ),      
               .std__pe42__lane23_strm1_data_mask     ( std__pe42__lane23_strm1_data_mask  ),      

               // PE 42, Lane 24                 
               .pe42__std__lane24_strm0_ready         ( pe42__std__lane24_strm0_ready      ),      
               .std__pe42__lane24_strm0_cntl          ( std__pe42__lane24_strm0_cntl       ),      
               .std__pe42__lane24_strm0_data          ( std__pe42__lane24_strm0_data       ),      
               .std__pe42__lane24_strm0_data_valid    ( std__pe42__lane24_strm0_data_valid ),      
               .std__pe42__lane24_strm0_data_mask     ( std__pe42__lane24_strm0_data_mask  ),      

               .pe42__std__lane24_strm1_ready         ( pe42__std__lane24_strm1_ready      ),      
               .std__pe42__lane24_strm1_cntl          ( std__pe42__lane24_strm1_cntl       ),      
               .std__pe42__lane24_strm1_data          ( std__pe42__lane24_strm1_data       ),      
               .std__pe42__lane24_strm1_data_valid    ( std__pe42__lane24_strm1_data_valid ),      
               .std__pe42__lane24_strm1_data_mask     ( std__pe42__lane24_strm1_data_mask  ),      

               // PE 42, Lane 25                 
               .pe42__std__lane25_strm0_ready         ( pe42__std__lane25_strm0_ready      ),      
               .std__pe42__lane25_strm0_cntl          ( std__pe42__lane25_strm0_cntl       ),      
               .std__pe42__lane25_strm0_data          ( std__pe42__lane25_strm0_data       ),      
               .std__pe42__lane25_strm0_data_valid    ( std__pe42__lane25_strm0_data_valid ),      
               .std__pe42__lane25_strm0_data_mask     ( std__pe42__lane25_strm0_data_mask  ),      

               .pe42__std__lane25_strm1_ready         ( pe42__std__lane25_strm1_ready      ),      
               .std__pe42__lane25_strm1_cntl          ( std__pe42__lane25_strm1_cntl       ),      
               .std__pe42__lane25_strm1_data          ( std__pe42__lane25_strm1_data       ),      
               .std__pe42__lane25_strm1_data_valid    ( std__pe42__lane25_strm1_data_valid ),      
               .std__pe42__lane25_strm1_data_mask     ( std__pe42__lane25_strm1_data_mask  ),      

               // PE 42, Lane 26                 
               .pe42__std__lane26_strm0_ready         ( pe42__std__lane26_strm0_ready      ),      
               .std__pe42__lane26_strm0_cntl          ( std__pe42__lane26_strm0_cntl       ),      
               .std__pe42__lane26_strm0_data          ( std__pe42__lane26_strm0_data       ),      
               .std__pe42__lane26_strm0_data_valid    ( std__pe42__lane26_strm0_data_valid ),      
               .std__pe42__lane26_strm0_data_mask     ( std__pe42__lane26_strm0_data_mask  ),      

               .pe42__std__lane26_strm1_ready         ( pe42__std__lane26_strm1_ready      ),      
               .std__pe42__lane26_strm1_cntl          ( std__pe42__lane26_strm1_cntl       ),      
               .std__pe42__lane26_strm1_data          ( std__pe42__lane26_strm1_data       ),      
               .std__pe42__lane26_strm1_data_valid    ( std__pe42__lane26_strm1_data_valid ),      
               .std__pe42__lane26_strm1_data_mask     ( std__pe42__lane26_strm1_data_mask  ),      

               // PE 42, Lane 27                 
               .pe42__std__lane27_strm0_ready         ( pe42__std__lane27_strm0_ready      ),      
               .std__pe42__lane27_strm0_cntl          ( std__pe42__lane27_strm0_cntl       ),      
               .std__pe42__lane27_strm0_data          ( std__pe42__lane27_strm0_data       ),      
               .std__pe42__lane27_strm0_data_valid    ( std__pe42__lane27_strm0_data_valid ),      
               .std__pe42__lane27_strm0_data_mask     ( std__pe42__lane27_strm0_data_mask  ),      

               .pe42__std__lane27_strm1_ready         ( pe42__std__lane27_strm1_ready      ),      
               .std__pe42__lane27_strm1_cntl          ( std__pe42__lane27_strm1_cntl       ),      
               .std__pe42__lane27_strm1_data          ( std__pe42__lane27_strm1_data       ),      
               .std__pe42__lane27_strm1_data_valid    ( std__pe42__lane27_strm1_data_valid ),      
               .std__pe42__lane27_strm1_data_mask     ( std__pe42__lane27_strm1_data_mask  ),      

               // PE 42, Lane 28                 
               .pe42__std__lane28_strm0_ready         ( pe42__std__lane28_strm0_ready      ),      
               .std__pe42__lane28_strm0_cntl          ( std__pe42__lane28_strm0_cntl       ),      
               .std__pe42__lane28_strm0_data          ( std__pe42__lane28_strm0_data       ),      
               .std__pe42__lane28_strm0_data_valid    ( std__pe42__lane28_strm0_data_valid ),      
               .std__pe42__lane28_strm0_data_mask     ( std__pe42__lane28_strm0_data_mask  ),      

               .pe42__std__lane28_strm1_ready         ( pe42__std__lane28_strm1_ready      ),      
               .std__pe42__lane28_strm1_cntl          ( std__pe42__lane28_strm1_cntl       ),      
               .std__pe42__lane28_strm1_data          ( std__pe42__lane28_strm1_data       ),      
               .std__pe42__lane28_strm1_data_valid    ( std__pe42__lane28_strm1_data_valid ),      
               .std__pe42__lane28_strm1_data_mask     ( std__pe42__lane28_strm1_data_mask  ),      

               // PE 42, Lane 29                 
               .pe42__std__lane29_strm0_ready         ( pe42__std__lane29_strm0_ready      ),      
               .std__pe42__lane29_strm0_cntl          ( std__pe42__lane29_strm0_cntl       ),      
               .std__pe42__lane29_strm0_data          ( std__pe42__lane29_strm0_data       ),      
               .std__pe42__lane29_strm0_data_valid    ( std__pe42__lane29_strm0_data_valid ),      
               .std__pe42__lane29_strm0_data_mask     ( std__pe42__lane29_strm0_data_mask  ),      

               .pe42__std__lane29_strm1_ready         ( pe42__std__lane29_strm1_ready      ),      
               .std__pe42__lane29_strm1_cntl          ( std__pe42__lane29_strm1_cntl       ),      
               .std__pe42__lane29_strm1_data          ( std__pe42__lane29_strm1_data       ),      
               .std__pe42__lane29_strm1_data_valid    ( std__pe42__lane29_strm1_data_valid ),      
               .std__pe42__lane29_strm1_data_mask     ( std__pe42__lane29_strm1_data_mask  ),      

               // PE 42, Lane 30                 
               .pe42__std__lane30_strm0_ready         ( pe42__std__lane30_strm0_ready      ),      
               .std__pe42__lane30_strm0_cntl          ( std__pe42__lane30_strm0_cntl       ),      
               .std__pe42__lane30_strm0_data          ( std__pe42__lane30_strm0_data       ),      
               .std__pe42__lane30_strm0_data_valid    ( std__pe42__lane30_strm0_data_valid ),      
               .std__pe42__lane30_strm0_data_mask     ( std__pe42__lane30_strm0_data_mask  ),      

               .pe42__std__lane30_strm1_ready         ( pe42__std__lane30_strm1_ready      ),      
               .std__pe42__lane30_strm1_cntl          ( std__pe42__lane30_strm1_cntl       ),      
               .std__pe42__lane30_strm1_data          ( std__pe42__lane30_strm1_data       ),      
               .std__pe42__lane30_strm1_data_valid    ( std__pe42__lane30_strm1_data_valid ),      
               .std__pe42__lane30_strm1_data_mask     ( std__pe42__lane30_strm1_data_mask  ),      

               // PE 42, Lane 31                 
               .pe42__std__lane31_strm0_ready         ( pe42__std__lane31_strm0_ready      ),      
               .std__pe42__lane31_strm0_cntl          ( std__pe42__lane31_strm0_cntl       ),      
               .std__pe42__lane31_strm0_data          ( std__pe42__lane31_strm0_data       ),      
               .std__pe42__lane31_strm0_data_valid    ( std__pe42__lane31_strm0_data_valid ),      
               .std__pe42__lane31_strm0_data_mask     ( std__pe42__lane31_strm0_data_mask  ),      

               .pe42__std__lane31_strm1_ready         ( pe42__std__lane31_strm1_ready      ),      
               .std__pe42__lane31_strm1_cntl          ( std__pe42__lane31_strm1_cntl       ),      
               .std__pe42__lane31_strm1_data          ( std__pe42__lane31_strm1_data       ),      
               .std__pe42__lane31_strm1_data_valid    ( std__pe42__lane31_strm1_data_valid ),      
               .std__pe42__lane31_strm1_data_mask     ( std__pe42__lane31_strm1_data_mask  ),      

               // PE 43, Lane 0                 
               .pe43__std__lane0_strm0_ready         ( pe43__std__lane0_strm0_ready      ),      
               .std__pe43__lane0_strm0_cntl          ( std__pe43__lane0_strm0_cntl       ),      
               .std__pe43__lane0_strm0_data          ( std__pe43__lane0_strm0_data       ),      
               .std__pe43__lane0_strm0_data_valid    ( std__pe43__lane0_strm0_data_valid ),      
               .std__pe43__lane0_strm0_data_mask     ( std__pe43__lane0_strm0_data_mask  ),      

               .pe43__std__lane0_strm1_ready         ( pe43__std__lane0_strm1_ready      ),      
               .std__pe43__lane0_strm1_cntl          ( std__pe43__lane0_strm1_cntl       ),      
               .std__pe43__lane0_strm1_data          ( std__pe43__lane0_strm1_data       ),      
               .std__pe43__lane0_strm1_data_valid    ( std__pe43__lane0_strm1_data_valid ),      
               .std__pe43__lane0_strm1_data_mask     ( std__pe43__lane0_strm1_data_mask  ),      

               // PE 43, Lane 1                 
               .pe43__std__lane1_strm0_ready         ( pe43__std__lane1_strm0_ready      ),      
               .std__pe43__lane1_strm0_cntl          ( std__pe43__lane1_strm0_cntl       ),      
               .std__pe43__lane1_strm0_data          ( std__pe43__lane1_strm0_data       ),      
               .std__pe43__lane1_strm0_data_valid    ( std__pe43__lane1_strm0_data_valid ),      
               .std__pe43__lane1_strm0_data_mask     ( std__pe43__lane1_strm0_data_mask  ),      

               .pe43__std__lane1_strm1_ready         ( pe43__std__lane1_strm1_ready      ),      
               .std__pe43__lane1_strm1_cntl          ( std__pe43__lane1_strm1_cntl       ),      
               .std__pe43__lane1_strm1_data          ( std__pe43__lane1_strm1_data       ),      
               .std__pe43__lane1_strm1_data_valid    ( std__pe43__lane1_strm1_data_valid ),      
               .std__pe43__lane1_strm1_data_mask     ( std__pe43__lane1_strm1_data_mask  ),      

               // PE 43, Lane 2                 
               .pe43__std__lane2_strm0_ready         ( pe43__std__lane2_strm0_ready      ),      
               .std__pe43__lane2_strm0_cntl          ( std__pe43__lane2_strm0_cntl       ),      
               .std__pe43__lane2_strm0_data          ( std__pe43__lane2_strm0_data       ),      
               .std__pe43__lane2_strm0_data_valid    ( std__pe43__lane2_strm0_data_valid ),      
               .std__pe43__lane2_strm0_data_mask     ( std__pe43__lane2_strm0_data_mask  ),      

               .pe43__std__lane2_strm1_ready         ( pe43__std__lane2_strm1_ready      ),      
               .std__pe43__lane2_strm1_cntl          ( std__pe43__lane2_strm1_cntl       ),      
               .std__pe43__lane2_strm1_data          ( std__pe43__lane2_strm1_data       ),      
               .std__pe43__lane2_strm1_data_valid    ( std__pe43__lane2_strm1_data_valid ),      
               .std__pe43__lane2_strm1_data_mask     ( std__pe43__lane2_strm1_data_mask  ),      

               // PE 43, Lane 3                 
               .pe43__std__lane3_strm0_ready         ( pe43__std__lane3_strm0_ready      ),      
               .std__pe43__lane3_strm0_cntl          ( std__pe43__lane3_strm0_cntl       ),      
               .std__pe43__lane3_strm0_data          ( std__pe43__lane3_strm0_data       ),      
               .std__pe43__lane3_strm0_data_valid    ( std__pe43__lane3_strm0_data_valid ),      
               .std__pe43__lane3_strm0_data_mask     ( std__pe43__lane3_strm0_data_mask  ),      

               .pe43__std__lane3_strm1_ready         ( pe43__std__lane3_strm1_ready      ),      
               .std__pe43__lane3_strm1_cntl          ( std__pe43__lane3_strm1_cntl       ),      
               .std__pe43__lane3_strm1_data          ( std__pe43__lane3_strm1_data       ),      
               .std__pe43__lane3_strm1_data_valid    ( std__pe43__lane3_strm1_data_valid ),      
               .std__pe43__lane3_strm1_data_mask     ( std__pe43__lane3_strm1_data_mask  ),      

               // PE 43, Lane 4                 
               .pe43__std__lane4_strm0_ready         ( pe43__std__lane4_strm0_ready      ),      
               .std__pe43__lane4_strm0_cntl          ( std__pe43__lane4_strm0_cntl       ),      
               .std__pe43__lane4_strm0_data          ( std__pe43__lane4_strm0_data       ),      
               .std__pe43__lane4_strm0_data_valid    ( std__pe43__lane4_strm0_data_valid ),      
               .std__pe43__lane4_strm0_data_mask     ( std__pe43__lane4_strm0_data_mask  ),      

               .pe43__std__lane4_strm1_ready         ( pe43__std__lane4_strm1_ready      ),      
               .std__pe43__lane4_strm1_cntl          ( std__pe43__lane4_strm1_cntl       ),      
               .std__pe43__lane4_strm1_data          ( std__pe43__lane4_strm1_data       ),      
               .std__pe43__lane4_strm1_data_valid    ( std__pe43__lane4_strm1_data_valid ),      
               .std__pe43__lane4_strm1_data_mask     ( std__pe43__lane4_strm1_data_mask  ),      

               // PE 43, Lane 5                 
               .pe43__std__lane5_strm0_ready         ( pe43__std__lane5_strm0_ready      ),      
               .std__pe43__lane5_strm0_cntl          ( std__pe43__lane5_strm0_cntl       ),      
               .std__pe43__lane5_strm0_data          ( std__pe43__lane5_strm0_data       ),      
               .std__pe43__lane5_strm0_data_valid    ( std__pe43__lane5_strm0_data_valid ),      
               .std__pe43__lane5_strm0_data_mask     ( std__pe43__lane5_strm0_data_mask  ),      

               .pe43__std__lane5_strm1_ready         ( pe43__std__lane5_strm1_ready      ),      
               .std__pe43__lane5_strm1_cntl          ( std__pe43__lane5_strm1_cntl       ),      
               .std__pe43__lane5_strm1_data          ( std__pe43__lane5_strm1_data       ),      
               .std__pe43__lane5_strm1_data_valid    ( std__pe43__lane5_strm1_data_valid ),      
               .std__pe43__lane5_strm1_data_mask     ( std__pe43__lane5_strm1_data_mask  ),      

               // PE 43, Lane 6                 
               .pe43__std__lane6_strm0_ready         ( pe43__std__lane6_strm0_ready      ),      
               .std__pe43__lane6_strm0_cntl          ( std__pe43__lane6_strm0_cntl       ),      
               .std__pe43__lane6_strm0_data          ( std__pe43__lane6_strm0_data       ),      
               .std__pe43__lane6_strm0_data_valid    ( std__pe43__lane6_strm0_data_valid ),      
               .std__pe43__lane6_strm0_data_mask     ( std__pe43__lane6_strm0_data_mask  ),      

               .pe43__std__lane6_strm1_ready         ( pe43__std__lane6_strm1_ready      ),      
               .std__pe43__lane6_strm1_cntl          ( std__pe43__lane6_strm1_cntl       ),      
               .std__pe43__lane6_strm1_data          ( std__pe43__lane6_strm1_data       ),      
               .std__pe43__lane6_strm1_data_valid    ( std__pe43__lane6_strm1_data_valid ),      
               .std__pe43__lane6_strm1_data_mask     ( std__pe43__lane6_strm1_data_mask  ),      

               // PE 43, Lane 7                 
               .pe43__std__lane7_strm0_ready         ( pe43__std__lane7_strm0_ready      ),      
               .std__pe43__lane7_strm0_cntl          ( std__pe43__lane7_strm0_cntl       ),      
               .std__pe43__lane7_strm0_data          ( std__pe43__lane7_strm0_data       ),      
               .std__pe43__lane7_strm0_data_valid    ( std__pe43__lane7_strm0_data_valid ),      
               .std__pe43__lane7_strm0_data_mask     ( std__pe43__lane7_strm0_data_mask  ),      

               .pe43__std__lane7_strm1_ready         ( pe43__std__lane7_strm1_ready      ),      
               .std__pe43__lane7_strm1_cntl          ( std__pe43__lane7_strm1_cntl       ),      
               .std__pe43__lane7_strm1_data          ( std__pe43__lane7_strm1_data       ),      
               .std__pe43__lane7_strm1_data_valid    ( std__pe43__lane7_strm1_data_valid ),      
               .std__pe43__lane7_strm1_data_mask     ( std__pe43__lane7_strm1_data_mask  ),      

               // PE 43, Lane 8                 
               .pe43__std__lane8_strm0_ready         ( pe43__std__lane8_strm0_ready      ),      
               .std__pe43__lane8_strm0_cntl          ( std__pe43__lane8_strm0_cntl       ),      
               .std__pe43__lane8_strm0_data          ( std__pe43__lane8_strm0_data       ),      
               .std__pe43__lane8_strm0_data_valid    ( std__pe43__lane8_strm0_data_valid ),      
               .std__pe43__lane8_strm0_data_mask     ( std__pe43__lane8_strm0_data_mask  ),      

               .pe43__std__lane8_strm1_ready         ( pe43__std__lane8_strm1_ready      ),      
               .std__pe43__lane8_strm1_cntl          ( std__pe43__lane8_strm1_cntl       ),      
               .std__pe43__lane8_strm1_data          ( std__pe43__lane8_strm1_data       ),      
               .std__pe43__lane8_strm1_data_valid    ( std__pe43__lane8_strm1_data_valid ),      
               .std__pe43__lane8_strm1_data_mask     ( std__pe43__lane8_strm1_data_mask  ),      

               // PE 43, Lane 9                 
               .pe43__std__lane9_strm0_ready         ( pe43__std__lane9_strm0_ready      ),      
               .std__pe43__lane9_strm0_cntl          ( std__pe43__lane9_strm0_cntl       ),      
               .std__pe43__lane9_strm0_data          ( std__pe43__lane9_strm0_data       ),      
               .std__pe43__lane9_strm0_data_valid    ( std__pe43__lane9_strm0_data_valid ),      
               .std__pe43__lane9_strm0_data_mask     ( std__pe43__lane9_strm0_data_mask  ),      

               .pe43__std__lane9_strm1_ready         ( pe43__std__lane9_strm1_ready      ),      
               .std__pe43__lane9_strm1_cntl          ( std__pe43__lane9_strm1_cntl       ),      
               .std__pe43__lane9_strm1_data          ( std__pe43__lane9_strm1_data       ),      
               .std__pe43__lane9_strm1_data_valid    ( std__pe43__lane9_strm1_data_valid ),      
               .std__pe43__lane9_strm1_data_mask     ( std__pe43__lane9_strm1_data_mask  ),      

               // PE 43, Lane 10                 
               .pe43__std__lane10_strm0_ready         ( pe43__std__lane10_strm0_ready      ),      
               .std__pe43__lane10_strm0_cntl          ( std__pe43__lane10_strm0_cntl       ),      
               .std__pe43__lane10_strm0_data          ( std__pe43__lane10_strm0_data       ),      
               .std__pe43__lane10_strm0_data_valid    ( std__pe43__lane10_strm0_data_valid ),      
               .std__pe43__lane10_strm0_data_mask     ( std__pe43__lane10_strm0_data_mask  ),      

               .pe43__std__lane10_strm1_ready         ( pe43__std__lane10_strm1_ready      ),      
               .std__pe43__lane10_strm1_cntl          ( std__pe43__lane10_strm1_cntl       ),      
               .std__pe43__lane10_strm1_data          ( std__pe43__lane10_strm1_data       ),      
               .std__pe43__lane10_strm1_data_valid    ( std__pe43__lane10_strm1_data_valid ),      
               .std__pe43__lane10_strm1_data_mask     ( std__pe43__lane10_strm1_data_mask  ),      

               // PE 43, Lane 11                 
               .pe43__std__lane11_strm0_ready         ( pe43__std__lane11_strm0_ready      ),      
               .std__pe43__lane11_strm0_cntl          ( std__pe43__lane11_strm0_cntl       ),      
               .std__pe43__lane11_strm0_data          ( std__pe43__lane11_strm0_data       ),      
               .std__pe43__lane11_strm0_data_valid    ( std__pe43__lane11_strm0_data_valid ),      
               .std__pe43__lane11_strm0_data_mask     ( std__pe43__lane11_strm0_data_mask  ),      

               .pe43__std__lane11_strm1_ready         ( pe43__std__lane11_strm1_ready      ),      
               .std__pe43__lane11_strm1_cntl          ( std__pe43__lane11_strm1_cntl       ),      
               .std__pe43__lane11_strm1_data          ( std__pe43__lane11_strm1_data       ),      
               .std__pe43__lane11_strm1_data_valid    ( std__pe43__lane11_strm1_data_valid ),      
               .std__pe43__lane11_strm1_data_mask     ( std__pe43__lane11_strm1_data_mask  ),      

               // PE 43, Lane 12                 
               .pe43__std__lane12_strm0_ready         ( pe43__std__lane12_strm0_ready      ),      
               .std__pe43__lane12_strm0_cntl          ( std__pe43__lane12_strm0_cntl       ),      
               .std__pe43__lane12_strm0_data          ( std__pe43__lane12_strm0_data       ),      
               .std__pe43__lane12_strm0_data_valid    ( std__pe43__lane12_strm0_data_valid ),      
               .std__pe43__lane12_strm0_data_mask     ( std__pe43__lane12_strm0_data_mask  ),      

               .pe43__std__lane12_strm1_ready         ( pe43__std__lane12_strm1_ready      ),      
               .std__pe43__lane12_strm1_cntl          ( std__pe43__lane12_strm1_cntl       ),      
               .std__pe43__lane12_strm1_data          ( std__pe43__lane12_strm1_data       ),      
               .std__pe43__lane12_strm1_data_valid    ( std__pe43__lane12_strm1_data_valid ),      
               .std__pe43__lane12_strm1_data_mask     ( std__pe43__lane12_strm1_data_mask  ),      

               // PE 43, Lane 13                 
               .pe43__std__lane13_strm0_ready         ( pe43__std__lane13_strm0_ready      ),      
               .std__pe43__lane13_strm0_cntl          ( std__pe43__lane13_strm0_cntl       ),      
               .std__pe43__lane13_strm0_data          ( std__pe43__lane13_strm0_data       ),      
               .std__pe43__lane13_strm0_data_valid    ( std__pe43__lane13_strm0_data_valid ),      
               .std__pe43__lane13_strm0_data_mask     ( std__pe43__lane13_strm0_data_mask  ),      

               .pe43__std__lane13_strm1_ready         ( pe43__std__lane13_strm1_ready      ),      
               .std__pe43__lane13_strm1_cntl          ( std__pe43__lane13_strm1_cntl       ),      
               .std__pe43__lane13_strm1_data          ( std__pe43__lane13_strm1_data       ),      
               .std__pe43__lane13_strm1_data_valid    ( std__pe43__lane13_strm1_data_valid ),      
               .std__pe43__lane13_strm1_data_mask     ( std__pe43__lane13_strm1_data_mask  ),      

               // PE 43, Lane 14                 
               .pe43__std__lane14_strm0_ready         ( pe43__std__lane14_strm0_ready      ),      
               .std__pe43__lane14_strm0_cntl          ( std__pe43__lane14_strm0_cntl       ),      
               .std__pe43__lane14_strm0_data          ( std__pe43__lane14_strm0_data       ),      
               .std__pe43__lane14_strm0_data_valid    ( std__pe43__lane14_strm0_data_valid ),      
               .std__pe43__lane14_strm0_data_mask     ( std__pe43__lane14_strm0_data_mask  ),      

               .pe43__std__lane14_strm1_ready         ( pe43__std__lane14_strm1_ready      ),      
               .std__pe43__lane14_strm1_cntl          ( std__pe43__lane14_strm1_cntl       ),      
               .std__pe43__lane14_strm1_data          ( std__pe43__lane14_strm1_data       ),      
               .std__pe43__lane14_strm1_data_valid    ( std__pe43__lane14_strm1_data_valid ),      
               .std__pe43__lane14_strm1_data_mask     ( std__pe43__lane14_strm1_data_mask  ),      

               // PE 43, Lane 15                 
               .pe43__std__lane15_strm0_ready         ( pe43__std__lane15_strm0_ready      ),      
               .std__pe43__lane15_strm0_cntl          ( std__pe43__lane15_strm0_cntl       ),      
               .std__pe43__lane15_strm0_data          ( std__pe43__lane15_strm0_data       ),      
               .std__pe43__lane15_strm0_data_valid    ( std__pe43__lane15_strm0_data_valid ),      
               .std__pe43__lane15_strm0_data_mask     ( std__pe43__lane15_strm0_data_mask  ),      

               .pe43__std__lane15_strm1_ready         ( pe43__std__lane15_strm1_ready      ),      
               .std__pe43__lane15_strm1_cntl          ( std__pe43__lane15_strm1_cntl       ),      
               .std__pe43__lane15_strm1_data          ( std__pe43__lane15_strm1_data       ),      
               .std__pe43__lane15_strm1_data_valid    ( std__pe43__lane15_strm1_data_valid ),      
               .std__pe43__lane15_strm1_data_mask     ( std__pe43__lane15_strm1_data_mask  ),      

               // PE 43, Lane 16                 
               .pe43__std__lane16_strm0_ready         ( pe43__std__lane16_strm0_ready      ),      
               .std__pe43__lane16_strm0_cntl          ( std__pe43__lane16_strm0_cntl       ),      
               .std__pe43__lane16_strm0_data          ( std__pe43__lane16_strm0_data       ),      
               .std__pe43__lane16_strm0_data_valid    ( std__pe43__lane16_strm0_data_valid ),      
               .std__pe43__lane16_strm0_data_mask     ( std__pe43__lane16_strm0_data_mask  ),      

               .pe43__std__lane16_strm1_ready         ( pe43__std__lane16_strm1_ready      ),      
               .std__pe43__lane16_strm1_cntl          ( std__pe43__lane16_strm1_cntl       ),      
               .std__pe43__lane16_strm1_data          ( std__pe43__lane16_strm1_data       ),      
               .std__pe43__lane16_strm1_data_valid    ( std__pe43__lane16_strm1_data_valid ),      
               .std__pe43__lane16_strm1_data_mask     ( std__pe43__lane16_strm1_data_mask  ),      

               // PE 43, Lane 17                 
               .pe43__std__lane17_strm0_ready         ( pe43__std__lane17_strm0_ready      ),      
               .std__pe43__lane17_strm0_cntl          ( std__pe43__lane17_strm0_cntl       ),      
               .std__pe43__lane17_strm0_data          ( std__pe43__lane17_strm0_data       ),      
               .std__pe43__lane17_strm0_data_valid    ( std__pe43__lane17_strm0_data_valid ),      
               .std__pe43__lane17_strm0_data_mask     ( std__pe43__lane17_strm0_data_mask  ),      

               .pe43__std__lane17_strm1_ready         ( pe43__std__lane17_strm1_ready      ),      
               .std__pe43__lane17_strm1_cntl          ( std__pe43__lane17_strm1_cntl       ),      
               .std__pe43__lane17_strm1_data          ( std__pe43__lane17_strm1_data       ),      
               .std__pe43__lane17_strm1_data_valid    ( std__pe43__lane17_strm1_data_valid ),      
               .std__pe43__lane17_strm1_data_mask     ( std__pe43__lane17_strm1_data_mask  ),      

               // PE 43, Lane 18                 
               .pe43__std__lane18_strm0_ready         ( pe43__std__lane18_strm0_ready      ),      
               .std__pe43__lane18_strm0_cntl          ( std__pe43__lane18_strm0_cntl       ),      
               .std__pe43__lane18_strm0_data          ( std__pe43__lane18_strm0_data       ),      
               .std__pe43__lane18_strm0_data_valid    ( std__pe43__lane18_strm0_data_valid ),      
               .std__pe43__lane18_strm0_data_mask     ( std__pe43__lane18_strm0_data_mask  ),      

               .pe43__std__lane18_strm1_ready         ( pe43__std__lane18_strm1_ready      ),      
               .std__pe43__lane18_strm1_cntl          ( std__pe43__lane18_strm1_cntl       ),      
               .std__pe43__lane18_strm1_data          ( std__pe43__lane18_strm1_data       ),      
               .std__pe43__lane18_strm1_data_valid    ( std__pe43__lane18_strm1_data_valid ),      
               .std__pe43__lane18_strm1_data_mask     ( std__pe43__lane18_strm1_data_mask  ),      

               // PE 43, Lane 19                 
               .pe43__std__lane19_strm0_ready         ( pe43__std__lane19_strm0_ready      ),      
               .std__pe43__lane19_strm0_cntl          ( std__pe43__lane19_strm0_cntl       ),      
               .std__pe43__lane19_strm0_data          ( std__pe43__lane19_strm0_data       ),      
               .std__pe43__lane19_strm0_data_valid    ( std__pe43__lane19_strm0_data_valid ),      
               .std__pe43__lane19_strm0_data_mask     ( std__pe43__lane19_strm0_data_mask  ),      

               .pe43__std__lane19_strm1_ready         ( pe43__std__lane19_strm1_ready      ),      
               .std__pe43__lane19_strm1_cntl          ( std__pe43__lane19_strm1_cntl       ),      
               .std__pe43__lane19_strm1_data          ( std__pe43__lane19_strm1_data       ),      
               .std__pe43__lane19_strm1_data_valid    ( std__pe43__lane19_strm1_data_valid ),      
               .std__pe43__lane19_strm1_data_mask     ( std__pe43__lane19_strm1_data_mask  ),      

               // PE 43, Lane 20                 
               .pe43__std__lane20_strm0_ready         ( pe43__std__lane20_strm0_ready      ),      
               .std__pe43__lane20_strm0_cntl          ( std__pe43__lane20_strm0_cntl       ),      
               .std__pe43__lane20_strm0_data          ( std__pe43__lane20_strm0_data       ),      
               .std__pe43__lane20_strm0_data_valid    ( std__pe43__lane20_strm0_data_valid ),      
               .std__pe43__lane20_strm0_data_mask     ( std__pe43__lane20_strm0_data_mask  ),      

               .pe43__std__lane20_strm1_ready         ( pe43__std__lane20_strm1_ready      ),      
               .std__pe43__lane20_strm1_cntl          ( std__pe43__lane20_strm1_cntl       ),      
               .std__pe43__lane20_strm1_data          ( std__pe43__lane20_strm1_data       ),      
               .std__pe43__lane20_strm1_data_valid    ( std__pe43__lane20_strm1_data_valid ),      
               .std__pe43__lane20_strm1_data_mask     ( std__pe43__lane20_strm1_data_mask  ),      

               // PE 43, Lane 21                 
               .pe43__std__lane21_strm0_ready         ( pe43__std__lane21_strm0_ready      ),      
               .std__pe43__lane21_strm0_cntl          ( std__pe43__lane21_strm0_cntl       ),      
               .std__pe43__lane21_strm0_data          ( std__pe43__lane21_strm0_data       ),      
               .std__pe43__lane21_strm0_data_valid    ( std__pe43__lane21_strm0_data_valid ),      
               .std__pe43__lane21_strm0_data_mask     ( std__pe43__lane21_strm0_data_mask  ),      

               .pe43__std__lane21_strm1_ready         ( pe43__std__lane21_strm1_ready      ),      
               .std__pe43__lane21_strm1_cntl          ( std__pe43__lane21_strm1_cntl       ),      
               .std__pe43__lane21_strm1_data          ( std__pe43__lane21_strm1_data       ),      
               .std__pe43__lane21_strm1_data_valid    ( std__pe43__lane21_strm1_data_valid ),      
               .std__pe43__lane21_strm1_data_mask     ( std__pe43__lane21_strm1_data_mask  ),      

               // PE 43, Lane 22                 
               .pe43__std__lane22_strm0_ready         ( pe43__std__lane22_strm0_ready      ),      
               .std__pe43__lane22_strm0_cntl          ( std__pe43__lane22_strm0_cntl       ),      
               .std__pe43__lane22_strm0_data          ( std__pe43__lane22_strm0_data       ),      
               .std__pe43__lane22_strm0_data_valid    ( std__pe43__lane22_strm0_data_valid ),      
               .std__pe43__lane22_strm0_data_mask     ( std__pe43__lane22_strm0_data_mask  ),      

               .pe43__std__lane22_strm1_ready         ( pe43__std__lane22_strm1_ready      ),      
               .std__pe43__lane22_strm1_cntl          ( std__pe43__lane22_strm1_cntl       ),      
               .std__pe43__lane22_strm1_data          ( std__pe43__lane22_strm1_data       ),      
               .std__pe43__lane22_strm1_data_valid    ( std__pe43__lane22_strm1_data_valid ),      
               .std__pe43__lane22_strm1_data_mask     ( std__pe43__lane22_strm1_data_mask  ),      

               // PE 43, Lane 23                 
               .pe43__std__lane23_strm0_ready         ( pe43__std__lane23_strm0_ready      ),      
               .std__pe43__lane23_strm0_cntl          ( std__pe43__lane23_strm0_cntl       ),      
               .std__pe43__lane23_strm0_data          ( std__pe43__lane23_strm0_data       ),      
               .std__pe43__lane23_strm0_data_valid    ( std__pe43__lane23_strm0_data_valid ),      
               .std__pe43__lane23_strm0_data_mask     ( std__pe43__lane23_strm0_data_mask  ),      

               .pe43__std__lane23_strm1_ready         ( pe43__std__lane23_strm1_ready      ),      
               .std__pe43__lane23_strm1_cntl          ( std__pe43__lane23_strm1_cntl       ),      
               .std__pe43__lane23_strm1_data          ( std__pe43__lane23_strm1_data       ),      
               .std__pe43__lane23_strm1_data_valid    ( std__pe43__lane23_strm1_data_valid ),      
               .std__pe43__lane23_strm1_data_mask     ( std__pe43__lane23_strm1_data_mask  ),      

               // PE 43, Lane 24                 
               .pe43__std__lane24_strm0_ready         ( pe43__std__lane24_strm0_ready      ),      
               .std__pe43__lane24_strm0_cntl          ( std__pe43__lane24_strm0_cntl       ),      
               .std__pe43__lane24_strm0_data          ( std__pe43__lane24_strm0_data       ),      
               .std__pe43__lane24_strm0_data_valid    ( std__pe43__lane24_strm0_data_valid ),      
               .std__pe43__lane24_strm0_data_mask     ( std__pe43__lane24_strm0_data_mask  ),      

               .pe43__std__lane24_strm1_ready         ( pe43__std__lane24_strm1_ready      ),      
               .std__pe43__lane24_strm1_cntl          ( std__pe43__lane24_strm1_cntl       ),      
               .std__pe43__lane24_strm1_data          ( std__pe43__lane24_strm1_data       ),      
               .std__pe43__lane24_strm1_data_valid    ( std__pe43__lane24_strm1_data_valid ),      
               .std__pe43__lane24_strm1_data_mask     ( std__pe43__lane24_strm1_data_mask  ),      

               // PE 43, Lane 25                 
               .pe43__std__lane25_strm0_ready         ( pe43__std__lane25_strm0_ready      ),      
               .std__pe43__lane25_strm0_cntl          ( std__pe43__lane25_strm0_cntl       ),      
               .std__pe43__lane25_strm0_data          ( std__pe43__lane25_strm0_data       ),      
               .std__pe43__lane25_strm0_data_valid    ( std__pe43__lane25_strm0_data_valid ),      
               .std__pe43__lane25_strm0_data_mask     ( std__pe43__lane25_strm0_data_mask  ),      

               .pe43__std__lane25_strm1_ready         ( pe43__std__lane25_strm1_ready      ),      
               .std__pe43__lane25_strm1_cntl          ( std__pe43__lane25_strm1_cntl       ),      
               .std__pe43__lane25_strm1_data          ( std__pe43__lane25_strm1_data       ),      
               .std__pe43__lane25_strm1_data_valid    ( std__pe43__lane25_strm1_data_valid ),      
               .std__pe43__lane25_strm1_data_mask     ( std__pe43__lane25_strm1_data_mask  ),      

               // PE 43, Lane 26                 
               .pe43__std__lane26_strm0_ready         ( pe43__std__lane26_strm0_ready      ),      
               .std__pe43__lane26_strm0_cntl          ( std__pe43__lane26_strm0_cntl       ),      
               .std__pe43__lane26_strm0_data          ( std__pe43__lane26_strm0_data       ),      
               .std__pe43__lane26_strm0_data_valid    ( std__pe43__lane26_strm0_data_valid ),      
               .std__pe43__lane26_strm0_data_mask     ( std__pe43__lane26_strm0_data_mask  ),      

               .pe43__std__lane26_strm1_ready         ( pe43__std__lane26_strm1_ready      ),      
               .std__pe43__lane26_strm1_cntl          ( std__pe43__lane26_strm1_cntl       ),      
               .std__pe43__lane26_strm1_data          ( std__pe43__lane26_strm1_data       ),      
               .std__pe43__lane26_strm1_data_valid    ( std__pe43__lane26_strm1_data_valid ),      
               .std__pe43__lane26_strm1_data_mask     ( std__pe43__lane26_strm1_data_mask  ),      

               // PE 43, Lane 27                 
               .pe43__std__lane27_strm0_ready         ( pe43__std__lane27_strm0_ready      ),      
               .std__pe43__lane27_strm0_cntl          ( std__pe43__lane27_strm0_cntl       ),      
               .std__pe43__lane27_strm0_data          ( std__pe43__lane27_strm0_data       ),      
               .std__pe43__lane27_strm0_data_valid    ( std__pe43__lane27_strm0_data_valid ),      
               .std__pe43__lane27_strm0_data_mask     ( std__pe43__lane27_strm0_data_mask  ),      

               .pe43__std__lane27_strm1_ready         ( pe43__std__lane27_strm1_ready      ),      
               .std__pe43__lane27_strm1_cntl          ( std__pe43__lane27_strm1_cntl       ),      
               .std__pe43__lane27_strm1_data          ( std__pe43__lane27_strm1_data       ),      
               .std__pe43__lane27_strm1_data_valid    ( std__pe43__lane27_strm1_data_valid ),      
               .std__pe43__lane27_strm1_data_mask     ( std__pe43__lane27_strm1_data_mask  ),      

               // PE 43, Lane 28                 
               .pe43__std__lane28_strm0_ready         ( pe43__std__lane28_strm0_ready      ),      
               .std__pe43__lane28_strm0_cntl          ( std__pe43__lane28_strm0_cntl       ),      
               .std__pe43__lane28_strm0_data          ( std__pe43__lane28_strm0_data       ),      
               .std__pe43__lane28_strm0_data_valid    ( std__pe43__lane28_strm0_data_valid ),      
               .std__pe43__lane28_strm0_data_mask     ( std__pe43__lane28_strm0_data_mask  ),      

               .pe43__std__lane28_strm1_ready         ( pe43__std__lane28_strm1_ready      ),      
               .std__pe43__lane28_strm1_cntl          ( std__pe43__lane28_strm1_cntl       ),      
               .std__pe43__lane28_strm1_data          ( std__pe43__lane28_strm1_data       ),      
               .std__pe43__lane28_strm1_data_valid    ( std__pe43__lane28_strm1_data_valid ),      
               .std__pe43__lane28_strm1_data_mask     ( std__pe43__lane28_strm1_data_mask  ),      

               // PE 43, Lane 29                 
               .pe43__std__lane29_strm0_ready         ( pe43__std__lane29_strm0_ready      ),      
               .std__pe43__lane29_strm0_cntl          ( std__pe43__lane29_strm0_cntl       ),      
               .std__pe43__lane29_strm0_data          ( std__pe43__lane29_strm0_data       ),      
               .std__pe43__lane29_strm0_data_valid    ( std__pe43__lane29_strm0_data_valid ),      
               .std__pe43__lane29_strm0_data_mask     ( std__pe43__lane29_strm0_data_mask  ),      

               .pe43__std__lane29_strm1_ready         ( pe43__std__lane29_strm1_ready      ),      
               .std__pe43__lane29_strm1_cntl          ( std__pe43__lane29_strm1_cntl       ),      
               .std__pe43__lane29_strm1_data          ( std__pe43__lane29_strm1_data       ),      
               .std__pe43__lane29_strm1_data_valid    ( std__pe43__lane29_strm1_data_valid ),      
               .std__pe43__lane29_strm1_data_mask     ( std__pe43__lane29_strm1_data_mask  ),      

               // PE 43, Lane 30                 
               .pe43__std__lane30_strm0_ready         ( pe43__std__lane30_strm0_ready      ),      
               .std__pe43__lane30_strm0_cntl          ( std__pe43__lane30_strm0_cntl       ),      
               .std__pe43__lane30_strm0_data          ( std__pe43__lane30_strm0_data       ),      
               .std__pe43__lane30_strm0_data_valid    ( std__pe43__lane30_strm0_data_valid ),      
               .std__pe43__lane30_strm0_data_mask     ( std__pe43__lane30_strm0_data_mask  ),      

               .pe43__std__lane30_strm1_ready         ( pe43__std__lane30_strm1_ready      ),      
               .std__pe43__lane30_strm1_cntl          ( std__pe43__lane30_strm1_cntl       ),      
               .std__pe43__lane30_strm1_data          ( std__pe43__lane30_strm1_data       ),      
               .std__pe43__lane30_strm1_data_valid    ( std__pe43__lane30_strm1_data_valid ),      
               .std__pe43__lane30_strm1_data_mask     ( std__pe43__lane30_strm1_data_mask  ),      

               // PE 43, Lane 31                 
               .pe43__std__lane31_strm0_ready         ( pe43__std__lane31_strm0_ready      ),      
               .std__pe43__lane31_strm0_cntl          ( std__pe43__lane31_strm0_cntl       ),      
               .std__pe43__lane31_strm0_data          ( std__pe43__lane31_strm0_data       ),      
               .std__pe43__lane31_strm0_data_valid    ( std__pe43__lane31_strm0_data_valid ),      
               .std__pe43__lane31_strm0_data_mask     ( std__pe43__lane31_strm0_data_mask  ),      

               .pe43__std__lane31_strm1_ready         ( pe43__std__lane31_strm1_ready      ),      
               .std__pe43__lane31_strm1_cntl          ( std__pe43__lane31_strm1_cntl       ),      
               .std__pe43__lane31_strm1_data          ( std__pe43__lane31_strm1_data       ),      
               .std__pe43__lane31_strm1_data_valid    ( std__pe43__lane31_strm1_data_valid ),      
               .std__pe43__lane31_strm1_data_mask     ( std__pe43__lane31_strm1_data_mask  ),      

               // PE 44, Lane 0                 
               .pe44__std__lane0_strm0_ready         ( pe44__std__lane0_strm0_ready      ),      
               .std__pe44__lane0_strm0_cntl          ( std__pe44__lane0_strm0_cntl       ),      
               .std__pe44__lane0_strm0_data          ( std__pe44__lane0_strm0_data       ),      
               .std__pe44__lane0_strm0_data_valid    ( std__pe44__lane0_strm0_data_valid ),      
               .std__pe44__lane0_strm0_data_mask     ( std__pe44__lane0_strm0_data_mask  ),      

               .pe44__std__lane0_strm1_ready         ( pe44__std__lane0_strm1_ready      ),      
               .std__pe44__lane0_strm1_cntl          ( std__pe44__lane0_strm1_cntl       ),      
               .std__pe44__lane0_strm1_data          ( std__pe44__lane0_strm1_data       ),      
               .std__pe44__lane0_strm1_data_valid    ( std__pe44__lane0_strm1_data_valid ),      
               .std__pe44__lane0_strm1_data_mask     ( std__pe44__lane0_strm1_data_mask  ),      

               // PE 44, Lane 1                 
               .pe44__std__lane1_strm0_ready         ( pe44__std__lane1_strm0_ready      ),      
               .std__pe44__lane1_strm0_cntl          ( std__pe44__lane1_strm0_cntl       ),      
               .std__pe44__lane1_strm0_data          ( std__pe44__lane1_strm0_data       ),      
               .std__pe44__lane1_strm0_data_valid    ( std__pe44__lane1_strm0_data_valid ),      
               .std__pe44__lane1_strm0_data_mask     ( std__pe44__lane1_strm0_data_mask  ),      

               .pe44__std__lane1_strm1_ready         ( pe44__std__lane1_strm1_ready      ),      
               .std__pe44__lane1_strm1_cntl          ( std__pe44__lane1_strm1_cntl       ),      
               .std__pe44__lane1_strm1_data          ( std__pe44__lane1_strm1_data       ),      
               .std__pe44__lane1_strm1_data_valid    ( std__pe44__lane1_strm1_data_valid ),      
               .std__pe44__lane1_strm1_data_mask     ( std__pe44__lane1_strm1_data_mask  ),      

               // PE 44, Lane 2                 
               .pe44__std__lane2_strm0_ready         ( pe44__std__lane2_strm0_ready      ),      
               .std__pe44__lane2_strm0_cntl          ( std__pe44__lane2_strm0_cntl       ),      
               .std__pe44__lane2_strm0_data          ( std__pe44__lane2_strm0_data       ),      
               .std__pe44__lane2_strm0_data_valid    ( std__pe44__lane2_strm0_data_valid ),      
               .std__pe44__lane2_strm0_data_mask     ( std__pe44__lane2_strm0_data_mask  ),      

               .pe44__std__lane2_strm1_ready         ( pe44__std__lane2_strm1_ready      ),      
               .std__pe44__lane2_strm1_cntl          ( std__pe44__lane2_strm1_cntl       ),      
               .std__pe44__lane2_strm1_data          ( std__pe44__lane2_strm1_data       ),      
               .std__pe44__lane2_strm1_data_valid    ( std__pe44__lane2_strm1_data_valid ),      
               .std__pe44__lane2_strm1_data_mask     ( std__pe44__lane2_strm1_data_mask  ),      

               // PE 44, Lane 3                 
               .pe44__std__lane3_strm0_ready         ( pe44__std__lane3_strm0_ready      ),      
               .std__pe44__lane3_strm0_cntl          ( std__pe44__lane3_strm0_cntl       ),      
               .std__pe44__lane3_strm0_data          ( std__pe44__lane3_strm0_data       ),      
               .std__pe44__lane3_strm0_data_valid    ( std__pe44__lane3_strm0_data_valid ),      
               .std__pe44__lane3_strm0_data_mask     ( std__pe44__lane3_strm0_data_mask  ),      

               .pe44__std__lane3_strm1_ready         ( pe44__std__lane3_strm1_ready      ),      
               .std__pe44__lane3_strm1_cntl          ( std__pe44__lane3_strm1_cntl       ),      
               .std__pe44__lane3_strm1_data          ( std__pe44__lane3_strm1_data       ),      
               .std__pe44__lane3_strm1_data_valid    ( std__pe44__lane3_strm1_data_valid ),      
               .std__pe44__lane3_strm1_data_mask     ( std__pe44__lane3_strm1_data_mask  ),      

               // PE 44, Lane 4                 
               .pe44__std__lane4_strm0_ready         ( pe44__std__lane4_strm0_ready      ),      
               .std__pe44__lane4_strm0_cntl          ( std__pe44__lane4_strm0_cntl       ),      
               .std__pe44__lane4_strm0_data          ( std__pe44__lane4_strm0_data       ),      
               .std__pe44__lane4_strm0_data_valid    ( std__pe44__lane4_strm0_data_valid ),      
               .std__pe44__lane4_strm0_data_mask     ( std__pe44__lane4_strm0_data_mask  ),      

               .pe44__std__lane4_strm1_ready         ( pe44__std__lane4_strm1_ready      ),      
               .std__pe44__lane4_strm1_cntl          ( std__pe44__lane4_strm1_cntl       ),      
               .std__pe44__lane4_strm1_data          ( std__pe44__lane4_strm1_data       ),      
               .std__pe44__lane4_strm1_data_valid    ( std__pe44__lane4_strm1_data_valid ),      
               .std__pe44__lane4_strm1_data_mask     ( std__pe44__lane4_strm1_data_mask  ),      

               // PE 44, Lane 5                 
               .pe44__std__lane5_strm0_ready         ( pe44__std__lane5_strm0_ready      ),      
               .std__pe44__lane5_strm0_cntl          ( std__pe44__lane5_strm0_cntl       ),      
               .std__pe44__lane5_strm0_data          ( std__pe44__lane5_strm0_data       ),      
               .std__pe44__lane5_strm0_data_valid    ( std__pe44__lane5_strm0_data_valid ),      
               .std__pe44__lane5_strm0_data_mask     ( std__pe44__lane5_strm0_data_mask  ),      

               .pe44__std__lane5_strm1_ready         ( pe44__std__lane5_strm1_ready      ),      
               .std__pe44__lane5_strm1_cntl          ( std__pe44__lane5_strm1_cntl       ),      
               .std__pe44__lane5_strm1_data          ( std__pe44__lane5_strm1_data       ),      
               .std__pe44__lane5_strm1_data_valid    ( std__pe44__lane5_strm1_data_valid ),      
               .std__pe44__lane5_strm1_data_mask     ( std__pe44__lane5_strm1_data_mask  ),      

               // PE 44, Lane 6                 
               .pe44__std__lane6_strm0_ready         ( pe44__std__lane6_strm0_ready      ),      
               .std__pe44__lane6_strm0_cntl          ( std__pe44__lane6_strm0_cntl       ),      
               .std__pe44__lane6_strm0_data          ( std__pe44__lane6_strm0_data       ),      
               .std__pe44__lane6_strm0_data_valid    ( std__pe44__lane6_strm0_data_valid ),      
               .std__pe44__lane6_strm0_data_mask     ( std__pe44__lane6_strm0_data_mask  ),      

               .pe44__std__lane6_strm1_ready         ( pe44__std__lane6_strm1_ready      ),      
               .std__pe44__lane6_strm1_cntl          ( std__pe44__lane6_strm1_cntl       ),      
               .std__pe44__lane6_strm1_data          ( std__pe44__lane6_strm1_data       ),      
               .std__pe44__lane6_strm1_data_valid    ( std__pe44__lane6_strm1_data_valid ),      
               .std__pe44__lane6_strm1_data_mask     ( std__pe44__lane6_strm1_data_mask  ),      

               // PE 44, Lane 7                 
               .pe44__std__lane7_strm0_ready         ( pe44__std__lane7_strm0_ready      ),      
               .std__pe44__lane7_strm0_cntl          ( std__pe44__lane7_strm0_cntl       ),      
               .std__pe44__lane7_strm0_data          ( std__pe44__lane7_strm0_data       ),      
               .std__pe44__lane7_strm0_data_valid    ( std__pe44__lane7_strm0_data_valid ),      
               .std__pe44__lane7_strm0_data_mask     ( std__pe44__lane7_strm0_data_mask  ),      

               .pe44__std__lane7_strm1_ready         ( pe44__std__lane7_strm1_ready      ),      
               .std__pe44__lane7_strm1_cntl          ( std__pe44__lane7_strm1_cntl       ),      
               .std__pe44__lane7_strm1_data          ( std__pe44__lane7_strm1_data       ),      
               .std__pe44__lane7_strm1_data_valid    ( std__pe44__lane7_strm1_data_valid ),      
               .std__pe44__lane7_strm1_data_mask     ( std__pe44__lane7_strm1_data_mask  ),      

               // PE 44, Lane 8                 
               .pe44__std__lane8_strm0_ready         ( pe44__std__lane8_strm0_ready      ),      
               .std__pe44__lane8_strm0_cntl          ( std__pe44__lane8_strm0_cntl       ),      
               .std__pe44__lane8_strm0_data          ( std__pe44__lane8_strm0_data       ),      
               .std__pe44__lane8_strm0_data_valid    ( std__pe44__lane8_strm0_data_valid ),      
               .std__pe44__lane8_strm0_data_mask     ( std__pe44__lane8_strm0_data_mask  ),      

               .pe44__std__lane8_strm1_ready         ( pe44__std__lane8_strm1_ready      ),      
               .std__pe44__lane8_strm1_cntl          ( std__pe44__lane8_strm1_cntl       ),      
               .std__pe44__lane8_strm1_data          ( std__pe44__lane8_strm1_data       ),      
               .std__pe44__lane8_strm1_data_valid    ( std__pe44__lane8_strm1_data_valid ),      
               .std__pe44__lane8_strm1_data_mask     ( std__pe44__lane8_strm1_data_mask  ),      

               // PE 44, Lane 9                 
               .pe44__std__lane9_strm0_ready         ( pe44__std__lane9_strm0_ready      ),      
               .std__pe44__lane9_strm0_cntl          ( std__pe44__lane9_strm0_cntl       ),      
               .std__pe44__lane9_strm0_data          ( std__pe44__lane9_strm0_data       ),      
               .std__pe44__lane9_strm0_data_valid    ( std__pe44__lane9_strm0_data_valid ),      
               .std__pe44__lane9_strm0_data_mask     ( std__pe44__lane9_strm0_data_mask  ),      

               .pe44__std__lane9_strm1_ready         ( pe44__std__lane9_strm1_ready      ),      
               .std__pe44__lane9_strm1_cntl          ( std__pe44__lane9_strm1_cntl       ),      
               .std__pe44__lane9_strm1_data          ( std__pe44__lane9_strm1_data       ),      
               .std__pe44__lane9_strm1_data_valid    ( std__pe44__lane9_strm1_data_valid ),      
               .std__pe44__lane9_strm1_data_mask     ( std__pe44__lane9_strm1_data_mask  ),      

               // PE 44, Lane 10                 
               .pe44__std__lane10_strm0_ready         ( pe44__std__lane10_strm0_ready      ),      
               .std__pe44__lane10_strm0_cntl          ( std__pe44__lane10_strm0_cntl       ),      
               .std__pe44__lane10_strm0_data          ( std__pe44__lane10_strm0_data       ),      
               .std__pe44__lane10_strm0_data_valid    ( std__pe44__lane10_strm0_data_valid ),      
               .std__pe44__lane10_strm0_data_mask     ( std__pe44__lane10_strm0_data_mask  ),      

               .pe44__std__lane10_strm1_ready         ( pe44__std__lane10_strm1_ready      ),      
               .std__pe44__lane10_strm1_cntl          ( std__pe44__lane10_strm1_cntl       ),      
               .std__pe44__lane10_strm1_data          ( std__pe44__lane10_strm1_data       ),      
               .std__pe44__lane10_strm1_data_valid    ( std__pe44__lane10_strm1_data_valid ),      
               .std__pe44__lane10_strm1_data_mask     ( std__pe44__lane10_strm1_data_mask  ),      

               // PE 44, Lane 11                 
               .pe44__std__lane11_strm0_ready         ( pe44__std__lane11_strm0_ready      ),      
               .std__pe44__lane11_strm0_cntl          ( std__pe44__lane11_strm0_cntl       ),      
               .std__pe44__lane11_strm0_data          ( std__pe44__lane11_strm0_data       ),      
               .std__pe44__lane11_strm0_data_valid    ( std__pe44__lane11_strm0_data_valid ),      
               .std__pe44__lane11_strm0_data_mask     ( std__pe44__lane11_strm0_data_mask  ),      

               .pe44__std__lane11_strm1_ready         ( pe44__std__lane11_strm1_ready      ),      
               .std__pe44__lane11_strm1_cntl          ( std__pe44__lane11_strm1_cntl       ),      
               .std__pe44__lane11_strm1_data          ( std__pe44__lane11_strm1_data       ),      
               .std__pe44__lane11_strm1_data_valid    ( std__pe44__lane11_strm1_data_valid ),      
               .std__pe44__lane11_strm1_data_mask     ( std__pe44__lane11_strm1_data_mask  ),      

               // PE 44, Lane 12                 
               .pe44__std__lane12_strm0_ready         ( pe44__std__lane12_strm0_ready      ),      
               .std__pe44__lane12_strm0_cntl          ( std__pe44__lane12_strm0_cntl       ),      
               .std__pe44__lane12_strm0_data          ( std__pe44__lane12_strm0_data       ),      
               .std__pe44__lane12_strm0_data_valid    ( std__pe44__lane12_strm0_data_valid ),      
               .std__pe44__lane12_strm0_data_mask     ( std__pe44__lane12_strm0_data_mask  ),      

               .pe44__std__lane12_strm1_ready         ( pe44__std__lane12_strm1_ready      ),      
               .std__pe44__lane12_strm1_cntl          ( std__pe44__lane12_strm1_cntl       ),      
               .std__pe44__lane12_strm1_data          ( std__pe44__lane12_strm1_data       ),      
               .std__pe44__lane12_strm1_data_valid    ( std__pe44__lane12_strm1_data_valid ),      
               .std__pe44__lane12_strm1_data_mask     ( std__pe44__lane12_strm1_data_mask  ),      

               // PE 44, Lane 13                 
               .pe44__std__lane13_strm0_ready         ( pe44__std__lane13_strm0_ready      ),      
               .std__pe44__lane13_strm0_cntl          ( std__pe44__lane13_strm0_cntl       ),      
               .std__pe44__lane13_strm0_data          ( std__pe44__lane13_strm0_data       ),      
               .std__pe44__lane13_strm0_data_valid    ( std__pe44__lane13_strm0_data_valid ),      
               .std__pe44__lane13_strm0_data_mask     ( std__pe44__lane13_strm0_data_mask  ),      

               .pe44__std__lane13_strm1_ready         ( pe44__std__lane13_strm1_ready      ),      
               .std__pe44__lane13_strm1_cntl          ( std__pe44__lane13_strm1_cntl       ),      
               .std__pe44__lane13_strm1_data          ( std__pe44__lane13_strm1_data       ),      
               .std__pe44__lane13_strm1_data_valid    ( std__pe44__lane13_strm1_data_valid ),      
               .std__pe44__lane13_strm1_data_mask     ( std__pe44__lane13_strm1_data_mask  ),      

               // PE 44, Lane 14                 
               .pe44__std__lane14_strm0_ready         ( pe44__std__lane14_strm0_ready      ),      
               .std__pe44__lane14_strm0_cntl          ( std__pe44__lane14_strm0_cntl       ),      
               .std__pe44__lane14_strm0_data          ( std__pe44__lane14_strm0_data       ),      
               .std__pe44__lane14_strm0_data_valid    ( std__pe44__lane14_strm0_data_valid ),      
               .std__pe44__lane14_strm0_data_mask     ( std__pe44__lane14_strm0_data_mask  ),      

               .pe44__std__lane14_strm1_ready         ( pe44__std__lane14_strm1_ready      ),      
               .std__pe44__lane14_strm1_cntl          ( std__pe44__lane14_strm1_cntl       ),      
               .std__pe44__lane14_strm1_data          ( std__pe44__lane14_strm1_data       ),      
               .std__pe44__lane14_strm1_data_valid    ( std__pe44__lane14_strm1_data_valid ),      
               .std__pe44__lane14_strm1_data_mask     ( std__pe44__lane14_strm1_data_mask  ),      

               // PE 44, Lane 15                 
               .pe44__std__lane15_strm0_ready         ( pe44__std__lane15_strm0_ready      ),      
               .std__pe44__lane15_strm0_cntl          ( std__pe44__lane15_strm0_cntl       ),      
               .std__pe44__lane15_strm0_data          ( std__pe44__lane15_strm0_data       ),      
               .std__pe44__lane15_strm0_data_valid    ( std__pe44__lane15_strm0_data_valid ),      
               .std__pe44__lane15_strm0_data_mask     ( std__pe44__lane15_strm0_data_mask  ),      

               .pe44__std__lane15_strm1_ready         ( pe44__std__lane15_strm1_ready      ),      
               .std__pe44__lane15_strm1_cntl          ( std__pe44__lane15_strm1_cntl       ),      
               .std__pe44__lane15_strm1_data          ( std__pe44__lane15_strm1_data       ),      
               .std__pe44__lane15_strm1_data_valid    ( std__pe44__lane15_strm1_data_valid ),      
               .std__pe44__lane15_strm1_data_mask     ( std__pe44__lane15_strm1_data_mask  ),      

               // PE 44, Lane 16                 
               .pe44__std__lane16_strm0_ready         ( pe44__std__lane16_strm0_ready      ),      
               .std__pe44__lane16_strm0_cntl          ( std__pe44__lane16_strm0_cntl       ),      
               .std__pe44__lane16_strm0_data          ( std__pe44__lane16_strm0_data       ),      
               .std__pe44__lane16_strm0_data_valid    ( std__pe44__lane16_strm0_data_valid ),      
               .std__pe44__lane16_strm0_data_mask     ( std__pe44__lane16_strm0_data_mask  ),      

               .pe44__std__lane16_strm1_ready         ( pe44__std__lane16_strm1_ready      ),      
               .std__pe44__lane16_strm1_cntl          ( std__pe44__lane16_strm1_cntl       ),      
               .std__pe44__lane16_strm1_data          ( std__pe44__lane16_strm1_data       ),      
               .std__pe44__lane16_strm1_data_valid    ( std__pe44__lane16_strm1_data_valid ),      
               .std__pe44__lane16_strm1_data_mask     ( std__pe44__lane16_strm1_data_mask  ),      

               // PE 44, Lane 17                 
               .pe44__std__lane17_strm0_ready         ( pe44__std__lane17_strm0_ready      ),      
               .std__pe44__lane17_strm0_cntl          ( std__pe44__lane17_strm0_cntl       ),      
               .std__pe44__lane17_strm0_data          ( std__pe44__lane17_strm0_data       ),      
               .std__pe44__lane17_strm0_data_valid    ( std__pe44__lane17_strm0_data_valid ),      
               .std__pe44__lane17_strm0_data_mask     ( std__pe44__lane17_strm0_data_mask  ),      

               .pe44__std__lane17_strm1_ready         ( pe44__std__lane17_strm1_ready      ),      
               .std__pe44__lane17_strm1_cntl          ( std__pe44__lane17_strm1_cntl       ),      
               .std__pe44__lane17_strm1_data          ( std__pe44__lane17_strm1_data       ),      
               .std__pe44__lane17_strm1_data_valid    ( std__pe44__lane17_strm1_data_valid ),      
               .std__pe44__lane17_strm1_data_mask     ( std__pe44__lane17_strm1_data_mask  ),      

               // PE 44, Lane 18                 
               .pe44__std__lane18_strm0_ready         ( pe44__std__lane18_strm0_ready      ),      
               .std__pe44__lane18_strm0_cntl          ( std__pe44__lane18_strm0_cntl       ),      
               .std__pe44__lane18_strm0_data          ( std__pe44__lane18_strm0_data       ),      
               .std__pe44__lane18_strm0_data_valid    ( std__pe44__lane18_strm0_data_valid ),      
               .std__pe44__lane18_strm0_data_mask     ( std__pe44__lane18_strm0_data_mask  ),      

               .pe44__std__lane18_strm1_ready         ( pe44__std__lane18_strm1_ready      ),      
               .std__pe44__lane18_strm1_cntl          ( std__pe44__lane18_strm1_cntl       ),      
               .std__pe44__lane18_strm1_data          ( std__pe44__lane18_strm1_data       ),      
               .std__pe44__lane18_strm1_data_valid    ( std__pe44__lane18_strm1_data_valid ),      
               .std__pe44__lane18_strm1_data_mask     ( std__pe44__lane18_strm1_data_mask  ),      

               // PE 44, Lane 19                 
               .pe44__std__lane19_strm0_ready         ( pe44__std__lane19_strm0_ready      ),      
               .std__pe44__lane19_strm0_cntl          ( std__pe44__lane19_strm0_cntl       ),      
               .std__pe44__lane19_strm0_data          ( std__pe44__lane19_strm0_data       ),      
               .std__pe44__lane19_strm0_data_valid    ( std__pe44__lane19_strm0_data_valid ),      
               .std__pe44__lane19_strm0_data_mask     ( std__pe44__lane19_strm0_data_mask  ),      

               .pe44__std__lane19_strm1_ready         ( pe44__std__lane19_strm1_ready      ),      
               .std__pe44__lane19_strm1_cntl          ( std__pe44__lane19_strm1_cntl       ),      
               .std__pe44__lane19_strm1_data          ( std__pe44__lane19_strm1_data       ),      
               .std__pe44__lane19_strm1_data_valid    ( std__pe44__lane19_strm1_data_valid ),      
               .std__pe44__lane19_strm1_data_mask     ( std__pe44__lane19_strm1_data_mask  ),      

               // PE 44, Lane 20                 
               .pe44__std__lane20_strm0_ready         ( pe44__std__lane20_strm0_ready      ),      
               .std__pe44__lane20_strm0_cntl          ( std__pe44__lane20_strm0_cntl       ),      
               .std__pe44__lane20_strm0_data          ( std__pe44__lane20_strm0_data       ),      
               .std__pe44__lane20_strm0_data_valid    ( std__pe44__lane20_strm0_data_valid ),      
               .std__pe44__lane20_strm0_data_mask     ( std__pe44__lane20_strm0_data_mask  ),      

               .pe44__std__lane20_strm1_ready         ( pe44__std__lane20_strm1_ready      ),      
               .std__pe44__lane20_strm1_cntl          ( std__pe44__lane20_strm1_cntl       ),      
               .std__pe44__lane20_strm1_data          ( std__pe44__lane20_strm1_data       ),      
               .std__pe44__lane20_strm1_data_valid    ( std__pe44__lane20_strm1_data_valid ),      
               .std__pe44__lane20_strm1_data_mask     ( std__pe44__lane20_strm1_data_mask  ),      

               // PE 44, Lane 21                 
               .pe44__std__lane21_strm0_ready         ( pe44__std__lane21_strm0_ready      ),      
               .std__pe44__lane21_strm0_cntl          ( std__pe44__lane21_strm0_cntl       ),      
               .std__pe44__lane21_strm0_data          ( std__pe44__lane21_strm0_data       ),      
               .std__pe44__lane21_strm0_data_valid    ( std__pe44__lane21_strm0_data_valid ),      
               .std__pe44__lane21_strm0_data_mask     ( std__pe44__lane21_strm0_data_mask  ),      

               .pe44__std__lane21_strm1_ready         ( pe44__std__lane21_strm1_ready      ),      
               .std__pe44__lane21_strm1_cntl          ( std__pe44__lane21_strm1_cntl       ),      
               .std__pe44__lane21_strm1_data          ( std__pe44__lane21_strm1_data       ),      
               .std__pe44__lane21_strm1_data_valid    ( std__pe44__lane21_strm1_data_valid ),      
               .std__pe44__lane21_strm1_data_mask     ( std__pe44__lane21_strm1_data_mask  ),      

               // PE 44, Lane 22                 
               .pe44__std__lane22_strm0_ready         ( pe44__std__lane22_strm0_ready      ),      
               .std__pe44__lane22_strm0_cntl          ( std__pe44__lane22_strm0_cntl       ),      
               .std__pe44__lane22_strm0_data          ( std__pe44__lane22_strm0_data       ),      
               .std__pe44__lane22_strm0_data_valid    ( std__pe44__lane22_strm0_data_valid ),      
               .std__pe44__lane22_strm0_data_mask     ( std__pe44__lane22_strm0_data_mask  ),      

               .pe44__std__lane22_strm1_ready         ( pe44__std__lane22_strm1_ready      ),      
               .std__pe44__lane22_strm1_cntl          ( std__pe44__lane22_strm1_cntl       ),      
               .std__pe44__lane22_strm1_data          ( std__pe44__lane22_strm1_data       ),      
               .std__pe44__lane22_strm1_data_valid    ( std__pe44__lane22_strm1_data_valid ),      
               .std__pe44__lane22_strm1_data_mask     ( std__pe44__lane22_strm1_data_mask  ),      

               // PE 44, Lane 23                 
               .pe44__std__lane23_strm0_ready         ( pe44__std__lane23_strm0_ready      ),      
               .std__pe44__lane23_strm0_cntl          ( std__pe44__lane23_strm0_cntl       ),      
               .std__pe44__lane23_strm0_data          ( std__pe44__lane23_strm0_data       ),      
               .std__pe44__lane23_strm0_data_valid    ( std__pe44__lane23_strm0_data_valid ),      
               .std__pe44__lane23_strm0_data_mask     ( std__pe44__lane23_strm0_data_mask  ),      

               .pe44__std__lane23_strm1_ready         ( pe44__std__lane23_strm1_ready      ),      
               .std__pe44__lane23_strm1_cntl          ( std__pe44__lane23_strm1_cntl       ),      
               .std__pe44__lane23_strm1_data          ( std__pe44__lane23_strm1_data       ),      
               .std__pe44__lane23_strm1_data_valid    ( std__pe44__lane23_strm1_data_valid ),      
               .std__pe44__lane23_strm1_data_mask     ( std__pe44__lane23_strm1_data_mask  ),      

               // PE 44, Lane 24                 
               .pe44__std__lane24_strm0_ready         ( pe44__std__lane24_strm0_ready      ),      
               .std__pe44__lane24_strm0_cntl          ( std__pe44__lane24_strm0_cntl       ),      
               .std__pe44__lane24_strm0_data          ( std__pe44__lane24_strm0_data       ),      
               .std__pe44__lane24_strm0_data_valid    ( std__pe44__lane24_strm0_data_valid ),      
               .std__pe44__lane24_strm0_data_mask     ( std__pe44__lane24_strm0_data_mask  ),      

               .pe44__std__lane24_strm1_ready         ( pe44__std__lane24_strm1_ready      ),      
               .std__pe44__lane24_strm1_cntl          ( std__pe44__lane24_strm1_cntl       ),      
               .std__pe44__lane24_strm1_data          ( std__pe44__lane24_strm1_data       ),      
               .std__pe44__lane24_strm1_data_valid    ( std__pe44__lane24_strm1_data_valid ),      
               .std__pe44__lane24_strm1_data_mask     ( std__pe44__lane24_strm1_data_mask  ),      

               // PE 44, Lane 25                 
               .pe44__std__lane25_strm0_ready         ( pe44__std__lane25_strm0_ready      ),      
               .std__pe44__lane25_strm0_cntl          ( std__pe44__lane25_strm0_cntl       ),      
               .std__pe44__lane25_strm0_data          ( std__pe44__lane25_strm0_data       ),      
               .std__pe44__lane25_strm0_data_valid    ( std__pe44__lane25_strm0_data_valid ),      
               .std__pe44__lane25_strm0_data_mask     ( std__pe44__lane25_strm0_data_mask  ),      

               .pe44__std__lane25_strm1_ready         ( pe44__std__lane25_strm1_ready      ),      
               .std__pe44__lane25_strm1_cntl          ( std__pe44__lane25_strm1_cntl       ),      
               .std__pe44__lane25_strm1_data          ( std__pe44__lane25_strm1_data       ),      
               .std__pe44__lane25_strm1_data_valid    ( std__pe44__lane25_strm1_data_valid ),      
               .std__pe44__lane25_strm1_data_mask     ( std__pe44__lane25_strm1_data_mask  ),      

               // PE 44, Lane 26                 
               .pe44__std__lane26_strm0_ready         ( pe44__std__lane26_strm0_ready      ),      
               .std__pe44__lane26_strm0_cntl          ( std__pe44__lane26_strm0_cntl       ),      
               .std__pe44__lane26_strm0_data          ( std__pe44__lane26_strm0_data       ),      
               .std__pe44__lane26_strm0_data_valid    ( std__pe44__lane26_strm0_data_valid ),      
               .std__pe44__lane26_strm0_data_mask     ( std__pe44__lane26_strm0_data_mask  ),      

               .pe44__std__lane26_strm1_ready         ( pe44__std__lane26_strm1_ready      ),      
               .std__pe44__lane26_strm1_cntl          ( std__pe44__lane26_strm1_cntl       ),      
               .std__pe44__lane26_strm1_data          ( std__pe44__lane26_strm1_data       ),      
               .std__pe44__lane26_strm1_data_valid    ( std__pe44__lane26_strm1_data_valid ),      
               .std__pe44__lane26_strm1_data_mask     ( std__pe44__lane26_strm1_data_mask  ),      

               // PE 44, Lane 27                 
               .pe44__std__lane27_strm0_ready         ( pe44__std__lane27_strm0_ready      ),      
               .std__pe44__lane27_strm0_cntl          ( std__pe44__lane27_strm0_cntl       ),      
               .std__pe44__lane27_strm0_data          ( std__pe44__lane27_strm0_data       ),      
               .std__pe44__lane27_strm0_data_valid    ( std__pe44__lane27_strm0_data_valid ),      
               .std__pe44__lane27_strm0_data_mask     ( std__pe44__lane27_strm0_data_mask  ),      

               .pe44__std__lane27_strm1_ready         ( pe44__std__lane27_strm1_ready      ),      
               .std__pe44__lane27_strm1_cntl          ( std__pe44__lane27_strm1_cntl       ),      
               .std__pe44__lane27_strm1_data          ( std__pe44__lane27_strm1_data       ),      
               .std__pe44__lane27_strm1_data_valid    ( std__pe44__lane27_strm1_data_valid ),      
               .std__pe44__lane27_strm1_data_mask     ( std__pe44__lane27_strm1_data_mask  ),      

               // PE 44, Lane 28                 
               .pe44__std__lane28_strm0_ready         ( pe44__std__lane28_strm0_ready      ),      
               .std__pe44__lane28_strm0_cntl          ( std__pe44__lane28_strm0_cntl       ),      
               .std__pe44__lane28_strm0_data          ( std__pe44__lane28_strm0_data       ),      
               .std__pe44__lane28_strm0_data_valid    ( std__pe44__lane28_strm0_data_valid ),      
               .std__pe44__lane28_strm0_data_mask     ( std__pe44__lane28_strm0_data_mask  ),      

               .pe44__std__lane28_strm1_ready         ( pe44__std__lane28_strm1_ready      ),      
               .std__pe44__lane28_strm1_cntl          ( std__pe44__lane28_strm1_cntl       ),      
               .std__pe44__lane28_strm1_data          ( std__pe44__lane28_strm1_data       ),      
               .std__pe44__lane28_strm1_data_valid    ( std__pe44__lane28_strm1_data_valid ),      
               .std__pe44__lane28_strm1_data_mask     ( std__pe44__lane28_strm1_data_mask  ),      

               // PE 44, Lane 29                 
               .pe44__std__lane29_strm0_ready         ( pe44__std__lane29_strm0_ready      ),      
               .std__pe44__lane29_strm0_cntl          ( std__pe44__lane29_strm0_cntl       ),      
               .std__pe44__lane29_strm0_data          ( std__pe44__lane29_strm0_data       ),      
               .std__pe44__lane29_strm0_data_valid    ( std__pe44__lane29_strm0_data_valid ),      
               .std__pe44__lane29_strm0_data_mask     ( std__pe44__lane29_strm0_data_mask  ),      

               .pe44__std__lane29_strm1_ready         ( pe44__std__lane29_strm1_ready      ),      
               .std__pe44__lane29_strm1_cntl          ( std__pe44__lane29_strm1_cntl       ),      
               .std__pe44__lane29_strm1_data          ( std__pe44__lane29_strm1_data       ),      
               .std__pe44__lane29_strm1_data_valid    ( std__pe44__lane29_strm1_data_valid ),      
               .std__pe44__lane29_strm1_data_mask     ( std__pe44__lane29_strm1_data_mask  ),      

               // PE 44, Lane 30                 
               .pe44__std__lane30_strm0_ready         ( pe44__std__lane30_strm0_ready      ),      
               .std__pe44__lane30_strm0_cntl          ( std__pe44__lane30_strm0_cntl       ),      
               .std__pe44__lane30_strm0_data          ( std__pe44__lane30_strm0_data       ),      
               .std__pe44__lane30_strm0_data_valid    ( std__pe44__lane30_strm0_data_valid ),      
               .std__pe44__lane30_strm0_data_mask     ( std__pe44__lane30_strm0_data_mask  ),      

               .pe44__std__lane30_strm1_ready         ( pe44__std__lane30_strm1_ready      ),      
               .std__pe44__lane30_strm1_cntl          ( std__pe44__lane30_strm1_cntl       ),      
               .std__pe44__lane30_strm1_data          ( std__pe44__lane30_strm1_data       ),      
               .std__pe44__lane30_strm1_data_valid    ( std__pe44__lane30_strm1_data_valid ),      
               .std__pe44__lane30_strm1_data_mask     ( std__pe44__lane30_strm1_data_mask  ),      

               // PE 44, Lane 31                 
               .pe44__std__lane31_strm0_ready         ( pe44__std__lane31_strm0_ready      ),      
               .std__pe44__lane31_strm0_cntl          ( std__pe44__lane31_strm0_cntl       ),      
               .std__pe44__lane31_strm0_data          ( std__pe44__lane31_strm0_data       ),      
               .std__pe44__lane31_strm0_data_valid    ( std__pe44__lane31_strm0_data_valid ),      
               .std__pe44__lane31_strm0_data_mask     ( std__pe44__lane31_strm0_data_mask  ),      

               .pe44__std__lane31_strm1_ready         ( pe44__std__lane31_strm1_ready      ),      
               .std__pe44__lane31_strm1_cntl          ( std__pe44__lane31_strm1_cntl       ),      
               .std__pe44__lane31_strm1_data          ( std__pe44__lane31_strm1_data       ),      
               .std__pe44__lane31_strm1_data_valid    ( std__pe44__lane31_strm1_data_valid ),      
               .std__pe44__lane31_strm1_data_mask     ( std__pe44__lane31_strm1_data_mask  ),      

               // PE 45, Lane 0                 
               .pe45__std__lane0_strm0_ready         ( pe45__std__lane0_strm0_ready      ),      
               .std__pe45__lane0_strm0_cntl          ( std__pe45__lane0_strm0_cntl       ),      
               .std__pe45__lane0_strm0_data          ( std__pe45__lane0_strm0_data       ),      
               .std__pe45__lane0_strm0_data_valid    ( std__pe45__lane0_strm0_data_valid ),      
               .std__pe45__lane0_strm0_data_mask     ( std__pe45__lane0_strm0_data_mask  ),      

               .pe45__std__lane0_strm1_ready         ( pe45__std__lane0_strm1_ready      ),      
               .std__pe45__lane0_strm1_cntl          ( std__pe45__lane0_strm1_cntl       ),      
               .std__pe45__lane0_strm1_data          ( std__pe45__lane0_strm1_data       ),      
               .std__pe45__lane0_strm1_data_valid    ( std__pe45__lane0_strm1_data_valid ),      
               .std__pe45__lane0_strm1_data_mask     ( std__pe45__lane0_strm1_data_mask  ),      

               // PE 45, Lane 1                 
               .pe45__std__lane1_strm0_ready         ( pe45__std__lane1_strm0_ready      ),      
               .std__pe45__lane1_strm0_cntl          ( std__pe45__lane1_strm0_cntl       ),      
               .std__pe45__lane1_strm0_data          ( std__pe45__lane1_strm0_data       ),      
               .std__pe45__lane1_strm0_data_valid    ( std__pe45__lane1_strm0_data_valid ),      
               .std__pe45__lane1_strm0_data_mask     ( std__pe45__lane1_strm0_data_mask  ),      

               .pe45__std__lane1_strm1_ready         ( pe45__std__lane1_strm1_ready      ),      
               .std__pe45__lane1_strm1_cntl          ( std__pe45__lane1_strm1_cntl       ),      
               .std__pe45__lane1_strm1_data          ( std__pe45__lane1_strm1_data       ),      
               .std__pe45__lane1_strm1_data_valid    ( std__pe45__lane1_strm1_data_valid ),      
               .std__pe45__lane1_strm1_data_mask     ( std__pe45__lane1_strm1_data_mask  ),      

               // PE 45, Lane 2                 
               .pe45__std__lane2_strm0_ready         ( pe45__std__lane2_strm0_ready      ),      
               .std__pe45__lane2_strm0_cntl          ( std__pe45__lane2_strm0_cntl       ),      
               .std__pe45__lane2_strm0_data          ( std__pe45__lane2_strm0_data       ),      
               .std__pe45__lane2_strm0_data_valid    ( std__pe45__lane2_strm0_data_valid ),      
               .std__pe45__lane2_strm0_data_mask     ( std__pe45__lane2_strm0_data_mask  ),      

               .pe45__std__lane2_strm1_ready         ( pe45__std__lane2_strm1_ready      ),      
               .std__pe45__lane2_strm1_cntl          ( std__pe45__lane2_strm1_cntl       ),      
               .std__pe45__lane2_strm1_data          ( std__pe45__lane2_strm1_data       ),      
               .std__pe45__lane2_strm1_data_valid    ( std__pe45__lane2_strm1_data_valid ),      
               .std__pe45__lane2_strm1_data_mask     ( std__pe45__lane2_strm1_data_mask  ),      

               // PE 45, Lane 3                 
               .pe45__std__lane3_strm0_ready         ( pe45__std__lane3_strm0_ready      ),      
               .std__pe45__lane3_strm0_cntl          ( std__pe45__lane3_strm0_cntl       ),      
               .std__pe45__lane3_strm0_data          ( std__pe45__lane3_strm0_data       ),      
               .std__pe45__lane3_strm0_data_valid    ( std__pe45__lane3_strm0_data_valid ),      
               .std__pe45__lane3_strm0_data_mask     ( std__pe45__lane3_strm0_data_mask  ),      

               .pe45__std__lane3_strm1_ready         ( pe45__std__lane3_strm1_ready      ),      
               .std__pe45__lane3_strm1_cntl          ( std__pe45__lane3_strm1_cntl       ),      
               .std__pe45__lane3_strm1_data          ( std__pe45__lane3_strm1_data       ),      
               .std__pe45__lane3_strm1_data_valid    ( std__pe45__lane3_strm1_data_valid ),      
               .std__pe45__lane3_strm1_data_mask     ( std__pe45__lane3_strm1_data_mask  ),      

               // PE 45, Lane 4                 
               .pe45__std__lane4_strm0_ready         ( pe45__std__lane4_strm0_ready      ),      
               .std__pe45__lane4_strm0_cntl          ( std__pe45__lane4_strm0_cntl       ),      
               .std__pe45__lane4_strm0_data          ( std__pe45__lane4_strm0_data       ),      
               .std__pe45__lane4_strm0_data_valid    ( std__pe45__lane4_strm0_data_valid ),      
               .std__pe45__lane4_strm0_data_mask     ( std__pe45__lane4_strm0_data_mask  ),      

               .pe45__std__lane4_strm1_ready         ( pe45__std__lane4_strm1_ready      ),      
               .std__pe45__lane4_strm1_cntl          ( std__pe45__lane4_strm1_cntl       ),      
               .std__pe45__lane4_strm1_data          ( std__pe45__lane4_strm1_data       ),      
               .std__pe45__lane4_strm1_data_valid    ( std__pe45__lane4_strm1_data_valid ),      
               .std__pe45__lane4_strm1_data_mask     ( std__pe45__lane4_strm1_data_mask  ),      

               // PE 45, Lane 5                 
               .pe45__std__lane5_strm0_ready         ( pe45__std__lane5_strm0_ready      ),      
               .std__pe45__lane5_strm0_cntl          ( std__pe45__lane5_strm0_cntl       ),      
               .std__pe45__lane5_strm0_data          ( std__pe45__lane5_strm0_data       ),      
               .std__pe45__lane5_strm0_data_valid    ( std__pe45__lane5_strm0_data_valid ),      
               .std__pe45__lane5_strm0_data_mask     ( std__pe45__lane5_strm0_data_mask  ),      

               .pe45__std__lane5_strm1_ready         ( pe45__std__lane5_strm1_ready      ),      
               .std__pe45__lane5_strm1_cntl          ( std__pe45__lane5_strm1_cntl       ),      
               .std__pe45__lane5_strm1_data          ( std__pe45__lane5_strm1_data       ),      
               .std__pe45__lane5_strm1_data_valid    ( std__pe45__lane5_strm1_data_valid ),      
               .std__pe45__lane5_strm1_data_mask     ( std__pe45__lane5_strm1_data_mask  ),      

               // PE 45, Lane 6                 
               .pe45__std__lane6_strm0_ready         ( pe45__std__lane6_strm0_ready      ),      
               .std__pe45__lane6_strm0_cntl          ( std__pe45__lane6_strm0_cntl       ),      
               .std__pe45__lane6_strm0_data          ( std__pe45__lane6_strm0_data       ),      
               .std__pe45__lane6_strm0_data_valid    ( std__pe45__lane6_strm0_data_valid ),      
               .std__pe45__lane6_strm0_data_mask     ( std__pe45__lane6_strm0_data_mask  ),      

               .pe45__std__lane6_strm1_ready         ( pe45__std__lane6_strm1_ready      ),      
               .std__pe45__lane6_strm1_cntl          ( std__pe45__lane6_strm1_cntl       ),      
               .std__pe45__lane6_strm1_data          ( std__pe45__lane6_strm1_data       ),      
               .std__pe45__lane6_strm1_data_valid    ( std__pe45__lane6_strm1_data_valid ),      
               .std__pe45__lane6_strm1_data_mask     ( std__pe45__lane6_strm1_data_mask  ),      

               // PE 45, Lane 7                 
               .pe45__std__lane7_strm0_ready         ( pe45__std__lane7_strm0_ready      ),      
               .std__pe45__lane7_strm0_cntl          ( std__pe45__lane7_strm0_cntl       ),      
               .std__pe45__lane7_strm0_data          ( std__pe45__lane7_strm0_data       ),      
               .std__pe45__lane7_strm0_data_valid    ( std__pe45__lane7_strm0_data_valid ),      
               .std__pe45__lane7_strm0_data_mask     ( std__pe45__lane7_strm0_data_mask  ),      

               .pe45__std__lane7_strm1_ready         ( pe45__std__lane7_strm1_ready      ),      
               .std__pe45__lane7_strm1_cntl          ( std__pe45__lane7_strm1_cntl       ),      
               .std__pe45__lane7_strm1_data          ( std__pe45__lane7_strm1_data       ),      
               .std__pe45__lane7_strm1_data_valid    ( std__pe45__lane7_strm1_data_valid ),      
               .std__pe45__lane7_strm1_data_mask     ( std__pe45__lane7_strm1_data_mask  ),      

               // PE 45, Lane 8                 
               .pe45__std__lane8_strm0_ready         ( pe45__std__lane8_strm0_ready      ),      
               .std__pe45__lane8_strm0_cntl          ( std__pe45__lane8_strm0_cntl       ),      
               .std__pe45__lane8_strm0_data          ( std__pe45__lane8_strm0_data       ),      
               .std__pe45__lane8_strm0_data_valid    ( std__pe45__lane8_strm0_data_valid ),      
               .std__pe45__lane8_strm0_data_mask     ( std__pe45__lane8_strm0_data_mask  ),      

               .pe45__std__lane8_strm1_ready         ( pe45__std__lane8_strm1_ready      ),      
               .std__pe45__lane8_strm1_cntl          ( std__pe45__lane8_strm1_cntl       ),      
               .std__pe45__lane8_strm1_data          ( std__pe45__lane8_strm1_data       ),      
               .std__pe45__lane8_strm1_data_valid    ( std__pe45__lane8_strm1_data_valid ),      
               .std__pe45__lane8_strm1_data_mask     ( std__pe45__lane8_strm1_data_mask  ),      

               // PE 45, Lane 9                 
               .pe45__std__lane9_strm0_ready         ( pe45__std__lane9_strm0_ready      ),      
               .std__pe45__lane9_strm0_cntl          ( std__pe45__lane9_strm0_cntl       ),      
               .std__pe45__lane9_strm0_data          ( std__pe45__lane9_strm0_data       ),      
               .std__pe45__lane9_strm0_data_valid    ( std__pe45__lane9_strm0_data_valid ),      
               .std__pe45__lane9_strm0_data_mask     ( std__pe45__lane9_strm0_data_mask  ),      

               .pe45__std__lane9_strm1_ready         ( pe45__std__lane9_strm1_ready      ),      
               .std__pe45__lane9_strm1_cntl          ( std__pe45__lane9_strm1_cntl       ),      
               .std__pe45__lane9_strm1_data          ( std__pe45__lane9_strm1_data       ),      
               .std__pe45__lane9_strm1_data_valid    ( std__pe45__lane9_strm1_data_valid ),      
               .std__pe45__lane9_strm1_data_mask     ( std__pe45__lane9_strm1_data_mask  ),      

               // PE 45, Lane 10                 
               .pe45__std__lane10_strm0_ready         ( pe45__std__lane10_strm0_ready      ),      
               .std__pe45__lane10_strm0_cntl          ( std__pe45__lane10_strm0_cntl       ),      
               .std__pe45__lane10_strm0_data          ( std__pe45__lane10_strm0_data       ),      
               .std__pe45__lane10_strm0_data_valid    ( std__pe45__lane10_strm0_data_valid ),      
               .std__pe45__lane10_strm0_data_mask     ( std__pe45__lane10_strm0_data_mask  ),      

               .pe45__std__lane10_strm1_ready         ( pe45__std__lane10_strm1_ready      ),      
               .std__pe45__lane10_strm1_cntl          ( std__pe45__lane10_strm1_cntl       ),      
               .std__pe45__lane10_strm1_data          ( std__pe45__lane10_strm1_data       ),      
               .std__pe45__lane10_strm1_data_valid    ( std__pe45__lane10_strm1_data_valid ),      
               .std__pe45__lane10_strm1_data_mask     ( std__pe45__lane10_strm1_data_mask  ),      

               // PE 45, Lane 11                 
               .pe45__std__lane11_strm0_ready         ( pe45__std__lane11_strm0_ready      ),      
               .std__pe45__lane11_strm0_cntl          ( std__pe45__lane11_strm0_cntl       ),      
               .std__pe45__lane11_strm0_data          ( std__pe45__lane11_strm0_data       ),      
               .std__pe45__lane11_strm0_data_valid    ( std__pe45__lane11_strm0_data_valid ),      
               .std__pe45__lane11_strm0_data_mask     ( std__pe45__lane11_strm0_data_mask  ),      

               .pe45__std__lane11_strm1_ready         ( pe45__std__lane11_strm1_ready      ),      
               .std__pe45__lane11_strm1_cntl          ( std__pe45__lane11_strm1_cntl       ),      
               .std__pe45__lane11_strm1_data          ( std__pe45__lane11_strm1_data       ),      
               .std__pe45__lane11_strm1_data_valid    ( std__pe45__lane11_strm1_data_valid ),      
               .std__pe45__lane11_strm1_data_mask     ( std__pe45__lane11_strm1_data_mask  ),      

               // PE 45, Lane 12                 
               .pe45__std__lane12_strm0_ready         ( pe45__std__lane12_strm0_ready      ),      
               .std__pe45__lane12_strm0_cntl          ( std__pe45__lane12_strm0_cntl       ),      
               .std__pe45__lane12_strm0_data          ( std__pe45__lane12_strm0_data       ),      
               .std__pe45__lane12_strm0_data_valid    ( std__pe45__lane12_strm0_data_valid ),      
               .std__pe45__lane12_strm0_data_mask     ( std__pe45__lane12_strm0_data_mask  ),      

               .pe45__std__lane12_strm1_ready         ( pe45__std__lane12_strm1_ready      ),      
               .std__pe45__lane12_strm1_cntl          ( std__pe45__lane12_strm1_cntl       ),      
               .std__pe45__lane12_strm1_data          ( std__pe45__lane12_strm1_data       ),      
               .std__pe45__lane12_strm1_data_valid    ( std__pe45__lane12_strm1_data_valid ),      
               .std__pe45__lane12_strm1_data_mask     ( std__pe45__lane12_strm1_data_mask  ),      

               // PE 45, Lane 13                 
               .pe45__std__lane13_strm0_ready         ( pe45__std__lane13_strm0_ready      ),      
               .std__pe45__lane13_strm0_cntl          ( std__pe45__lane13_strm0_cntl       ),      
               .std__pe45__lane13_strm0_data          ( std__pe45__lane13_strm0_data       ),      
               .std__pe45__lane13_strm0_data_valid    ( std__pe45__lane13_strm0_data_valid ),      
               .std__pe45__lane13_strm0_data_mask     ( std__pe45__lane13_strm0_data_mask  ),      

               .pe45__std__lane13_strm1_ready         ( pe45__std__lane13_strm1_ready      ),      
               .std__pe45__lane13_strm1_cntl          ( std__pe45__lane13_strm1_cntl       ),      
               .std__pe45__lane13_strm1_data          ( std__pe45__lane13_strm1_data       ),      
               .std__pe45__lane13_strm1_data_valid    ( std__pe45__lane13_strm1_data_valid ),      
               .std__pe45__lane13_strm1_data_mask     ( std__pe45__lane13_strm1_data_mask  ),      

               // PE 45, Lane 14                 
               .pe45__std__lane14_strm0_ready         ( pe45__std__lane14_strm0_ready      ),      
               .std__pe45__lane14_strm0_cntl          ( std__pe45__lane14_strm0_cntl       ),      
               .std__pe45__lane14_strm0_data          ( std__pe45__lane14_strm0_data       ),      
               .std__pe45__lane14_strm0_data_valid    ( std__pe45__lane14_strm0_data_valid ),      
               .std__pe45__lane14_strm0_data_mask     ( std__pe45__lane14_strm0_data_mask  ),      

               .pe45__std__lane14_strm1_ready         ( pe45__std__lane14_strm1_ready      ),      
               .std__pe45__lane14_strm1_cntl          ( std__pe45__lane14_strm1_cntl       ),      
               .std__pe45__lane14_strm1_data          ( std__pe45__lane14_strm1_data       ),      
               .std__pe45__lane14_strm1_data_valid    ( std__pe45__lane14_strm1_data_valid ),      
               .std__pe45__lane14_strm1_data_mask     ( std__pe45__lane14_strm1_data_mask  ),      

               // PE 45, Lane 15                 
               .pe45__std__lane15_strm0_ready         ( pe45__std__lane15_strm0_ready      ),      
               .std__pe45__lane15_strm0_cntl          ( std__pe45__lane15_strm0_cntl       ),      
               .std__pe45__lane15_strm0_data          ( std__pe45__lane15_strm0_data       ),      
               .std__pe45__lane15_strm0_data_valid    ( std__pe45__lane15_strm0_data_valid ),      
               .std__pe45__lane15_strm0_data_mask     ( std__pe45__lane15_strm0_data_mask  ),      

               .pe45__std__lane15_strm1_ready         ( pe45__std__lane15_strm1_ready      ),      
               .std__pe45__lane15_strm1_cntl          ( std__pe45__lane15_strm1_cntl       ),      
               .std__pe45__lane15_strm1_data          ( std__pe45__lane15_strm1_data       ),      
               .std__pe45__lane15_strm1_data_valid    ( std__pe45__lane15_strm1_data_valid ),      
               .std__pe45__lane15_strm1_data_mask     ( std__pe45__lane15_strm1_data_mask  ),      

               // PE 45, Lane 16                 
               .pe45__std__lane16_strm0_ready         ( pe45__std__lane16_strm0_ready      ),      
               .std__pe45__lane16_strm0_cntl          ( std__pe45__lane16_strm0_cntl       ),      
               .std__pe45__lane16_strm0_data          ( std__pe45__lane16_strm0_data       ),      
               .std__pe45__lane16_strm0_data_valid    ( std__pe45__lane16_strm0_data_valid ),      
               .std__pe45__lane16_strm0_data_mask     ( std__pe45__lane16_strm0_data_mask  ),      

               .pe45__std__lane16_strm1_ready         ( pe45__std__lane16_strm1_ready      ),      
               .std__pe45__lane16_strm1_cntl          ( std__pe45__lane16_strm1_cntl       ),      
               .std__pe45__lane16_strm1_data          ( std__pe45__lane16_strm1_data       ),      
               .std__pe45__lane16_strm1_data_valid    ( std__pe45__lane16_strm1_data_valid ),      
               .std__pe45__lane16_strm1_data_mask     ( std__pe45__lane16_strm1_data_mask  ),      

               // PE 45, Lane 17                 
               .pe45__std__lane17_strm0_ready         ( pe45__std__lane17_strm0_ready      ),      
               .std__pe45__lane17_strm0_cntl          ( std__pe45__lane17_strm0_cntl       ),      
               .std__pe45__lane17_strm0_data          ( std__pe45__lane17_strm0_data       ),      
               .std__pe45__lane17_strm0_data_valid    ( std__pe45__lane17_strm0_data_valid ),      
               .std__pe45__lane17_strm0_data_mask     ( std__pe45__lane17_strm0_data_mask  ),      

               .pe45__std__lane17_strm1_ready         ( pe45__std__lane17_strm1_ready      ),      
               .std__pe45__lane17_strm1_cntl          ( std__pe45__lane17_strm1_cntl       ),      
               .std__pe45__lane17_strm1_data          ( std__pe45__lane17_strm1_data       ),      
               .std__pe45__lane17_strm1_data_valid    ( std__pe45__lane17_strm1_data_valid ),      
               .std__pe45__lane17_strm1_data_mask     ( std__pe45__lane17_strm1_data_mask  ),      

               // PE 45, Lane 18                 
               .pe45__std__lane18_strm0_ready         ( pe45__std__lane18_strm0_ready      ),      
               .std__pe45__lane18_strm0_cntl          ( std__pe45__lane18_strm0_cntl       ),      
               .std__pe45__lane18_strm0_data          ( std__pe45__lane18_strm0_data       ),      
               .std__pe45__lane18_strm0_data_valid    ( std__pe45__lane18_strm0_data_valid ),      
               .std__pe45__lane18_strm0_data_mask     ( std__pe45__lane18_strm0_data_mask  ),      

               .pe45__std__lane18_strm1_ready         ( pe45__std__lane18_strm1_ready      ),      
               .std__pe45__lane18_strm1_cntl          ( std__pe45__lane18_strm1_cntl       ),      
               .std__pe45__lane18_strm1_data          ( std__pe45__lane18_strm1_data       ),      
               .std__pe45__lane18_strm1_data_valid    ( std__pe45__lane18_strm1_data_valid ),      
               .std__pe45__lane18_strm1_data_mask     ( std__pe45__lane18_strm1_data_mask  ),      

               // PE 45, Lane 19                 
               .pe45__std__lane19_strm0_ready         ( pe45__std__lane19_strm0_ready      ),      
               .std__pe45__lane19_strm0_cntl          ( std__pe45__lane19_strm0_cntl       ),      
               .std__pe45__lane19_strm0_data          ( std__pe45__lane19_strm0_data       ),      
               .std__pe45__lane19_strm0_data_valid    ( std__pe45__lane19_strm0_data_valid ),      
               .std__pe45__lane19_strm0_data_mask     ( std__pe45__lane19_strm0_data_mask  ),      

               .pe45__std__lane19_strm1_ready         ( pe45__std__lane19_strm1_ready      ),      
               .std__pe45__lane19_strm1_cntl          ( std__pe45__lane19_strm1_cntl       ),      
               .std__pe45__lane19_strm1_data          ( std__pe45__lane19_strm1_data       ),      
               .std__pe45__lane19_strm1_data_valid    ( std__pe45__lane19_strm1_data_valid ),      
               .std__pe45__lane19_strm1_data_mask     ( std__pe45__lane19_strm1_data_mask  ),      

               // PE 45, Lane 20                 
               .pe45__std__lane20_strm0_ready         ( pe45__std__lane20_strm0_ready      ),      
               .std__pe45__lane20_strm0_cntl          ( std__pe45__lane20_strm0_cntl       ),      
               .std__pe45__lane20_strm0_data          ( std__pe45__lane20_strm0_data       ),      
               .std__pe45__lane20_strm0_data_valid    ( std__pe45__lane20_strm0_data_valid ),      
               .std__pe45__lane20_strm0_data_mask     ( std__pe45__lane20_strm0_data_mask  ),      

               .pe45__std__lane20_strm1_ready         ( pe45__std__lane20_strm1_ready      ),      
               .std__pe45__lane20_strm1_cntl          ( std__pe45__lane20_strm1_cntl       ),      
               .std__pe45__lane20_strm1_data          ( std__pe45__lane20_strm1_data       ),      
               .std__pe45__lane20_strm1_data_valid    ( std__pe45__lane20_strm1_data_valid ),      
               .std__pe45__lane20_strm1_data_mask     ( std__pe45__lane20_strm1_data_mask  ),      

               // PE 45, Lane 21                 
               .pe45__std__lane21_strm0_ready         ( pe45__std__lane21_strm0_ready      ),      
               .std__pe45__lane21_strm0_cntl          ( std__pe45__lane21_strm0_cntl       ),      
               .std__pe45__lane21_strm0_data          ( std__pe45__lane21_strm0_data       ),      
               .std__pe45__lane21_strm0_data_valid    ( std__pe45__lane21_strm0_data_valid ),      
               .std__pe45__lane21_strm0_data_mask     ( std__pe45__lane21_strm0_data_mask  ),      

               .pe45__std__lane21_strm1_ready         ( pe45__std__lane21_strm1_ready      ),      
               .std__pe45__lane21_strm1_cntl          ( std__pe45__lane21_strm1_cntl       ),      
               .std__pe45__lane21_strm1_data          ( std__pe45__lane21_strm1_data       ),      
               .std__pe45__lane21_strm1_data_valid    ( std__pe45__lane21_strm1_data_valid ),      
               .std__pe45__lane21_strm1_data_mask     ( std__pe45__lane21_strm1_data_mask  ),      

               // PE 45, Lane 22                 
               .pe45__std__lane22_strm0_ready         ( pe45__std__lane22_strm0_ready      ),      
               .std__pe45__lane22_strm0_cntl          ( std__pe45__lane22_strm0_cntl       ),      
               .std__pe45__lane22_strm0_data          ( std__pe45__lane22_strm0_data       ),      
               .std__pe45__lane22_strm0_data_valid    ( std__pe45__lane22_strm0_data_valid ),      
               .std__pe45__lane22_strm0_data_mask     ( std__pe45__lane22_strm0_data_mask  ),      

               .pe45__std__lane22_strm1_ready         ( pe45__std__lane22_strm1_ready      ),      
               .std__pe45__lane22_strm1_cntl          ( std__pe45__lane22_strm1_cntl       ),      
               .std__pe45__lane22_strm1_data          ( std__pe45__lane22_strm1_data       ),      
               .std__pe45__lane22_strm1_data_valid    ( std__pe45__lane22_strm1_data_valid ),      
               .std__pe45__lane22_strm1_data_mask     ( std__pe45__lane22_strm1_data_mask  ),      

               // PE 45, Lane 23                 
               .pe45__std__lane23_strm0_ready         ( pe45__std__lane23_strm0_ready      ),      
               .std__pe45__lane23_strm0_cntl          ( std__pe45__lane23_strm0_cntl       ),      
               .std__pe45__lane23_strm0_data          ( std__pe45__lane23_strm0_data       ),      
               .std__pe45__lane23_strm0_data_valid    ( std__pe45__lane23_strm0_data_valid ),      
               .std__pe45__lane23_strm0_data_mask     ( std__pe45__lane23_strm0_data_mask  ),      

               .pe45__std__lane23_strm1_ready         ( pe45__std__lane23_strm1_ready      ),      
               .std__pe45__lane23_strm1_cntl          ( std__pe45__lane23_strm1_cntl       ),      
               .std__pe45__lane23_strm1_data          ( std__pe45__lane23_strm1_data       ),      
               .std__pe45__lane23_strm1_data_valid    ( std__pe45__lane23_strm1_data_valid ),      
               .std__pe45__lane23_strm1_data_mask     ( std__pe45__lane23_strm1_data_mask  ),      

               // PE 45, Lane 24                 
               .pe45__std__lane24_strm0_ready         ( pe45__std__lane24_strm0_ready      ),      
               .std__pe45__lane24_strm0_cntl          ( std__pe45__lane24_strm0_cntl       ),      
               .std__pe45__lane24_strm0_data          ( std__pe45__lane24_strm0_data       ),      
               .std__pe45__lane24_strm0_data_valid    ( std__pe45__lane24_strm0_data_valid ),      
               .std__pe45__lane24_strm0_data_mask     ( std__pe45__lane24_strm0_data_mask  ),      

               .pe45__std__lane24_strm1_ready         ( pe45__std__lane24_strm1_ready      ),      
               .std__pe45__lane24_strm1_cntl          ( std__pe45__lane24_strm1_cntl       ),      
               .std__pe45__lane24_strm1_data          ( std__pe45__lane24_strm1_data       ),      
               .std__pe45__lane24_strm1_data_valid    ( std__pe45__lane24_strm1_data_valid ),      
               .std__pe45__lane24_strm1_data_mask     ( std__pe45__lane24_strm1_data_mask  ),      

               // PE 45, Lane 25                 
               .pe45__std__lane25_strm0_ready         ( pe45__std__lane25_strm0_ready      ),      
               .std__pe45__lane25_strm0_cntl          ( std__pe45__lane25_strm0_cntl       ),      
               .std__pe45__lane25_strm0_data          ( std__pe45__lane25_strm0_data       ),      
               .std__pe45__lane25_strm0_data_valid    ( std__pe45__lane25_strm0_data_valid ),      
               .std__pe45__lane25_strm0_data_mask     ( std__pe45__lane25_strm0_data_mask  ),      

               .pe45__std__lane25_strm1_ready         ( pe45__std__lane25_strm1_ready      ),      
               .std__pe45__lane25_strm1_cntl          ( std__pe45__lane25_strm1_cntl       ),      
               .std__pe45__lane25_strm1_data          ( std__pe45__lane25_strm1_data       ),      
               .std__pe45__lane25_strm1_data_valid    ( std__pe45__lane25_strm1_data_valid ),      
               .std__pe45__lane25_strm1_data_mask     ( std__pe45__lane25_strm1_data_mask  ),      

               // PE 45, Lane 26                 
               .pe45__std__lane26_strm0_ready         ( pe45__std__lane26_strm0_ready      ),      
               .std__pe45__lane26_strm0_cntl          ( std__pe45__lane26_strm0_cntl       ),      
               .std__pe45__lane26_strm0_data          ( std__pe45__lane26_strm0_data       ),      
               .std__pe45__lane26_strm0_data_valid    ( std__pe45__lane26_strm0_data_valid ),      
               .std__pe45__lane26_strm0_data_mask     ( std__pe45__lane26_strm0_data_mask  ),      

               .pe45__std__lane26_strm1_ready         ( pe45__std__lane26_strm1_ready      ),      
               .std__pe45__lane26_strm1_cntl          ( std__pe45__lane26_strm1_cntl       ),      
               .std__pe45__lane26_strm1_data          ( std__pe45__lane26_strm1_data       ),      
               .std__pe45__lane26_strm1_data_valid    ( std__pe45__lane26_strm1_data_valid ),      
               .std__pe45__lane26_strm1_data_mask     ( std__pe45__lane26_strm1_data_mask  ),      

               // PE 45, Lane 27                 
               .pe45__std__lane27_strm0_ready         ( pe45__std__lane27_strm0_ready      ),      
               .std__pe45__lane27_strm0_cntl          ( std__pe45__lane27_strm0_cntl       ),      
               .std__pe45__lane27_strm0_data          ( std__pe45__lane27_strm0_data       ),      
               .std__pe45__lane27_strm0_data_valid    ( std__pe45__lane27_strm0_data_valid ),      
               .std__pe45__lane27_strm0_data_mask     ( std__pe45__lane27_strm0_data_mask  ),      

               .pe45__std__lane27_strm1_ready         ( pe45__std__lane27_strm1_ready      ),      
               .std__pe45__lane27_strm1_cntl          ( std__pe45__lane27_strm1_cntl       ),      
               .std__pe45__lane27_strm1_data          ( std__pe45__lane27_strm1_data       ),      
               .std__pe45__lane27_strm1_data_valid    ( std__pe45__lane27_strm1_data_valid ),      
               .std__pe45__lane27_strm1_data_mask     ( std__pe45__lane27_strm1_data_mask  ),      

               // PE 45, Lane 28                 
               .pe45__std__lane28_strm0_ready         ( pe45__std__lane28_strm0_ready      ),      
               .std__pe45__lane28_strm0_cntl          ( std__pe45__lane28_strm0_cntl       ),      
               .std__pe45__lane28_strm0_data          ( std__pe45__lane28_strm0_data       ),      
               .std__pe45__lane28_strm0_data_valid    ( std__pe45__lane28_strm0_data_valid ),      
               .std__pe45__lane28_strm0_data_mask     ( std__pe45__lane28_strm0_data_mask  ),      

               .pe45__std__lane28_strm1_ready         ( pe45__std__lane28_strm1_ready      ),      
               .std__pe45__lane28_strm1_cntl          ( std__pe45__lane28_strm1_cntl       ),      
               .std__pe45__lane28_strm1_data          ( std__pe45__lane28_strm1_data       ),      
               .std__pe45__lane28_strm1_data_valid    ( std__pe45__lane28_strm1_data_valid ),      
               .std__pe45__lane28_strm1_data_mask     ( std__pe45__lane28_strm1_data_mask  ),      

               // PE 45, Lane 29                 
               .pe45__std__lane29_strm0_ready         ( pe45__std__lane29_strm0_ready      ),      
               .std__pe45__lane29_strm0_cntl          ( std__pe45__lane29_strm0_cntl       ),      
               .std__pe45__lane29_strm0_data          ( std__pe45__lane29_strm0_data       ),      
               .std__pe45__lane29_strm0_data_valid    ( std__pe45__lane29_strm0_data_valid ),      
               .std__pe45__lane29_strm0_data_mask     ( std__pe45__lane29_strm0_data_mask  ),      

               .pe45__std__lane29_strm1_ready         ( pe45__std__lane29_strm1_ready      ),      
               .std__pe45__lane29_strm1_cntl          ( std__pe45__lane29_strm1_cntl       ),      
               .std__pe45__lane29_strm1_data          ( std__pe45__lane29_strm1_data       ),      
               .std__pe45__lane29_strm1_data_valid    ( std__pe45__lane29_strm1_data_valid ),      
               .std__pe45__lane29_strm1_data_mask     ( std__pe45__lane29_strm1_data_mask  ),      

               // PE 45, Lane 30                 
               .pe45__std__lane30_strm0_ready         ( pe45__std__lane30_strm0_ready      ),      
               .std__pe45__lane30_strm0_cntl          ( std__pe45__lane30_strm0_cntl       ),      
               .std__pe45__lane30_strm0_data          ( std__pe45__lane30_strm0_data       ),      
               .std__pe45__lane30_strm0_data_valid    ( std__pe45__lane30_strm0_data_valid ),      
               .std__pe45__lane30_strm0_data_mask     ( std__pe45__lane30_strm0_data_mask  ),      

               .pe45__std__lane30_strm1_ready         ( pe45__std__lane30_strm1_ready      ),      
               .std__pe45__lane30_strm1_cntl          ( std__pe45__lane30_strm1_cntl       ),      
               .std__pe45__lane30_strm1_data          ( std__pe45__lane30_strm1_data       ),      
               .std__pe45__lane30_strm1_data_valid    ( std__pe45__lane30_strm1_data_valid ),      
               .std__pe45__lane30_strm1_data_mask     ( std__pe45__lane30_strm1_data_mask  ),      

               // PE 45, Lane 31                 
               .pe45__std__lane31_strm0_ready         ( pe45__std__lane31_strm0_ready      ),      
               .std__pe45__lane31_strm0_cntl          ( std__pe45__lane31_strm0_cntl       ),      
               .std__pe45__lane31_strm0_data          ( std__pe45__lane31_strm0_data       ),      
               .std__pe45__lane31_strm0_data_valid    ( std__pe45__lane31_strm0_data_valid ),      
               .std__pe45__lane31_strm0_data_mask     ( std__pe45__lane31_strm0_data_mask  ),      

               .pe45__std__lane31_strm1_ready         ( pe45__std__lane31_strm1_ready      ),      
               .std__pe45__lane31_strm1_cntl          ( std__pe45__lane31_strm1_cntl       ),      
               .std__pe45__lane31_strm1_data          ( std__pe45__lane31_strm1_data       ),      
               .std__pe45__lane31_strm1_data_valid    ( std__pe45__lane31_strm1_data_valid ),      
               .std__pe45__lane31_strm1_data_mask     ( std__pe45__lane31_strm1_data_mask  ),      

               // PE 46, Lane 0                 
               .pe46__std__lane0_strm0_ready         ( pe46__std__lane0_strm0_ready      ),      
               .std__pe46__lane0_strm0_cntl          ( std__pe46__lane0_strm0_cntl       ),      
               .std__pe46__lane0_strm0_data          ( std__pe46__lane0_strm0_data       ),      
               .std__pe46__lane0_strm0_data_valid    ( std__pe46__lane0_strm0_data_valid ),      
               .std__pe46__lane0_strm0_data_mask     ( std__pe46__lane0_strm0_data_mask  ),      

               .pe46__std__lane0_strm1_ready         ( pe46__std__lane0_strm1_ready      ),      
               .std__pe46__lane0_strm1_cntl          ( std__pe46__lane0_strm1_cntl       ),      
               .std__pe46__lane0_strm1_data          ( std__pe46__lane0_strm1_data       ),      
               .std__pe46__lane0_strm1_data_valid    ( std__pe46__lane0_strm1_data_valid ),      
               .std__pe46__lane0_strm1_data_mask     ( std__pe46__lane0_strm1_data_mask  ),      

               // PE 46, Lane 1                 
               .pe46__std__lane1_strm0_ready         ( pe46__std__lane1_strm0_ready      ),      
               .std__pe46__lane1_strm0_cntl          ( std__pe46__lane1_strm0_cntl       ),      
               .std__pe46__lane1_strm0_data          ( std__pe46__lane1_strm0_data       ),      
               .std__pe46__lane1_strm0_data_valid    ( std__pe46__lane1_strm0_data_valid ),      
               .std__pe46__lane1_strm0_data_mask     ( std__pe46__lane1_strm0_data_mask  ),      

               .pe46__std__lane1_strm1_ready         ( pe46__std__lane1_strm1_ready      ),      
               .std__pe46__lane1_strm1_cntl          ( std__pe46__lane1_strm1_cntl       ),      
               .std__pe46__lane1_strm1_data          ( std__pe46__lane1_strm1_data       ),      
               .std__pe46__lane1_strm1_data_valid    ( std__pe46__lane1_strm1_data_valid ),      
               .std__pe46__lane1_strm1_data_mask     ( std__pe46__lane1_strm1_data_mask  ),      

               // PE 46, Lane 2                 
               .pe46__std__lane2_strm0_ready         ( pe46__std__lane2_strm0_ready      ),      
               .std__pe46__lane2_strm0_cntl          ( std__pe46__lane2_strm0_cntl       ),      
               .std__pe46__lane2_strm0_data          ( std__pe46__lane2_strm0_data       ),      
               .std__pe46__lane2_strm0_data_valid    ( std__pe46__lane2_strm0_data_valid ),      
               .std__pe46__lane2_strm0_data_mask     ( std__pe46__lane2_strm0_data_mask  ),      

               .pe46__std__lane2_strm1_ready         ( pe46__std__lane2_strm1_ready      ),      
               .std__pe46__lane2_strm1_cntl          ( std__pe46__lane2_strm1_cntl       ),      
               .std__pe46__lane2_strm1_data          ( std__pe46__lane2_strm1_data       ),      
               .std__pe46__lane2_strm1_data_valid    ( std__pe46__lane2_strm1_data_valid ),      
               .std__pe46__lane2_strm1_data_mask     ( std__pe46__lane2_strm1_data_mask  ),      

               // PE 46, Lane 3                 
               .pe46__std__lane3_strm0_ready         ( pe46__std__lane3_strm0_ready      ),      
               .std__pe46__lane3_strm0_cntl          ( std__pe46__lane3_strm0_cntl       ),      
               .std__pe46__lane3_strm0_data          ( std__pe46__lane3_strm0_data       ),      
               .std__pe46__lane3_strm0_data_valid    ( std__pe46__lane3_strm0_data_valid ),      
               .std__pe46__lane3_strm0_data_mask     ( std__pe46__lane3_strm0_data_mask  ),      

               .pe46__std__lane3_strm1_ready         ( pe46__std__lane3_strm1_ready      ),      
               .std__pe46__lane3_strm1_cntl          ( std__pe46__lane3_strm1_cntl       ),      
               .std__pe46__lane3_strm1_data          ( std__pe46__lane3_strm1_data       ),      
               .std__pe46__lane3_strm1_data_valid    ( std__pe46__lane3_strm1_data_valid ),      
               .std__pe46__lane3_strm1_data_mask     ( std__pe46__lane3_strm1_data_mask  ),      

               // PE 46, Lane 4                 
               .pe46__std__lane4_strm0_ready         ( pe46__std__lane4_strm0_ready      ),      
               .std__pe46__lane4_strm0_cntl          ( std__pe46__lane4_strm0_cntl       ),      
               .std__pe46__lane4_strm0_data          ( std__pe46__lane4_strm0_data       ),      
               .std__pe46__lane4_strm0_data_valid    ( std__pe46__lane4_strm0_data_valid ),      
               .std__pe46__lane4_strm0_data_mask     ( std__pe46__lane4_strm0_data_mask  ),      

               .pe46__std__lane4_strm1_ready         ( pe46__std__lane4_strm1_ready      ),      
               .std__pe46__lane4_strm1_cntl          ( std__pe46__lane4_strm1_cntl       ),      
               .std__pe46__lane4_strm1_data          ( std__pe46__lane4_strm1_data       ),      
               .std__pe46__lane4_strm1_data_valid    ( std__pe46__lane4_strm1_data_valid ),      
               .std__pe46__lane4_strm1_data_mask     ( std__pe46__lane4_strm1_data_mask  ),      

               // PE 46, Lane 5                 
               .pe46__std__lane5_strm0_ready         ( pe46__std__lane5_strm0_ready      ),      
               .std__pe46__lane5_strm0_cntl          ( std__pe46__lane5_strm0_cntl       ),      
               .std__pe46__lane5_strm0_data          ( std__pe46__lane5_strm0_data       ),      
               .std__pe46__lane5_strm0_data_valid    ( std__pe46__lane5_strm0_data_valid ),      
               .std__pe46__lane5_strm0_data_mask     ( std__pe46__lane5_strm0_data_mask  ),      

               .pe46__std__lane5_strm1_ready         ( pe46__std__lane5_strm1_ready      ),      
               .std__pe46__lane5_strm1_cntl          ( std__pe46__lane5_strm1_cntl       ),      
               .std__pe46__lane5_strm1_data          ( std__pe46__lane5_strm1_data       ),      
               .std__pe46__lane5_strm1_data_valid    ( std__pe46__lane5_strm1_data_valid ),      
               .std__pe46__lane5_strm1_data_mask     ( std__pe46__lane5_strm1_data_mask  ),      

               // PE 46, Lane 6                 
               .pe46__std__lane6_strm0_ready         ( pe46__std__lane6_strm0_ready      ),      
               .std__pe46__lane6_strm0_cntl          ( std__pe46__lane6_strm0_cntl       ),      
               .std__pe46__lane6_strm0_data          ( std__pe46__lane6_strm0_data       ),      
               .std__pe46__lane6_strm0_data_valid    ( std__pe46__lane6_strm0_data_valid ),      
               .std__pe46__lane6_strm0_data_mask     ( std__pe46__lane6_strm0_data_mask  ),      

               .pe46__std__lane6_strm1_ready         ( pe46__std__lane6_strm1_ready      ),      
               .std__pe46__lane6_strm1_cntl          ( std__pe46__lane6_strm1_cntl       ),      
               .std__pe46__lane6_strm1_data          ( std__pe46__lane6_strm1_data       ),      
               .std__pe46__lane6_strm1_data_valid    ( std__pe46__lane6_strm1_data_valid ),      
               .std__pe46__lane6_strm1_data_mask     ( std__pe46__lane6_strm1_data_mask  ),      

               // PE 46, Lane 7                 
               .pe46__std__lane7_strm0_ready         ( pe46__std__lane7_strm0_ready      ),      
               .std__pe46__lane7_strm0_cntl          ( std__pe46__lane7_strm0_cntl       ),      
               .std__pe46__lane7_strm0_data          ( std__pe46__lane7_strm0_data       ),      
               .std__pe46__lane7_strm0_data_valid    ( std__pe46__lane7_strm0_data_valid ),      
               .std__pe46__lane7_strm0_data_mask     ( std__pe46__lane7_strm0_data_mask  ),      

               .pe46__std__lane7_strm1_ready         ( pe46__std__lane7_strm1_ready      ),      
               .std__pe46__lane7_strm1_cntl          ( std__pe46__lane7_strm1_cntl       ),      
               .std__pe46__lane7_strm1_data          ( std__pe46__lane7_strm1_data       ),      
               .std__pe46__lane7_strm1_data_valid    ( std__pe46__lane7_strm1_data_valid ),      
               .std__pe46__lane7_strm1_data_mask     ( std__pe46__lane7_strm1_data_mask  ),      

               // PE 46, Lane 8                 
               .pe46__std__lane8_strm0_ready         ( pe46__std__lane8_strm0_ready      ),      
               .std__pe46__lane8_strm0_cntl          ( std__pe46__lane8_strm0_cntl       ),      
               .std__pe46__lane8_strm0_data          ( std__pe46__lane8_strm0_data       ),      
               .std__pe46__lane8_strm0_data_valid    ( std__pe46__lane8_strm0_data_valid ),      
               .std__pe46__lane8_strm0_data_mask     ( std__pe46__lane8_strm0_data_mask  ),      

               .pe46__std__lane8_strm1_ready         ( pe46__std__lane8_strm1_ready      ),      
               .std__pe46__lane8_strm1_cntl          ( std__pe46__lane8_strm1_cntl       ),      
               .std__pe46__lane8_strm1_data          ( std__pe46__lane8_strm1_data       ),      
               .std__pe46__lane8_strm1_data_valid    ( std__pe46__lane8_strm1_data_valid ),      
               .std__pe46__lane8_strm1_data_mask     ( std__pe46__lane8_strm1_data_mask  ),      

               // PE 46, Lane 9                 
               .pe46__std__lane9_strm0_ready         ( pe46__std__lane9_strm0_ready      ),      
               .std__pe46__lane9_strm0_cntl          ( std__pe46__lane9_strm0_cntl       ),      
               .std__pe46__lane9_strm0_data          ( std__pe46__lane9_strm0_data       ),      
               .std__pe46__lane9_strm0_data_valid    ( std__pe46__lane9_strm0_data_valid ),      
               .std__pe46__lane9_strm0_data_mask     ( std__pe46__lane9_strm0_data_mask  ),      

               .pe46__std__lane9_strm1_ready         ( pe46__std__lane9_strm1_ready      ),      
               .std__pe46__lane9_strm1_cntl          ( std__pe46__lane9_strm1_cntl       ),      
               .std__pe46__lane9_strm1_data          ( std__pe46__lane9_strm1_data       ),      
               .std__pe46__lane9_strm1_data_valid    ( std__pe46__lane9_strm1_data_valid ),      
               .std__pe46__lane9_strm1_data_mask     ( std__pe46__lane9_strm1_data_mask  ),      

               // PE 46, Lane 10                 
               .pe46__std__lane10_strm0_ready         ( pe46__std__lane10_strm0_ready      ),      
               .std__pe46__lane10_strm0_cntl          ( std__pe46__lane10_strm0_cntl       ),      
               .std__pe46__lane10_strm0_data          ( std__pe46__lane10_strm0_data       ),      
               .std__pe46__lane10_strm0_data_valid    ( std__pe46__lane10_strm0_data_valid ),      
               .std__pe46__lane10_strm0_data_mask     ( std__pe46__lane10_strm0_data_mask  ),      

               .pe46__std__lane10_strm1_ready         ( pe46__std__lane10_strm1_ready      ),      
               .std__pe46__lane10_strm1_cntl          ( std__pe46__lane10_strm1_cntl       ),      
               .std__pe46__lane10_strm1_data          ( std__pe46__lane10_strm1_data       ),      
               .std__pe46__lane10_strm1_data_valid    ( std__pe46__lane10_strm1_data_valid ),      
               .std__pe46__lane10_strm1_data_mask     ( std__pe46__lane10_strm1_data_mask  ),      

               // PE 46, Lane 11                 
               .pe46__std__lane11_strm0_ready         ( pe46__std__lane11_strm0_ready      ),      
               .std__pe46__lane11_strm0_cntl          ( std__pe46__lane11_strm0_cntl       ),      
               .std__pe46__lane11_strm0_data          ( std__pe46__lane11_strm0_data       ),      
               .std__pe46__lane11_strm0_data_valid    ( std__pe46__lane11_strm0_data_valid ),      
               .std__pe46__lane11_strm0_data_mask     ( std__pe46__lane11_strm0_data_mask  ),      

               .pe46__std__lane11_strm1_ready         ( pe46__std__lane11_strm1_ready      ),      
               .std__pe46__lane11_strm1_cntl          ( std__pe46__lane11_strm1_cntl       ),      
               .std__pe46__lane11_strm1_data          ( std__pe46__lane11_strm1_data       ),      
               .std__pe46__lane11_strm1_data_valid    ( std__pe46__lane11_strm1_data_valid ),      
               .std__pe46__lane11_strm1_data_mask     ( std__pe46__lane11_strm1_data_mask  ),      

               // PE 46, Lane 12                 
               .pe46__std__lane12_strm0_ready         ( pe46__std__lane12_strm0_ready      ),      
               .std__pe46__lane12_strm0_cntl          ( std__pe46__lane12_strm0_cntl       ),      
               .std__pe46__lane12_strm0_data          ( std__pe46__lane12_strm0_data       ),      
               .std__pe46__lane12_strm0_data_valid    ( std__pe46__lane12_strm0_data_valid ),      
               .std__pe46__lane12_strm0_data_mask     ( std__pe46__lane12_strm0_data_mask  ),      

               .pe46__std__lane12_strm1_ready         ( pe46__std__lane12_strm1_ready      ),      
               .std__pe46__lane12_strm1_cntl          ( std__pe46__lane12_strm1_cntl       ),      
               .std__pe46__lane12_strm1_data          ( std__pe46__lane12_strm1_data       ),      
               .std__pe46__lane12_strm1_data_valid    ( std__pe46__lane12_strm1_data_valid ),      
               .std__pe46__lane12_strm1_data_mask     ( std__pe46__lane12_strm1_data_mask  ),      

               // PE 46, Lane 13                 
               .pe46__std__lane13_strm0_ready         ( pe46__std__lane13_strm0_ready      ),      
               .std__pe46__lane13_strm0_cntl          ( std__pe46__lane13_strm0_cntl       ),      
               .std__pe46__lane13_strm0_data          ( std__pe46__lane13_strm0_data       ),      
               .std__pe46__lane13_strm0_data_valid    ( std__pe46__lane13_strm0_data_valid ),      
               .std__pe46__lane13_strm0_data_mask     ( std__pe46__lane13_strm0_data_mask  ),      

               .pe46__std__lane13_strm1_ready         ( pe46__std__lane13_strm1_ready      ),      
               .std__pe46__lane13_strm1_cntl          ( std__pe46__lane13_strm1_cntl       ),      
               .std__pe46__lane13_strm1_data          ( std__pe46__lane13_strm1_data       ),      
               .std__pe46__lane13_strm1_data_valid    ( std__pe46__lane13_strm1_data_valid ),      
               .std__pe46__lane13_strm1_data_mask     ( std__pe46__lane13_strm1_data_mask  ),      

               // PE 46, Lane 14                 
               .pe46__std__lane14_strm0_ready         ( pe46__std__lane14_strm0_ready      ),      
               .std__pe46__lane14_strm0_cntl          ( std__pe46__lane14_strm0_cntl       ),      
               .std__pe46__lane14_strm0_data          ( std__pe46__lane14_strm0_data       ),      
               .std__pe46__lane14_strm0_data_valid    ( std__pe46__lane14_strm0_data_valid ),      
               .std__pe46__lane14_strm0_data_mask     ( std__pe46__lane14_strm0_data_mask  ),      

               .pe46__std__lane14_strm1_ready         ( pe46__std__lane14_strm1_ready      ),      
               .std__pe46__lane14_strm1_cntl          ( std__pe46__lane14_strm1_cntl       ),      
               .std__pe46__lane14_strm1_data          ( std__pe46__lane14_strm1_data       ),      
               .std__pe46__lane14_strm1_data_valid    ( std__pe46__lane14_strm1_data_valid ),      
               .std__pe46__lane14_strm1_data_mask     ( std__pe46__lane14_strm1_data_mask  ),      

               // PE 46, Lane 15                 
               .pe46__std__lane15_strm0_ready         ( pe46__std__lane15_strm0_ready      ),      
               .std__pe46__lane15_strm0_cntl          ( std__pe46__lane15_strm0_cntl       ),      
               .std__pe46__lane15_strm0_data          ( std__pe46__lane15_strm0_data       ),      
               .std__pe46__lane15_strm0_data_valid    ( std__pe46__lane15_strm0_data_valid ),      
               .std__pe46__lane15_strm0_data_mask     ( std__pe46__lane15_strm0_data_mask  ),      

               .pe46__std__lane15_strm1_ready         ( pe46__std__lane15_strm1_ready      ),      
               .std__pe46__lane15_strm1_cntl          ( std__pe46__lane15_strm1_cntl       ),      
               .std__pe46__lane15_strm1_data          ( std__pe46__lane15_strm1_data       ),      
               .std__pe46__lane15_strm1_data_valid    ( std__pe46__lane15_strm1_data_valid ),      
               .std__pe46__lane15_strm1_data_mask     ( std__pe46__lane15_strm1_data_mask  ),      

               // PE 46, Lane 16                 
               .pe46__std__lane16_strm0_ready         ( pe46__std__lane16_strm0_ready      ),      
               .std__pe46__lane16_strm0_cntl          ( std__pe46__lane16_strm0_cntl       ),      
               .std__pe46__lane16_strm0_data          ( std__pe46__lane16_strm0_data       ),      
               .std__pe46__lane16_strm0_data_valid    ( std__pe46__lane16_strm0_data_valid ),      
               .std__pe46__lane16_strm0_data_mask     ( std__pe46__lane16_strm0_data_mask  ),      

               .pe46__std__lane16_strm1_ready         ( pe46__std__lane16_strm1_ready      ),      
               .std__pe46__lane16_strm1_cntl          ( std__pe46__lane16_strm1_cntl       ),      
               .std__pe46__lane16_strm1_data          ( std__pe46__lane16_strm1_data       ),      
               .std__pe46__lane16_strm1_data_valid    ( std__pe46__lane16_strm1_data_valid ),      
               .std__pe46__lane16_strm1_data_mask     ( std__pe46__lane16_strm1_data_mask  ),      

               // PE 46, Lane 17                 
               .pe46__std__lane17_strm0_ready         ( pe46__std__lane17_strm0_ready      ),      
               .std__pe46__lane17_strm0_cntl          ( std__pe46__lane17_strm0_cntl       ),      
               .std__pe46__lane17_strm0_data          ( std__pe46__lane17_strm0_data       ),      
               .std__pe46__lane17_strm0_data_valid    ( std__pe46__lane17_strm0_data_valid ),      
               .std__pe46__lane17_strm0_data_mask     ( std__pe46__lane17_strm0_data_mask  ),      

               .pe46__std__lane17_strm1_ready         ( pe46__std__lane17_strm1_ready      ),      
               .std__pe46__lane17_strm1_cntl          ( std__pe46__lane17_strm1_cntl       ),      
               .std__pe46__lane17_strm1_data          ( std__pe46__lane17_strm1_data       ),      
               .std__pe46__lane17_strm1_data_valid    ( std__pe46__lane17_strm1_data_valid ),      
               .std__pe46__lane17_strm1_data_mask     ( std__pe46__lane17_strm1_data_mask  ),      

               // PE 46, Lane 18                 
               .pe46__std__lane18_strm0_ready         ( pe46__std__lane18_strm0_ready      ),      
               .std__pe46__lane18_strm0_cntl          ( std__pe46__lane18_strm0_cntl       ),      
               .std__pe46__lane18_strm0_data          ( std__pe46__lane18_strm0_data       ),      
               .std__pe46__lane18_strm0_data_valid    ( std__pe46__lane18_strm0_data_valid ),      
               .std__pe46__lane18_strm0_data_mask     ( std__pe46__lane18_strm0_data_mask  ),      

               .pe46__std__lane18_strm1_ready         ( pe46__std__lane18_strm1_ready      ),      
               .std__pe46__lane18_strm1_cntl          ( std__pe46__lane18_strm1_cntl       ),      
               .std__pe46__lane18_strm1_data          ( std__pe46__lane18_strm1_data       ),      
               .std__pe46__lane18_strm1_data_valid    ( std__pe46__lane18_strm1_data_valid ),      
               .std__pe46__lane18_strm1_data_mask     ( std__pe46__lane18_strm1_data_mask  ),      

               // PE 46, Lane 19                 
               .pe46__std__lane19_strm0_ready         ( pe46__std__lane19_strm0_ready      ),      
               .std__pe46__lane19_strm0_cntl          ( std__pe46__lane19_strm0_cntl       ),      
               .std__pe46__lane19_strm0_data          ( std__pe46__lane19_strm0_data       ),      
               .std__pe46__lane19_strm0_data_valid    ( std__pe46__lane19_strm0_data_valid ),      
               .std__pe46__lane19_strm0_data_mask     ( std__pe46__lane19_strm0_data_mask  ),      

               .pe46__std__lane19_strm1_ready         ( pe46__std__lane19_strm1_ready      ),      
               .std__pe46__lane19_strm1_cntl          ( std__pe46__lane19_strm1_cntl       ),      
               .std__pe46__lane19_strm1_data          ( std__pe46__lane19_strm1_data       ),      
               .std__pe46__lane19_strm1_data_valid    ( std__pe46__lane19_strm1_data_valid ),      
               .std__pe46__lane19_strm1_data_mask     ( std__pe46__lane19_strm1_data_mask  ),      

               // PE 46, Lane 20                 
               .pe46__std__lane20_strm0_ready         ( pe46__std__lane20_strm0_ready      ),      
               .std__pe46__lane20_strm0_cntl          ( std__pe46__lane20_strm0_cntl       ),      
               .std__pe46__lane20_strm0_data          ( std__pe46__lane20_strm0_data       ),      
               .std__pe46__lane20_strm0_data_valid    ( std__pe46__lane20_strm0_data_valid ),      
               .std__pe46__lane20_strm0_data_mask     ( std__pe46__lane20_strm0_data_mask  ),      

               .pe46__std__lane20_strm1_ready         ( pe46__std__lane20_strm1_ready      ),      
               .std__pe46__lane20_strm1_cntl          ( std__pe46__lane20_strm1_cntl       ),      
               .std__pe46__lane20_strm1_data          ( std__pe46__lane20_strm1_data       ),      
               .std__pe46__lane20_strm1_data_valid    ( std__pe46__lane20_strm1_data_valid ),      
               .std__pe46__lane20_strm1_data_mask     ( std__pe46__lane20_strm1_data_mask  ),      

               // PE 46, Lane 21                 
               .pe46__std__lane21_strm0_ready         ( pe46__std__lane21_strm0_ready      ),      
               .std__pe46__lane21_strm0_cntl          ( std__pe46__lane21_strm0_cntl       ),      
               .std__pe46__lane21_strm0_data          ( std__pe46__lane21_strm0_data       ),      
               .std__pe46__lane21_strm0_data_valid    ( std__pe46__lane21_strm0_data_valid ),      
               .std__pe46__lane21_strm0_data_mask     ( std__pe46__lane21_strm0_data_mask  ),      

               .pe46__std__lane21_strm1_ready         ( pe46__std__lane21_strm1_ready      ),      
               .std__pe46__lane21_strm1_cntl          ( std__pe46__lane21_strm1_cntl       ),      
               .std__pe46__lane21_strm1_data          ( std__pe46__lane21_strm1_data       ),      
               .std__pe46__lane21_strm1_data_valid    ( std__pe46__lane21_strm1_data_valid ),      
               .std__pe46__lane21_strm1_data_mask     ( std__pe46__lane21_strm1_data_mask  ),      

               // PE 46, Lane 22                 
               .pe46__std__lane22_strm0_ready         ( pe46__std__lane22_strm0_ready      ),      
               .std__pe46__lane22_strm0_cntl          ( std__pe46__lane22_strm0_cntl       ),      
               .std__pe46__lane22_strm0_data          ( std__pe46__lane22_strm0_data       ),      
               .std__pe46__lane22_strm0_data_valid    ( std__pe46__lane22_strm0_data_valid ),      
               .std__pe46__lane22_strm0_data_mask     ( std__pe46__lane22_strm0_data_mask  ),      

               .pe46__std__lane22_strm1_ready         ( pe46__std__lane22_strm1_ready      ),      
               .std__pe46__lane22_strm1_cntl          ( std__pe46__lane22_strm1_cntl       ),      
               .std__pe46__lane22_strm1_data          ( std__pe46__lane22_strm1_data       ),      
               .std__pe46__lane22_strm1_data_valid    ( std__pe46__lane22_strm1_data_valid ),      
               .std__pe46__lane22_strm1_data_mask     ( std__pe46__lane22_strm1_data_mask  ),      

               // PE 46, Lane 23                 
               .pe46__std__lane23_strm0_ready         ( pe46__std__lane23_strm0_ready      ),      
               .std__pe46__lane23_strm0_cntl          ( std__pe46__lane23_strm0_cntl       ),      
               .std__pe46__lane23_strm0_data          ( std__pe46__lane23_strm0_data       ),      
               .std__pe46__lane23_strm0_data_valid    ( std__pe46__lane23_strm0_data_valid ),      
               .std__pe46__lane23_strm0_data_mask     ( std__pe46__lane23_strm0_data_mask  ),      

               .pe46__std__lane23_strm1_ready         ( pe46__std__lane23_strm1_ready      ),      
               .std__pe46__lane23_strm1_cntl          ( std__pe46__lane23_strm1_cntl       ),      
               .std__pe46__lane23_strm1_data          ( std__pe46__lane23_strm1_data       ),      
               .std__pe46__lane23_strm1_data_valid    ( std__pe46__lane23_strm1_data_valid ),      
               .std__pe46__lane23_strm1_data_mask     ( std__pe46__lane23_strm1_data_mask  ),      

               // PE 46, Lane 24                 
               .pe46__std__lane24_strm0_ready         ( pe46__std__lane24_strm0_ready      ),      
               .std__pe46__lane24_strm0_cntl          ( std__pe46__lane24_strm0_cntl       ),      
               .std__pe46__lane24_strm0_data          ( std__pe46__lane24_strm0_data       ),      
               .std__pe46__lane24_strm0_data_valid    ( std__pe46__lane24_strm0_data_valid ),      
               .std__pe46__lane24_strm0_data_mask     ( std__pe46__lane24_strm0_data_mask  ),      

               .pe46__std__lane24_strm1_ready         ( pe46__std__lane24_strm1_ready      ),      
               .std__pe46__lane24_strm1_cntl          ( std__pe46__lane24_strm1_cntl       ),      
               .std__pe46__lane24_strm1_data          ( std__pe46__lane24_strm1_data       ),      
               .std__pe46__lane24_strm1_data_valid    ( std__pe46__lane24_strm1_data_valid ),      
               .std__pe46__lane24_strm1_data_mask     ( std__pe46__lane24_strm1_data_mask  ),      

               // PE 46, Lane 25                 
               .pe46__std__lane25_strm0_ready         ( pe46__std__lane25_strm0_ready      ),      
               .std__pe46__lane25_strm0_cntl          ( std__pe46__lane25_strm0_cntl       ),      
               .std__pe46__lane25_strm0_data          ( std__pe46__lane25_strm0_data       ),      
               .std__pe46__lane25_strm0_data_valid    ( std__pe46__lane25_strm0_data_valid ),      
               .std__pe46__lane25_strm0_data_mask     ( std__pe46__lane25_strm0_data_mask  ),      

               .pe46__std__lane25_strm1_ready         ( pe46__std__lane25_strm1_ready      ),      
               .std__pe46__lane25_strm1_cntl          ( std__pe46__lane25_strm1_cntl       ),      
               .std__pe46__lane25_strm1_data          ( std__pe46__lane25_strm1_data       ),      
               .std__pe46__lane25_strm1_data_valid    ( std__pe46__lane25_strm1_data_valid ),      
               .std__pe46__lane25_strm1_data_mask     ( std__pe46__lane25_strm1_data_mask  ),      

               // PE 46, Lane 26                 
               .pe46__std__lane26_strm0_ready         ( pe46__std__lane26_strm0_ready      ),      
               .std__pe46__lane26_strm0_cntl          ( std__pe46__lane26_strm0_cntl       ),      
               .std__pe46__lane26_strm0_data          ( std__pe46__lane26_strm0_data       ),      
               .std__pe46__lane26_strm0_data_valid    ( std__pe46__lane26_strm0_data_valid ),      
               .std__pe46__lane26_strm0_data_mask     ( std__pe46__lane26_strm0_data_mask  ),      

               .pe46__std__lane26_strm1_ready         ( pe46__std__lane26_strm1_ready      ),      
               .std__pe46__lane26_strm1_cntl          ( std__pe46__lane26_strm1_cntl       ),      
               .std__pe46__lane26_strm1_data          ( std__pe46__lane26_strm1_data       ),      
               .std__pe46__lane26_strm1_data_valid    ( std__pe46__lane26_strm1_data_valid ),      
               .std__pe46__lane26_strm1_data_mask     ( std__pe46__lane26_strm1_data_mask  ),      

               // PE 46, Lane 27                 
               .pe46__std__lane27_strm0_ready         ( pe46__std__lane27_strm0_ready      ),      
               .std__pe46__lane27_strm0_cntl          ( std__pe46__lane27_strm0_cntl       ),      
               .std__pe46__lane27_strm0_data          ( std__pe46__lane27_strm0_data       ),      
               .std__pe46__lane27_strm0_data_valid    ( std__pe46__lane27_strm0_data_valid ),      
               .std__pe46__lane27_strm0_data_mask     ( std__pe46__lane27_strm0_data_mask  ),      

               .pe46__std__lane27_strm1_ready         ( pe46__std__lane27_strm1_ready      ),      
               .std__pe46__lane27_strm1_cntl          ( std__pe46__lane27_strm1_cntl       ),      
               .std__pe46__lane27_strm1_data          ( std__pe46__lane27_strm1_data       ),      
               .std__pe46__lane27_strm1_data_valid    ( std__pe46__lane27_strm1_data_valid ),      
               .std__pe46__lane27_strm1_data_mask     ( std__pe46__lane27_strm1_data_mask  ),      

               // PE 46, Lane 28                 
               .pe46__std__lane28_strm0_ready         ( pe46__std__lane28_strm0_ready      ),      
               .std__pe46__lane28_strm0_cntl          ( std__pe46__lane28_strm0_cntl       ),      
               .std__pe46__lane28_strm0_data          ( std__pe46__lane28_strm0_data       ),      
               .std__pe46__lane28_strm0_data_valid    ( std__pe46__lane28_strm0_data_valid ),      
               .std__pe46__lane28_strm0_data_mask     ( std__pe46__lane28_strm0_data_mask  ),      

               .pe46__std__lane28_strm1_ready         ( pe46__std__lane28_strm1_ready      ),      
               .std__pe46__lane28_strm1_cntl          ( std__pe46__lane28_strm1_cntl       ),      
               .std__pe46__lane28_strm1_data          ( std__pe46__lane28_strm1_data       ),      
               .std__pe46__lane28_strm1_data_valid    ( std__pe46__lane28_strm1_data_valid ),      
               .std__pe46__lane28_strm1_data_mask     ( std__pe46__lane28_strm1_data_mask  ),      

               // PE 46, Lane 29                 
               .pe46__std__lane29_strm0_ready         ( pe46__std__lane29_strm0_ready      ),      
               .std__pe46__lane29_strm0_cntl          ( std__pe46__lane29_strm0_cntl       ),      
               .std__pe46__lane29_strm0_data          ( std__pe46__lane29_strm0_data       ),      
               .std__pe46__lane29_strm0_data_valid    ( std__pe46__lane29_strm0_data_valid ),      
               .std__pe46__lane29_strm0_data_mask     ( std__pe46__lane29_strm0_data_mask  ),      

               .pe46__std__lane29_strm1_ready         ( pe46__std__lane29_strm1_ready      ),      
               .std__pe46__lane29_strm1_cntl          ( std__pe46__lane29_strm1_cntl       ),      
               .std__pe46__lane29_strm1_data          ( std__pe46__lane29_strm1_data       ),      
               .std__pe46__lane29_strm1_data_valid    ( std__pe46__lane29_strm1_data_valid ),      
               .std__pe46__lane29_strm1_data_mask     ( std__pe46__lane29_strm1_data_mask  ),      

               // PE 46, Lane 30                 
               .pe46__std__lane30_strm0_ready         ( pe46__std__lane30_strm0_ready      ),      
               .std__pe46__lane30_strm0_cntl          ( std__pe46__lane30_strm0_cntl       ),      
               .std__pe46__lane30_strm0_data          ( std__pe46__lane30_strm0_data       ),      
               .std__pe46__lane30_strm0_data_valid    ( std__pe46__lane30_strm0_data_valid ),      
               .std__pe46__lane30_strm0_data_mask     ( std__pe46__lane30_strm0_data_mask  ),      

               .pe46__std__lane30_strm1_ready         ( pe46__std__lane30_strm1_ready      ),      
               .std__pe46__lane30_strm1_cntl          ( std__pe46__lane30_strm1_cntl       ),      
               .std__pe46__lane30_strm1_data          ( std__pe46__lane30_strm1_data       ),      
               .std__pe46__lane30_strm1_data_valid    ( std__pe46__lane30_strm1_data_valid ),      
               .std__pe46__lane30_strm1_data_mask     ( std__pe46__lane30_strm1_data_mask  ),      

               // PE 46, Lane 31                 
               .pe46__std__lane31_strm0_ready         ( pe46__std__lane31_strm0_ready      ),      
               .std__pe46__lane31_strm0_cntl          ( std__pe46__lane31_strm0_cntl       ),      
               .std__pe46__lane31_strm0_data          ( std__pe46__lane31_strm0_data       ),      
               .std__pe46__lane31_strm0_data_valid    ( std__pe46__lane31_strm0_data_valid ),      
               .std__pe46__lane31_strm0_data_mask     ( std__pe46__lane31_strm0_data_mask  ),      

               .pe46__std__lane31_strm1_ready         ( pe46__std__lane31_strm1_ready      ),      
               .std__pe46__lane31_strm1_cntl          ( std__pe46__lane31_strm1_cntl       ),      
               .std__pe46__lane31_strm1_data          ( std__pe46__lane31_strm1_data       ),      
               .std__pe46__lane31_strm1_data_valid    ( std__pe46__lane31_strm1_data_valid ),      
               .std__pe46__lane31_strm1_data_mask     ( std__pe46__lane31_strm1_data_mask  ),      

               // PE 47, Lane 0                 
               .pe47__std__lane0_strm0_ready         ( pe47__std__lane0_strm0_ready      ),      
               .std__pe47__lane0_strm0_cntl          ( std__pe47__lane0_strm0_cntl       ),      
               .std__pe47__lane0_strm0_data          ( std__pe47__lane0_strm0_data       ),      
               .std__pe47__lane0_strm0_data_valid    ( std__pe47__lane0_strm0_data_valid ),      
               .std__pe47__lane0_strm0_data_mask     ( std__pe47__lane0_strm0_data_mask  ),      

               .pe47__std__lane0_strm1_ready         ( pe47__std__lane0_strm1_ready      ),      
               .std__pe47__lane0_strm1_cntl          ( std__pe47__lane0_strm1_cntl       ),      
               .std__pe47__lane0_strm1_data          ( std__pe47__lane0_strm1_data       ),      
               .std__pe47__lane0_strm1_data_valid    ( std__pe47__lane0_strm1_data_valid ),      
               .std__pe47__lane0_strm1_data_mask     ( std__pe47__lane0_strm1_data_mask  ),      

               // PE 47, Lane 1                 
               .pe47__std__lane1_strm0_ready         ( pe47__std__lane1_strm0_ready      ),      
               .std__pe47__lane1_strm0_cntl          ( std__pe47__lane1_strm0_cntl       ),      
               .std__pe47__lane1_strm0_data          ( std__pe47__lane1_strm0_data       ),      
               .std__pe47__lane1_strm0_data_valid    ( std__pe47__lane1_strm0_data_valid ),      
               .std__pe47__lane1_strm0_data_mask     ( std__pe47__lane1_strm0_data_mask  ),      

               .pe47__std__lane1_strm1_ready         ( pe47__std__lane1_strm1_ready      ),      
               .std__pe47__lane1_strm1_cntl          ( std__pe47__lane1_strm1_cntl       ),      
               .std__pe47__lane1_strm1_data          ( std__pe47__lane1_strm1_data       ),      
               .std__pe47__lane1_strm1_data_valid    ( std__pe47__lane1_strm1_data_valid ),      
               .std__pe47__lane1_strm1_data_mask     ( std__pe47__lane1_strm1_data_mask  ),      

               // PE 47, Lane 2                 
               .pe47__std__lane2_strm0_ready         ( pe47__std__lane2_strm0_ready      ),      
               .std__pe47__lane2_strm0_cntl          ( std__pe47__lane2_strm0_cntl       ),      
               .std__pe47__lane2_strm0_data          ( std__pe47__lane2_strm0_data       ),      
               .std__pe47__lane2_strm0_data_valid    ( std__pe47__lane2_strm0_data_valid ),      
               .std__pe47__lane2_strm0_data_mask     ( std__pe47__lane2_strm0_data_mask  ),      

               .pe47__std__lane2_strm1_ready         ( pe47__std__lane2_strm1_ready      ),      
               .std__pe47__lane2_strm1_cntl          ( std__pe47__lane2_strm1_cntl       ),      
               .std__pe47__lane2_strm1_data          ( std__pe47__lane2_strm1_data       ),      
               .std__pe47__lane2_strm1_data_valid    ( std__pe47__lane2_strm1_data_valid ),      
               .std__pe47__lane2_strm1_data_mask     ( std__pe47__lane2_strm1_data_mask  ),      

               // PE 47, Lane 3                 
               .pe47__std__lane3_strm0_ready         ( pe47__std__lane3_strm0_ready      ),      
               .std__pe47__lane3_strm0_cntl          ( std__pe47__lane3_strm0_cntl       ),      
               .std__pe47__lane3_strm0_data          ( std__pe47__lane3_strm0_data       ),      
               .std__pe47__lane3_strm0_data_valid    ( std__pe47__lane3_strm0_data_valid ),      
               .std__pe47__lane3_strm0_data_mask     ( std__pe47__lane3_strm0_data_mask  ),      

               .pe47__std__lane3_strm1_ready         ( pe47__std__lane3_strm1_ready      ),      
               .std__pe47__lane3_strm1_cntl          ( std__pe47__lane3_strm1_cntl       ),      
               .std__pe47__lane3_strm1_data          ( std__pe47__lane3_strm1_data       ),      
               .std__pe47__lane3_strm1_data_valid    ( std__pe47__lane3_strm1_data_valid ),      
               .std__pe47__lane3_strm1_data_mask     ( std__pe47__lane3_strm1_data_mask  ),      

               // PE 47, Lane 4                 
               .pe47__std__lane4_strm0_ready         ( pe47__std__lane4_strm0_ready      ),      
               .std__pe47__lane4_strm0_cntl          ( std__pe47__lane4_strm0_cntl       ),      
               .std__pe47__lane4_strm0_data          ( std__pe47__lane4_strm0_data       ),      
               .std__pe47__lane4_strm0_data_valid    ( std__pe47__lane4_strm0_data_valid ),      
               .std__pe47__lane4_strm0_data_mask     ( std__pe47__lane4_strm0_data_mask  ),      

               .pe47__std__lane4_strm1_ready         ( pe47__std__lane4_strm1_ready      ),      
               .std__pe47__lane4_strm1_cntl          ( std__pe47__lane4_strm1_cntl       ),      
               .std__pe47__lane4_strm1_data          ( std__pe47__lane4_strm1_data       ),      
               .std__pe47__lane4_strm1_data_valid    ( std__pe47__lane4_strm1_data_valid ),      
               .std__pe47__lane4_strm1_data_mask     ( std__pe47__lane4_strm1_data_mask  ),      

               // PE 47, Lane 5                 
               .pe47__std__lane5_strm0_ready         ( pe47__std__lane5_strm0_ready      ),      
               .std__pe47__lane5_strm0_cntl          ( std__pe47__lane5_strm0_cntl       ),      
               .std__pe47__lane5_strm0_data          ( std__pe47__lane5_strm0_data       ),      
               .std__pe47__lane5_strm0_data_valid    ( std__pe47__lane5_strm0_data_valid ),      
               .std__pe47__lane5_strm0_data_mask     ( std__pe47__lane5_strm0_data_mask  ),      

               .pe47__std__lane5_strm1_ready         ( pe47__std__lane5_strm1_ready      ),      
               .std__pe47__lane5_strm1_cntl          ( std__pe47__lane5_strm1_cntl       ),      
               .std__pe47__lane5_strm1_data          ( std__pe47__lane5_strm1_data       ),      
               .std__pe47__lane5_strm1_data_valid    ( std__pe47__lane5_strm1_data_valid ),      
               .std__pe47__lane5_strm1_data_mask     ( std__pe47__lane5_strm1_data_mask  ),      

               // PE 47, Lane 6                 
               .pe47__std__lane6_strm0_ready         ( pe47__std__lane6_strm0_ready      ),      
               .std__pe47__lane6_strm0_cntl          ( std__pe47__lane6_strm0_cntl       ),      
               .std__pe47__lane6_strm0_data          ( std__pe47__lane6_strm0_data       ),      
               .std__pe47__lane6_strm0_data_valid    ( std__pe47__lane6_strm0_data_valid ),      
               .std__pe47__lane6_strm0_data_mask     ( std__pe47__lane6_strm0_data_mask  ),      

               .pe47__std__lane6_strm1_ready         ( pe47__std__lane6_strm1_ready      ),      
               .std__pe47__lane6_strm1_cntl          ( std__pe47__lane6_strm1_cntl       ),      
               .std__pe47__lane6_strm1_data          ( std__pe47__lane6_strm1_data       ),      
               .std__pe47__lane6_strm1_data_valid    ( std__pe47__lane6_strm1_data_valid ),      
               .std__pe47__lane6_strm1_data_mask     ( std__pe47__lane6_strm1_data_mask  ),      

               // PE 47, Lane 7                 
               .pe47__std__lane7_strm0_ready         ( pe47__std__lane7_strm0_ready      ),      
               .std__pe47__lane7_strm0_cntl          ( std__pe47__lane7_strm0_cntl       ),      
               .std__pe47__lane7_strm0_data          ( std__pe47__lane7_strm0_data       ),      
               .std__pe47__lane7_strm0_data_valid    ( std__pe47__lane7_strm0_data_valid ),      
               .std__pe47__lane7_strm0_data_mask     ( std__pe47__lane7_strm0_data_mask  ),      

               .pe47__std__lane7_strm1_ready         ( pe47__std__lane7_strm1_ready      ),      
               .std__pe47__lane7_strm1_cntl          ( std__pe47__lane7_strm1_cntl       ),      
               .std__pe47__lane7_strm1_data          ( std__pe47__lane7_strm1_data       ),      
               .std__pe47__lane7_strm1_data_valid    ( std__pe47__lane7_strm1_data_valid ),      
               .std__pe47__lane7_strm1_data_mask     ( std__pe47__lane7_strm1_data_mask  ),      

               // PE 47, Lane 8                 
               .pe47__std__lane8_strm0_ready         ( pe47__std__lane8_strm0_ready      ),      
               .std__pe47__lane8_strm0_cntl          ( std__pe47__lane8_strm0_cntl       ),      
               .std__pe47__lane8_strm0_data          ( std__pe47__lane8_strm0_data       ),      
               .std__pe47__lane8_strm0_data_valid    ( std__pe47__lane8_strm0_data_valid ),      
               .std__pe47__lane8_strm0_data_mask     ( std__pe47__lane8_strm0_data_mask  ),      

               .pe47__std__lane8_strm1_ready         ( pe47__std__lane8_strm1_ready      ),      
               .std__pe47__lane8_strm1_cntl          ( std__pe47__lane8_strm1_cntl       ),      
               .std__pe47__lane8_strm1_data          ( std__pe47__lane8_strm1_data       ),      
               .std__pe47__lane8_strm1_data_valid    ( std__pe47__lane8_strm1_data_valid ),      
               .std__pe47__lane8_strm1_data_mask     ( std__pe47__lane8_strm1_data_mask  ),      

               // PE 47, Lane 9                 
               .pe47__std__lane9_strm0_ready         ( pe47__std__lane9_strm0_ready      ),      
               .std__pe47__lane9_strm0_cntl          ( std__pe47__lane9_strm0_cntl       ),      
               .std__pe47__lane9_strm0_data          ( std__pe47__lane9_strm0_data       ),      
               .std__pe47__lane9_strm0_data_valid    ( std__pe47__lane9_strm0_data_valid ),      
               .std__pe47__lane9_strm0_data_mask     ( std__pe47__lane9_strm0_data_mask  ),      

               .pe47__std__lane9_strm1_ready         ( pe47__std__lane9_strm1_ready      ),      
               .std__pe47__lane9_strm1_cntl          ( std__pe47__lane9_strm1_cntl       ),      
               .std__pe47__lane9_strm1_data          ( std__pe47__lane9_strm1_data       ),      
               .std__pe47__lane9_strm1_data_valid    ( std__pe47__lane9_strm1_data_valid ),      
               .std__pe47__lane9_strm1_data_mask     ( std__pe47__lane9_strm1_data_mask  ),      

               // PE 47, Lane 10                 
               .pe47__std__lane10_strm0_ready         ( pe47__std__lane10_strm0_ready      ),      
               .std__pe47__lane10_strm0_cntl          ( std__pe47__lane10_strm0_cntl       ),      
               .std__pe47__lane10_strm0_data          ( std__pe47__lane10_strm0_data       ),      
               .std__pe47__lane10_strm0_data_valid    ( std__pe47__lane10_strm0_data_valid ),      
               .std__pe47__lane10_strm0_data_mask     ( std__pe47__lane10_strm0_data_mask  ),      

               .pe47__std__lane10_strm1_ready         ( pe47__std__lane10_strm1_ready      ),      
               .std__pe47__lane10_strm1_cntl          ( std__pe47__lane10_strm1_cntl       ),      
               .std__pe47__lane10_strm1_data          ( std__pe47__lane10_strm1_data       ),      
               .std__pe47__lane10_strm1_data_valid    ( std__pe47__lane10_strm1_data_valid ),      
               .std__pe47__lane10_strm1_data_mask     ( std__pe47__lane10_strm1_data_mask  ),      

               // PE 47, Lane 11                 
               .pe47__std__lane11_strm0_ready         ( pe47__std__lane11_strm0_ready      ),      
               .std__pe47__lane11_strm0_cntl          ( std__pe47__lane11_strm0_cntl       ),      
               .std__pe47__lane11_strm0_data          ( std__pe47__lane11_strm0_data       ),      
               .std__pe47__lane11_strm0_data_valid    ( std__pe47__lane11_strm0_data_valid ),      
               .std__pe47__lane11_strm0_data_mask     ( std__pe47__lane11_strm0_data_mask  ),      

               .pe47__std__lane11_strm1_ready         ( pe47__std__lane11_strm1_ready      ),      
               .std__pe47__lane11_strm1_cntl          ( std__pe47__lane11_strm1_cntl       ),      
               .std__pe47__lane11_strm1_data          ( std__pe47__lane11_strm1_data       ),      
               .std__pe47__lane11_strm1_data_valid    ( std__pe47__lane11_strm1_data_valid ),      
               .std__pe47__lane11_strm1_data_mask     ( std__pe47__lane11_strm1_data_mask  ),      

               // PE 47, Lane 12                 
               .pe47__std__lane12_strm0_ready         ( pe47__std__lane12_strm0_ready      ),      
               .std__pe47__lane12_strm0_cntl          ( std__pe47__lane12_strm0_cntl       ),      
               .std__pe47__lane12_strm0_data          ( std__pe47__lane12_strm0_data       ),      
               .std__pe47__lane12_strm0_data_valid    ( std__pe47__lane12_strm0_data_valid ),      
               .std__pe47__lane12_strm0_data_mask     ( std__pe47__lane12_strm0_data_mask  ),      

               .pe47__std__lane12_strm1_ready         ( pe47__std__lane12_strm1_ready      ),      
               .std__pe47__lane12_strm1_cntl          ( std__pe47__lane12_strm1_cntl       ),      
               .std__pe47__lane12_strm1_data          ( std__pe47__lane12_strm1_data       ),      
               .std__pe47__lane12_strm1_data_valid    ( std__pe47__lane12_strm1_data_valid ),      
               .std__pe47__lane12_strm1_data_mask     ( std__pe47__lane12_strm1_data_mask  ),      

               // PE 47, Lane 13                 
               .pe47__std__lane13_strm0_ready         ( pe47__std__lane13_strm0_ready      ),      
               .std__pe47__lane13_strm0_cntl          ( std__pe47__lane13_strm0_cntl       ),      
               .std__pe47__lane13_strm0_data          ( std__pe47__lane13_strm0_data       ),      
               .std__pe47__lane13_strm0_data_valid    ( std__pe47__lane13_strm0_data_valid ),      
               .std__pe47__lane13_strm0_data_mask     ( std__pe47__lane13_strm0_data_mask  ),      

               .pe47__std__lane13_strm1_ready         ( pe47__std__lane13_strm1_ready      ),      
               .std__pe47__lane13_strm1_cntl          ( std__pe47__lane13_strm1_cntl       ),      
               .std__pe47__lane13_strm1_data          ( std__pe47__lane13_strm1_data       ),      
               .std__pe47__lane13_strm1_data_valid    ( std__pe47__lane13_strm1_data_valid ),      
               .std__pe47__lane13_strm1_data_mask     ( std__pe47__lane13_strm1_data_mask  ),      

               // PE 47, Lane 14                 
               .pe47__std__lane14_strm0_ready         ( pe47__std__lane14_strm0_ready      ),      
               .std__pe47__lane14_strm0_cntl          ( std__pe47__lane14_strm0_cntl       ),      
               .std__pe47__lane14_strm0_data          ( std__pe47__lane14_strm0_data       ),      
               .std__pe47__lane14_strm0_data_valid    ( std__pe47__lane14_strm0_data_valid ),      
               .std__pe47__lane14_strm0_data_mask     ( std__pe47__lane14_strm0_data_mask  ),      

               .pe47__std__lane14_strm1_ready         ( pe47__std__lane14_strm1_ready      ),      
               .std__pe47__lane14_strm1_cntl          ( std__pe47__lane14_strm1_cntl       ),      
               .std__pe47__lane14_strm1_data          ( std__pe47__lane14_strm1_data       ),      
               .std__pe47__lane14_strm1_data_valid    ( std__pe47__lane14_strm1_data_valid ),      
               .std__pe47__lane14_strm1_data_mask     ( std__pe47__lane14_strm1_data_mask  ),      

               // PE 47, Lane 15                 
               .pe47__std__lane15_strm0_ready         ( pe47__std__lane15_strm0_ready      ),      
               .std__pe47__lane15_strm0_cntl          ( std__pe47__lane15_strm0_cntl       ),      
               .std__pe47__lane15_strm0_data          ( std__pe47__lane15_strm0_data       ),      
               .std__pe47__lane15_strm0_data_valid    ( std__pe47__lane15_strm0_data_valid ),      
               .std__pe47__lane15_strm0_data_mask     ( std__pe47__lane15_strm0_data_mask  ),      

               .pe47__std__lane15_strm1_ready         ( pe47__std__lane15_strm1_ready      ),      
               .std__pe47__lane15_strm1_cntl          ( std__pe47__lane15_strm1_cntl       ),      
               .std__pe47__lane15_strm1_data          ( std__pe47__lane15_strm1_data       ),      
               .std__pe47__lane15_strm1_data_valid    ( std__pe47__lane15_strm1_data_valid ),      
               .std__pe47__lane15_strm1_data_mask     ( std__pe47__lane15_strm1_data_mask  ),      

               // PE 47, Lane 16                 
               .pe47__std__lane16_strm0_ready         ( pe47__std__lane16_strm0_ready      ),      
               .std__pe47__lane16_strm0_cntl          ( std__pe47__lane16_strm0_cntl       ),      
               .std__pe47__lane16_strm0_data          ( std__pe47__lane16_strm0_data       ),      
               .std__pe47__lane16_strm0_data_valid    ( std__pe47__lane16_strm0_data_valid ),      
               .std__pe47__lane16_strm0_data_mask     ( std__pe47__lane16_strm0_data_mask  ),      

               .pe47__std__lane16_strm1_ready         ( pe47__std__lane16_strm1_ready      ),      
               .std__pe47__lane16_strm1_cntl          ( std__pe47__lane16_strm1_cntl       ),      
               .std__pe47__lane16_strm1_data          ( std__pe47__lane16_strm1_data       ),      
               .std__pe47__lane16_strm1_data_valid    ( std__pe47__lane16_strm1_data_valid ),      
               .std__pe47__lane16_strm1_data_mask     ( std__pe47__lane16_strm1_data_mask  ),      

               // PE 47, Lane 17                 
               .pe47__std__lane17_strm0_ready         ( pe47__std__lane17_strm0_ready      ),      
               .std__pe47__lane17_strm0_cntl          ( std__pe47__lane17_strm0_cntl       ),      
               .std__pe47__lane17_strm0_data          ( std__pe47__lane17_strm0_data       ),      
               .std__pe47__lane17_strm0_data_valid    ( std__pe47__lane17_strm0_data_valid ),      
               .std__pe47__lane17_strm0_data_mask     ( std__pe47__lane17_strm0_data_mask  ),      

               .pe47__std__lane17_strm1_ready         ( pe47__std__lane17_strm1_ready      ),      
               .std__pe47__lane17_strm1_cntl          ( std__pe47__lane17_strm1_cntl       ),      
               .std__pe47__lane17_strm1_data          ( std__pe47__lane17_strm1_data       ),      
               .std__pe47__lane17_strm1_data_valid    ( std__pe47__lane17_strm1_data_valid ),      
               .std__pe47__lane17_strm1_data_mask     ( std__pe47__lane17_strm1_data_mask  ),      

               // PE 47, Lane 18                 
               .pe47__std__lane18_strm0_ready         ( pe47__std__lane18_strm0_ready      ),      
               .std__pe47__lane18_strm0_cntl          ( std__pe47__lane18_strm0_cntl       ),      
               .std__pe47__lane18_strm0_data          ( std__pe47__lane18_strm0_data       ),      
               .std__pe47__lane18_strm0_data_valid    ( std__pe47__lane18_strm0_data_valid ),      
               .std__pe47__lane18_strm0_data_mask     ( std__pe47__lane18_strm0_data_mask  ),      

               .pe47__std__lane18_strm1_ready         ( pe47__std__lane18_strm1_ready      ),      
               .std__pe47__lane18_strm1_cntl          ( std__pe47__lane18_strm1_cntl       ),      
               .std__pe47__lane18_strm1_data          ( std__pe47__lane18_strm1_data       ),      
               .std__pe47__lane18_strm1_data_valid    ( std__pe47__lane18_strm1_data_valid ),      
               .std__pe47__lane18_strm1_data_mask     ( std__pe47__lane18_strm1_data_mask  ),      

               // PE 47, Lane 19                 
               .pe47__std__lane19_strm0_ready         ( pe47__std__lane19_strm0_ready      ),      
               .std__pe47__lane19_strm0_cntl          ( std__pe47__lane19_strm0_cntl       ),      
               .std__pe47__lane19_strm0_data          ( std__pe47__lane19_strm0_data       ),      
               .std__pe47__lane19_strm0_data_valid    ( std__pe47__lane19_strm0_data_valid ),      
               .std__pe47__lane19_strm0_data_mask     ( std__pe47__lane19_strm0_data_mask  ),      

               .pe47__std__lane19_strm1_ready         ( pe47__std__lane19_strm1_ready      ),      
               .std__pe47__lane19_strm1_cntl          ( std__pe47__lane19_strm1_cntl       ),      
               .std__pe47__lane19_strm1_data          ( std__pe47__lane19_strm1_data       ),      
               .std__pe47__lane19_strm1_data_valid    ( std__pe47__lane19_strm1_data_valid ),      
               .std__pe47__lane19_strm1_data_mask     ( std__pe47__lane19_strm1_data_mask  ),      

               // PE 47, Lane 20                 
               .pe47__std__lane20_strm0_ready         ( pe47__std__lane20_strm0_ready      ),      
               .std__pe47__lane20_strm0_cntl          ( std__pe47__lane20_strm0_cntl       ),      
               .std__pe47__lane20_strm0_data          ( std__pe47__lane20_strm0_data       ),      
               .std__pe47__lane20_strm0_data_valid    ( std__pe47__lane20_strm0_data_valid ),      
               .std__pe47__lane20_strm0_data_mask     ( std__pe47__lane20_strm0_data_mask  ),      

               .pe47__std__lane20_strm1_ready         ( pe47__std__lane20_strm1_ready      ),      
               .std__pe47__lane20_strm1_cntl          ( std__pe47__lane20_strm1_cntl       ),      
               .std__pe47__lane20_strm1_data          ( std__pe47__lane20_strm1_data       ),      
               .std__pe47__lane20_strm1_data_valid    ( std__pe47__lane20_strm1_data_valid ),      
               .std__pe47__lane20_strm1_data_mask     ( std__pe47__lane20_strm1_data_mask  ),      

               // PE 47, Lane 21                 
               .pe47__std__lane21_strm0_ready         ( pe47__std__lane21_strm0_ready      ),      
               .std__pe47__lane21_strm0_cntl          ( std__pe47__lane21_strm0_cntl       ),      
               .std__pe47__lane21_strm0_data          ( std__pe47__lane21_strm0_data       ),      
               .std__pe47__lane21_strm0_data_valid    ( std__pe47__lane21_strm0_data_valid ),      
               .std__pe47__lane21_strm0_data_mask     ( std__pe47__lane21_strm0_data_mask  ),      

               .pe47__std__lane21_strm1_ready         ( pe47__std__lane21_strm1_ready      ),      
               .std__pe47__lane21_strm1_cntl          ( std__pe47__lane21_strm1_cntl       ),      
               .std__pe47__lane21_strm1_data          ( std__pe47__lane21_strm1_data       ),      
               .std__pe47__lane21_strm1_data_valid    ( std__pe47__lane21_strm1_data_valid ),      
               .std__pe47__lane21_strm1_data_mask     ( std__pe47__lane21_strm1_data_mask  ),      

               // PE 47, Lane 22                 
               .pe47__std__lane22_strm0_ready         ( pe47__std__lane22_strm0_ready      ),      
               .std__pe47__lane22_strm0_cntl          ( std__pe47__lane22_strm0_cntl       ),      
               .std__pe47__lane22_strm0_data          ( std__pe47__lane22_strm0_data       ),      
               .std__pe47__lane22_strm0_data_valid    ( std__pe47__lane22_strm0_data_valid ),      
               .std__pe47__lane22_strm0_data_mask     ( std__pe47__lane22_strm0_data_mask  ),      

               .pe47__std__lane22_strm1_ready         ( pe47__std__lane22_strm1_ready      ),      
               .std__pe47__lane22_strm1_cntl          ( std__pe47__lane22_strm1_cntl       ),      
               .std__pe47__lane22_strm1_data          ( std__pe47__lane22_strm1_data       ),      
               .std__pe47__lane22_strm1_data_valid    ( std__pe47__lane22_strm1_data_valid ),      
               .std__pe47__lane22_strm1_data_mask     ( std__pe47__lane22_strm1_data_mask  ),      

               // PE 47, Lane 23                 
               .pe47__std__lane23_strm0_ready         ( pe47__std__lane23_strm0_ready      ),      
               .std__pe47__lane23_strm0_cntl          ( std__pe47__lane23_strm0_cntl       ),      
               .std__pe47__lane23_strm0_data          ( std__pe47__lane23_strm0_data       ),      
               .std__pe47__lane23_strm0_data_valid    ( std__pe47__lane23_strm0_data_valid ),      
               .std__pe47__lane23_strm0_data_mask     ( std__pe47__lane23_strm0_data_mask  ),      

               .pe47__std__lane23_strm1_ready         ( pe47__std__lane23_strm1_ready      ),      
               .std__pe47__lane23_strm1_cntl          ( std__pe47__lane23_strm1_cntl       ),      
               .std__pe47__lane23_strm1_data          ( std__pe47__lane23_strm1_data       ),      
               .std__pe47__lane23_strm1_data_valid    ( std__pe47__lane23_strm1_data_valid ),      
               .std__pe47__lane23_strm1_data_mask     ( std__pe47__lane23_strm1_data_mask  ),      

               // PE 47, Lane 24                 
               .pe47__std__lane24_strm0_ready         ( pe47__std__lane24_strm0_ready      ),      
               .std__pe47__lane24_strm0_cntl          ( std__pe47__lane24_strm0_cntl       ),      
               .std__pe47__lane24_strm0_data          ( std__pe47__lane24_strm0_data       ),      
               .std__pe47__lane24_strm0_data_valid    ( std__pe47__lane24_strm0_data_valid ),      
               .std__pe47__lane24_strm0_data_mask     ( std__pe47__lane24_strm0_data_mask  ),      

               .pe47__std__lane24_strm1_ready         ( pe47__std__lane24_strm1_ready      ),      
               .std__pe47__lane24_strm1_cntl          ( std__pe47__lane24_strm1_cntl       ),      
               .std__pe47__lane24_strm1_data          ( std__pe47__lane24_strm1_data       ),      
               .std__pe47__lane24_strm1_data_valid    ( std__pe47__lane24_strm1_data_valid ),      
               .std__pe47__lane24_strm1_data_mask     ( std__pe47__lane24_strm1_data_mask  ),      

               // PE 47, Lane 25                 
               .pe47__std__lane25_strm0_ready         ( pe47__std__lane25_strm0_ready      ),      
               .std__pe47__lane25_strm0_cntl          ( std__pe47__lane25_strm0_cntl       ),      
               .std__pe47__lane25_strm0_data          ( std__pe47__lane25_strm0_data       ),      
               .std__pe47__lane25_strm0_data_valid    ( std__pe47__lane25_strm0_data_valid ),      
               .std__pe47__lane25_strm0_data_mask     ( std__pe47__lane25_strm0_data_mask  ),      

               .pe47__std__lane25_strm1_ready         ( pe47__std__lane25_strm1_ready      ),      
               .std__pe47__lane25_strm1_cntl          ( std__pe47__lane25_strm1_cntl       ),      
               .std__pe47__lane25_strm1_data          ( std__pe47__lane25_strm1_data       ),      
               .std__pe47__lane25_strm1_data_valid    ( std__pe47__lane25_strm1_data_valid ),      
               .std__pe47__lane25_strm1_data_mask     ( std__pe47__lane25_strm1_data_mask  ),      

               // PE 47, Lane 26                 
               .pe47__std__lane26_strm0_ready         ( pe47__std__lane26_strm0_ready      ),      
               .std__pe47__lane26_strm0_cntl          ( std__pe47__lane26_strm0_cntl       ),      
               .std__pe47__lane26_strm0_data          ( std__pe47__lane26_strm0_data       ),      
               .std__pe47__lane26_strm0_data_valid    ( std__pe47__lane26_strm0_data_valid ),      
               .std__pe47__lane26_strm0_data_mask     ( std__pe47__lane26_strm0_data_mask  ),      

               .pe47__std__lane26_strm1_ready         ( pe47__std__lane26_strm1_ready      ),      
               .std__pe47__lane26_strm1_cntl          ( std__pe47__lane26_strm1_cntl       ),      
               .std__pe47__lane26_strm1_data          ( std__pe47__lane26_strm1_data       ),      
               .std__pe47__lane26_strm1_data_valid    ( std__pe47__lane26_strm1_data_valid ),      
               .std__pe47__lane26_strm1_data_mask     ( std__pe47__lane26_strm1_data_mask  ),      

               // PE 47, Lane 27                 
               .pe47__std__lane27_strm0_ready         ( pe47__std__lane27_strm0_ready      ),      
               .std__pe47__lane27_strm0_cntl          ( std__pe47__lane27_strm0_cntl       ),      
               .std__pe47__lane27_strm0_data          ( std__pe47__lane27_strm0_data       ),      
               .std__pe47__lane27_strm0_data_valid    ( std__pe47__lane27_strm0_data_valid ),      
               .std__pe47__lane27_strm0_data_mask     ( std__pe47__lane27_strm0_data_mask  ),      

               .pe47__std__lane27_strm1_ready         ( pe47__std__lane27_strm1_ready      ),      
               .std__pe47__lane27_strm1_cntl          ( std__pe47__lane27_strm1_cntl       ),      
               .std__pe47__lane27_strm1_data          ( std__pe47__lane27_strm1_data       ),      
               .std__pe47__lane27_strm1_data_valid    ( std__pe47__lane27_strm1_data_valid ),      
               .std__pe47__lane27_strm1_data_mask     ( std__pe47__lane27_strm1_data_mask  ),      

               // PE 47, Lane 28                 
               .pe47__std__lane28_strm0_ready         ( pe47__std__lane28_strm0_ready      ),      
               .std__pe47__lane28_strm0_cntl          ( std__pe47__lane28_strm0_cntl       ),      
               .std__pe47__lane28_strm0_data          ( std__pe47__lane28_strm0_data       ),      
               .std__pe47__lane28_strm0_data_valid    ( std__pe47__lane28_strm0_data_valid ),      
               .std__pe47__lane28_strm0_data_mask     ( std__pe47__lane28_strm0_data_mask  ),      

               .pe47__std__lane28_strm1_ready         ( pe47__std__lane28_strm1_ready      ),      
               .std__pe47__lane28_strm1_cntl          ( std__pe47__lane28_strm1_cntl       ),      
               .std__pe47__lane28_strm1_data          ( std__pe47__lane28_strm1_data       ),      
               .std__pe47__lane28_strm1_data_valid    ( std__pe47__lane28_strm1_data_valid ),      
               .std__pe47__lane28_strm1_data_mask     ( std__pe47__lane28_strm1_data_mask  ),      

               // PE 47, Lane 29                 
               .pe47__std__lane29_strm0_ready         ( pe47__std__lane29_strm0_ready      ),      
               .std__pe47__lane29_strm0_cntl          ( std__pe47__lane29_strm0_cntl       ),      
               .std__pe47__lane29_strm0_data          ( std__pe47__lane29_strm0_data       ),      
               .std__pe47__lane29_strm0_data_valid    ( std__pe47__lane29_strm0_data_valid ),      
               .std__pe47__lane29_strm0_data_mask     ( std__pe47__lane29_strm0_data_mask  ),      

               .pe47__std__lane29_strm1_ready         ( pe47__std__lane29_strm1_ready      ),      
               .std__pe47__lane29_strm1_cntl          ( std__pe47__lane29_strm1_cntl       ),      
               .std__pe47__lane29_strm1_data          ( std__pe47__lane29_strm1_data       ),      
               .std__pe47__lane29_strm1_data_valid    ( std__pe47__lane29_strm1_data_valid ),      
               .std__pe47__lane29_strm1_data_mask     ( std__pe47__lane29_strm1_data_mask  ),      

               // PE 47, Lane 30                 
               .pe47__std__lane30_strm0_ready         ( pe47__std__lane30_strm0_ready      ),      
               .std__pe47__lane30_strm0_cntl          ( std__pe47__lane30_strm0_cntl       ),      
               .std__pe47__lane30_strm0_data          ( std__pe47__lane30_strm0_data       ),      
               .std__pe47__lane30_strm0_data_valid    ( std__pe47__lane30_strm0_data_valid ),      
               .std__pe47__lane30_strm0_data_mask     ( std__pe47__lane30_strm0_data_mask  ),      

               .pe47__std__lane30_strm1_ready         ( pe47__std__lane30_strm1_ready      ),      
               .std__pe47__lane30_strm1_cntl          ( std__pe47__lane30_strm1_cntl       ),      
               .std__pe47__lane30_strm1_data          ( std__pe47__lane30_strm1_data       ),      
               .std__pe47__lane30_strm1_data_valid    ( std__pe47__lane30_strm1_data_valid ),      
               .std__pe47__lane30_strm1_data_mask     ( std__pe47__lane30_strm1_data_mask  ),      

               // PE 47, Lane 31                 
               .pe47__std__lane31_strm0_ready         ( pe47__std__lane31_strm0_ready      ),      
               .std__pe47__lane31_strm0_cntl          ( std__pe47__lane31_strm0_cntl       ),      
               .std__pe47__lane31_strm0_data          ( std__pe47__lane31_strm0_data       ),      
               .std__pe47__lane31_strm0_data_valid    ( std__pe47__lane31_strm0_data_valid ),      
               .std__pe47__lane31_strm0_data_mask     ( std__pe47__lane31_strm0_data_mask  ),      

               .pe47__std__lane31_strm1_ready         ( pe47__std__lane31_strm1_ready      ),      
               .std__pe47__lane31_strm1_cntl          ( std__pe47__lane31_strm1_cntl       ),      
               .std__pe47__lane31_strm1_data          ( std__pe47__lane31_strm1_data       ),      
               .std__pe47__lane31_strm1_data_valid    ( std__pe47__lane31_strm1_data_valid ),      
               .std__pe47__lane31_strm1_data_mask     ( std__pe47__lane31_strm1_data_mask  ),      

               // PE 48, Lane 0                 
               .pe48__std__lane0_strm0_ready         ( pe48__std__lane0_strm0_ready      ),      
               .std__pe48__lane0_strm0_cntl          ( std__pe48__lane0_strm0_cntl       ),      
               .std__pe48__lane0_strm0_data          ( std__pe48__lane0_strm0_data       ),      
               .std__pe48__lane0_strm0_data_valid    ( std__pe48__lane0_strm0_data_valid ),      
               .std__pe48__lane0_strm0_data_mask     ( std__pe48__lane0_strm0_data_mask  ),      

               .pe48__std__lane0_strm1_ready         ( pe48__std__lane0_strm1_ready      ),      
               .std__pe48__lane0_strm1_cntl          ( std__pe48__lane0_strm1_cntl       ),      
               .std__pe48__lane0_strm1_data          ( std__pe48__lane0_strm1_data       ),      
               .std__pe48__lane0_strm1_data_valid    ( std__pe48__lane0_strm1_data_valid ),      
               .std__pe48__lane0_strm1_data_mask     ( std__pe48__lane0_strm1_data_mask  ),      

               // PE 48, Lane 1                 
               .pe48__std__lane1_strm0_ready         ( pe48__std__lane1_strm0_ready      ),      
               .std__pe48__lane1_strm0_cntl          ( std__pe48__lane1_strm0_cntl       ),      
               .std__pe48__lane1_strm0_data          ( std__pe48__lane1_strm0_data       ),      
               .std__pe48__lane1_strm0_data_valid    ( std__pe48__lane1_strm0_data_valid ),      
               .std__pe48__lane1_strm0_data_mask     ( std__pe48__lane1_strm0_data_mask  ),      

               .pe48__std__lane1_strm1_ready         ( pe48__std__lane1_strm1_ready      ),      
               .std__pe48__lane1_strm1_cntl          ( std__pe48__lane1_strm1_cntl       ),      
               .std__pe48__lane1_strm1_data          ( std__pe48__lane1_strm1_data       ),      
               .std__pe48__lane1_strm1_data_valid    ( std__pe48__lane1_strm1_data_valid ),      
               .std__pe48__lane1_strm1_data_mask     ( std__pe48__lane1_strm1_data_mask  ),      

               // PE 48, Lane 2                 
               .pe48__std__lane2_strm0_ready         ( pe48__std__lane2_strm0_ready      ),      
               .std__pe48__lane2_strm0_cntl          ( std__pe48__lane2_strm0_cntl       ),      
               .std__pe48__lane2_strm0_data          ( std__pe48__lane2_strm0_data       ),      
               .std__pe48__lane2_strm0_data_valid    ( std__pe48__lane2_strm0_data_valid ),      
               .std__pe48__lane2_strm0_data_mask     ( std__pe48__lane2_strm0_data_mask  ),      

               .pe48__std__lane2_strm1_ready         ( pe48__std__lane2_strm1_ready      ),      
               .std__pe48__lane2_strm1_cntl          ( std__pe48__lane2_strm1_cntl       ),      
               .std__pe48__lane2_strm1_data          ( std__pe48__lane2_strm1_data       ),      
               .std__pe48__lane2_strm1_data_valid    ( std__pe48__lane2_strm1_data_valid ),      
               .std__pe48__lane2_strm1_data_mask     ( std__pe48__lane2_strm1_data_mask  ),      

               // PE 48, Lane 3                 
               .pe48__std__lane3_strm0_ready         ( pe48__std__lane3_strm0_ready      ),      
               .std__pe48__lane3_strm0_cntl          ( std__pe48__lane3_strm0_cntl       ),      
               .std__pe48__lane3_strm0_data          ( std__pe48__lane3_strm0_data       ),      
               .std__pe48__lane3_strm0_data_valid    ( std__pe48__lane3_strm0_data_valid ),      
               .std__pe48__lane3_strm0_data_mask     ( std__pe48__lane3_strm0_data_mask  ),      

               .pe48__std__lane3_strm1_ready         ( pe48__std__lane3_strm1_ready      ),      
               .std__pe48__lane3_strm1_cntl          ( std__pe48__lane3_strm1_cntl       ),      
               .std__pe48__lane3_strm1_data          ( std__pe48__lane3_strm1_data       ),      
               .std__pe48__lane3_strm1_data_valid    ( std__pe48__lane3_strm1_data_valid ),      
               .std__pe48__lane3_strm1_data_mask     ( std__pe48__lane3_strm1_data_mask  ),      

               // PE 48, Lane 4                 
               .pe48__std__lane4_strm0_ready         ( pe48__std__lane4_strm0_ready      ),      
               .std__pe48__lane4_strm0_cntl          ( std__pe48__lane4_strm0_cntl       ),      
               .std__pe48__lane4_strm0_data          ( std__pe48__lane4_strm0_data       ),      
               .std__pe48__lane4_strm0_data_valid    ( std__pe48__lane4_strm0_data_valid ),      
               .std__pe48__lane4_strm0_data_mask     ( std__pe48__lane4_strm0_data_mask  ),      

               .pe48__std__lane4_strm1_ready         ( pe48__std__lane4_strm1_ready      ),      
               .std__pe48__lane4_strm1_cntl          ( std__pe48__lane4_strm1_cntl       ),      
               .std__pe48__lane4_strm1_data          ( std__pe48__lane4_strm1_data       ),      
               .std__pe48__lane4_strm1_data_valid    ( std__pe48__lane4_strm1_data_valid ),      
               .std__pe48__lane4_strm1_data_mask     ( std__pe48__lane4_strm1_data_mask  ),      

               // PE 48, Lane 5                 
               .pe48__std__lane5_strm0_ready         ( pe48__std__lane5_strm0_ready      ),      
               .std__pe48__lane5_strm0_cntl          ( std__pe48__lane5_strm0_cntl       ),      
               .std__pe48__lane5_strm0_data          ( std__pe48__lane5_strm0_data       ),      
               .std__pe48__lane5_strm0_data_valid    ( std__pe48__lane5_strm0_data_valid ),      
               .std__pe48__lane5_strm0_data_mask     ( std__pe48__lane5_strm0_data_mask  ),      

               .pe48__std__lane5_strm1_ready         ( pe48__std__lane5_strm1_ready      ),      
               .std__pe48__lane5_strm1_cntl          ( std__pe48__lane5_strm1_cntl       ),      
               .std__pe48__lane5_strm1_data          ( std__pe48__lane5_strm1_data       ),      
               .std__pe48__lane5_strm1_data_valid    ( std__pe48__lane5_strm1_data_valid ),      
               .std__pe48__lane5_strm1_data_mask     ( std__pe48__lane5_strm1_data_mask  ),      

               // PE 48, Lane 6                 
               .pe48__std__lane6_strm0_ready         ( pe48__std__lane6_strm0_ready      ),      
               .std__pe48__lane6_strm0_cntl          ( std__pe48__lane6_strm0_cntl       ),      
               .std__pe48__lane6_strm0_data          ( std__pe48__lane6_strm0_data       ),      
               .std__pe48__lane6_strm0_data_valid    ( std__pe48__lane6_strm0_data_valid ),      
               .std__pe48__lane6_strm0_data_mask     ( std__pe48__lane6_strm0_data_mask  ),      

               .pe48__std__lane6_strm1_ready         ( pe48__std__lane6_strm1_ready      ),      
               .std__pe48__lane6_strm1_cntl          ( std__pe48__lane6_strm1_cntl       ),      
               .std__pe48__lane6_strm1_data          ( std__pe48__lane6_strm1_data       ),      
               .std__pe48__lane6_strm1_data_valid    ( std__pe48__lane6_strm1_data_valid ),      
               .std__pe48__lane6_strm1_data_mask     ( std__pe48__lane6_strm1_data_mask  ),      

               // PE 48, Lane 7                 
               .pe48__std__lane7_strm0_ready         ( pe48__std__lane7_strm0_ready      ),      
               .std__pe48__lane7_strm0_cntl          ( std__pe48__lane7_strm0_cntl       ),      
               .std__pe48__lane7_strm0_data          ( std__pe48__lane7_strm0_data       ),      
               .std__pe48__lane7_strm0_data_valid    ( std__pe48__lane7_strm0_data_valid ),      
               .std__pe48__lane7_strm0_data_mask     ( std__pe48__lane7_strm0_data_mask  ),      

               .pe48__std__lane7_strm1_ready         ( pe48__std__lane7_strm1_ready      ),      
               .std__pe48__lane7_strm1_cntl          ( std__pe48__lane7_strm1_cntl       ),      
               .std__pe48__lane7_strm1_data          ( std__pe48__lane7_strm1_data       ),      
               .std__pe48__lane7_strm1_data_valid    ( std__pe48__lane7_strm1_data_valid ),      
               .std__pe48__lane7_strm1_data_mask     ( std__pe48__lane7_strm1_data_mask  ),      

               // PE 48, Lane 8                 
               .pe48__std__lane8_strm0_ready         ( pe48__std__lane8_strm0_ready      ),      
               .std__pe48__lane8_strm0_cntl          ( std__pe48__lane8_strm0_cntl       ),      
               .std__pe48__lane8_strm0_data          ( std__pe48__lane8_strm0_data       ),      
               .std__pe48__lane8_strm0_data_valid    ( std__pe48__lane8_strm0_data_valid ),      
               .std__pe48__lane8_strm0_data_mask     ( std__pe48__lane8_strm0_data_mask  ),      

               .pe48__std__lane8_strm1_ready         ( pe48__std__lane8_strm1_ready      ),      
               .std__pe48__lane8_strm1_cntl          ( std__pe48__lane8_strm1_cntl       ),      
               .std__pe48__lane8_strm1_data          ( std__pe48__lane8_strm1_data       ),      
               .std__pe48__lane8_strm1_data_valid    ( std__pe48__lane8_strm1_data_valid ),      
               .std__pe48__lane8_strm1_data_mask     ( std__pe48__lane8_strm1_data_mask  ),      

               // PE 48, Lane 9                 
               .pe48__std__lane9_strm0_ready         ( pe48__std__lane9_strm0_ready      ),      
               .std__pe48__lane9_strm0_cntl          ( std__pe48__lane9_strm0_cntl       ),      
               .std__pe48__lane9_strm0_data          ( std__pe48__lane9_strm0_data       ),      
               .std__pe48__lane9_strm0_data_valid    ( std__pe48__lane9_strm0_data_valid ),      
               .std__pe48__lane9_strm0_data_mask     ( std__pe48__lane9_strm0_data_mask  ),      

               .pe48__std__lane9_strm1_ready         ( pe48__std__lane9_strm1_ready      ),      
               .std__pe48__lane9_strm1_cntl          ( std__pe48__lane9_strm1_cntl       ),      
               .std__pe48__lane9_strm1_data          ( std__pe48__lane9_strm1_data       ),      
               .std__pe48__lane9_strm1_data_valid    ( std__pe48__lane9_strm1_data_valid ),      
               .std__pe48__lane9_strm1_data_mask     ( std__pe48__lane9_strm1_data_mask  ),      

               // PE 48, Lane 10                 
               .pe48__std__lane10_strm0_ready         ( pe48__std__lane10_strm0_ready      ),      
               .std__pe48__lane10_strm0_cntl          ( std__pe48__lane10_strm0_cntl       ),      
               .std__pe48__lane10_strm0_data          ( std__pe48__lane10_strm0_data       ),      
               .std__pe48__lane10_strm0_data_valid    ( std__pe48__lane10_strm0_data_valid ),      
               .std__pe48__lane10_strm0_data_mask     ( std__pe48__lane10_strm0_data_mask  ),      

               .pe48__std__lane10_strm1_ready         ( pe48__std__lane10_strm1_ready      ),      
               .std__pe48__lane10_strm1_cntl          ( std__pe48__lane10_strm1_cntl       ),      
               .std__pe48__lane10_strm1_data          ( std__pe48__lane10_strm1_data       ),      
               .std__pe48__lane10_strm1_data_valid    ( std__pe48__lane10_strm1_data_valid ),      
               .std__pe48__lane10_strm1_data_mask     ( std__pe48__lane10_strm1_data_mask  ),      

               // PE 48, Lane 11                 
               .pe48__std__lane11_strm0_ready         ( pe48__std__lane11_strm0_ready      ),      
               .std__pe48__lane11_strm0_cntl          ( std__pe48__lane11_strm0_cntl       ),      
               .std__pe48__lane11_strm0_data          ( std__pe48__lane11_strm0_data       ),      
               .std__pe48__lane11_strm0_data_valid    ( std__pe48__lane11_strm0_data_valid ),      
               .std__pe48__lane11_strm0_data_mask     ( std__pe48__lane11_strm0_data_mask  ),      

               .pe48__std__lane11_strm1_ready         ( pe48__std__lane11_strm1_ready      ),      
               .std__pe48__lane11_strm1_cntl          ( std__pe48__lane11_strm1_cntl       ),      
               .std__pe48__lane11_strm1_data          ( std__pe48__lane11_strm1_data       ),      
               .std__pe48__lane11_strm1_data_valid    ( std__pe48__lane11_strm1_data_valid ),      
               .std__pe48__lane11_strm1_data_mask     ( std__pe48__lane11_strm1_data_mask  ),      

               // PE 48, Lane 12                 
               .pe48__std__lane12_strm0_ready         ( pe48__std__lane12_strm0_ready      ),      
               .std__pe48__lane12_strm0_cntl          ( std__pe48__lane12_strm0_cntl       ),      
               .std__pe48__lane12_strm0_data          ( std__pe48__lane12_strm0_data       ),      
               .std__pe48__lane12_strm0_data_valid    ( std__pe48__lane12_strm0_data_valid ),      
               .std__pe48__lane12_strm0_data_mask     ( std__pe48__lane12_strm0_data_mask  ),      

               .pe48__std__lane12_strm1_ready         ( pe48__std__lane12_strm1_ready      ),      
               .std__pe48__lane12_strm1_cntl          ( std__pe48__lane12_strm1_cntl       ),      
               .std__pe48__lane12_strm1_data          ( std__pe48__lane12_strm1_data       ),      
               .std__pe48__lane12_strm1_data_valid    ( std__pe48__lane12_strm1_data_valid ),      
               .std__pe48__lane12_strm1_data_mask     ( std__pe48__lane12_strm1_data_mask  ),      

               // PE 48, Lane 13                 
               .pe48__std__lane13_strm0_ready         ( pe48__std__lane13_strm0_ready      ),      
               .std__pe48__lane13_strm0_cntl          ( std__pe48__lane13_strm0_cntl       ),      
               .std__pe48__lane13_strm0_data          ( std__pe48__lane13_strm0_data       ),      
               .std__pe48__lane13_strm0_data_valid    ( std__pe48__lane13_strm0_data_valid ),      
               .std__pe48__lane13_strm0_data_mask     ( std__pe48__lane13_strm0_data_mask  ),      

               .pe48__std__lane13_strm1_ready         ( pe48__std__lane13_strm1_ready      ),      
               .std__pe48__lane13_strm1_cntl          ( std__pe48__lane13_strm1_cntl       ),      
               .std__pe48__lane13_strm1_data          ( std__pe48__lane13_strm1_data       ),      
               .std__pe48__lane13_strm1_data_valid    ( std__pe48__lane13_strm1_data_valid ),      
               .std__pe48__lane13_strm1_data_mask     ( std__pe48__lane13_strm1_data_mask  ),      

               // PE 48, Lane 14                 
               .pe48__std__lane14_strm0_ready         ( pe48__std__lane14_strm0_ready      ),      
               .std__pe48__lane14_strm0_cntl          ( std__pe48__lane14_strm0_cntl       ),      
               .std__pe48__lane14_strm0_data          ( std__pe48__lane14_strm0_data       ),      
               .std__pe48__lane14_strm0_data_valid    ( std__pe48__lane14_strm0_data_valid ),      
               .std__pe48__lane14_strm0_data_mask     ( std__pe48__lane14_strm0_data_mask  ),      

               .pe48__std__lane14_strm1_ready         ( pe48__std__lane14_strm1_ready      ),      
               .std__pe48__lane14_strm1_cntl          ( std__pe48__lane14_strm1_cntl       ),      
               .std__pe48__lane14_strm1_data          ( std__pe48__lane14_strm1_data       ),      
               .std__pe48__lane14_strm1_data_valid    ( std__pe48__lane14_strm1_data_valid ),      
               .std__pe48__lane14_strm1_data_mask     ( std__pe48__lane14_strm1_data_mask  ),      

               // PE 48, Lane 15                 
               .pe48__std__lane15_strm0_ready         ( pe48__std__lane15_strm0_ready      ),      
               .std__pe48__lane15_strm0_cntl          ( std__pe48__lane15_strm0_cntl       ),      
               .std__pe48__lane15_strm0_data          ( std__pe48__lane15_strm0_data       ),      
               .std__pe48__lane15_strm0_data_valid    ( std__pe48__lane15_strm0_data_valid ),      
               .std__pe48__lane15_strm0_data_mask     ( std__pe48__lane15_strm0_data_mask  ),      

               .pe48__std__lane15_strm1_ready         ( pe48__std__lane15_strm1_ready      ),      
               .std__pe48__lane15_strm1_cntl          ( std__pe48__lane15_strm1_cntl       ),      
               .std__pe48__lane15_strm1_data          ( std__pe48__lane15_strm1_data       ),      
               .std__pe48__lane15_strm1_data_valid    ( std__pe48__lane15_strm1_data_valid ),      
               .std__pe48__lane15_strm1_data_mask     ( std__pe48__lane15_strm1_data_mask  ),      

               // PE 48, Lane 16                 
               .pe48__std__lane16_strm0_ready         ( pe48__std__lane16_strm0_ready      ),      
               .std__pe48__lane16_strm0_cntl          ( std__pe48__lane16_strm0_cntl       ),      
               .std__pe48__lane16_strm0_data          ( std__pe48__lane16_strm0_data       ),      
               .std__pe48__lane16_strm0_data_valid    ( std__pe48__lane16_strm0_data_valid ),      
               .std__pe48__lane16_strm0_data_mask     ( std__pe48__lane16_strm0_data_mask  ),      

               .pe48__std__lane16_strm1_ready         ( pe48__std__lane16_strm1_ready      ),      
               .std__pe48__lane16_strm1_cntl          ( std__pe48__lane16_strm1_cntl       ),      
               .std__pe48__lane16_strm1_data          ( std__pe48__lane16_strm1_data       ),      
               .std__pe48__lane16_strm1_data_valid    ( std__pe48__lane16_strm1_data_valid ),      
               .std__pe48__lane16_strm1_data_mask     ( std__pe48__lane16_strm1_data_mask  ),      

               // PE 48, Lane 17                 
               .pe48__std__lane17_strm0_ready         ( pe48__std__lane17_strm0_ready      ),      
               .std__pe48__lane17_strm0_cntl          ( std__pe48__lane17_strm0_cntl       ),      
               .std__pe48__lane17_strm0_data          ( std__pe48__lane17_strm0_data       ),      
               .std__pe48__lane17_strm0_data_valid    ( std__pe48__lane17_strm0_data_valid ),      
               .std__pe48__lane17_strm0_data_mask     ( std__pe48__lane17_strm0_data_mask  ),      

               .pe48__std__lane17_strm1_ready         ( pe48__std__lane17_strm1_ready      ),      
               .std__pe48__lane17_strm1_cntl          ( std__pe48__lane17_strm1_cntl       ),      
               .std__pe48__lane17_strm1_data          ( std__pe48__lane17_strm1_data       ),      
               .std__pe48__lane17_strm1_data_valid    ( std__pe48__lane17_strm1_data_valid ),      
               .std__pe48__lane17_strm1_data_mask     ( std__pe48__lane17_strm1_data_mask  ),      

               // PE 48, Lane 18                 
               .pe48__std__lane18_strm0_ready         ( pe48__std__lane18_strm0_ready      ),      
               .std__pe48__lane18_strm0_cntl          ( std__pe48__lane18_strm0_cntl       ),      
               .std__pe48__lane18_strm0_data          ( std__pe48__lane18_strm0_data       ),      
               .std__pe48__lane18_strm0_data_valid    ( std__pe48__lane18_strm0_data_valid ),      
               .std__pe48__lane18_strm0_data_mask     ( std__pe48__lane18_strm0_data_mask  ),      

               .pe48__std__lane18_strm1_ready         ( pe48__std__lane18_strm1_ready      ),      
               .std__pe48__lane18_strm1_cntl          ( std__pe48__lane18_strm1_cntl       ),      
               .std__pe48__lane18_strm1_data          ( std__pe48__lane18_strm1_data       ),      
               .std__pe48__lane18_strm1_data_valid    ( std__pe48__lane18_strm1_data_valid ),      
               .std__pe48__lane18_strm1_data_mask     ( std__pe48__lane18_strm1_data_mask  ),      

               // PE 48, Lane 19                 
               .pe48__std__lane19_strm0_ready         ( pe48__std__lane19_strm0_ready      ),      
               .std__pe48__lane19_strm0_cntl          ( std__pe48__lane19_strm0_cntl       ),      
               .std__pe48__lane19_strm0_data          ( std__pe48__lane19_strm0_data       ),      
               .std__pe48__lane19_strm0_data_valid    ( std__pe48__lane19_strm0_data_valid ),      
               .std__pe48__lane19_strm0_data_mask     ( std__pe48__lane19_strm0_data_mask  ),      

               .pe48__std__lane19_strm1_ready         ( pe48__std__lane19_strm1_ready      ),      
               .std__pe48__lane19_strm1_cntl          ( std__pe48__lane19_strm1_cntl       ),      
               .std__pe48__lane19_strm1_data          ( std__pe48__lane19_strm1_data       ),      
               .std__pe48__lane19_strm1_data_valid    ( std__pe48__lane19_strm1_data_valid ),      
               .std__pe48__lane19_strm1_data_mask     ( std__pe48__lane19_strm1_data_mask  ),      

               // PE 48, Lane 20                 
               .pe48__std__lane20_strm0_ready         ( pe48__std__lane20_strm0_ready      ),      
               .std__pe48__lane20_strm0_cntl          ( std__pe48__lane20_strm0_cntl       ),      
               .std__pe48__lane20_strm0_data          ( std__pe48__lane20_strm0_data       ),      
               .std__pe48__lane20_strm0_data_valid    ( std__pe48__lane20_strm0_data_valid ),      
               .std__pe48__lane20_strm0_data_mask     ( std__pe48__lane20_strm0_data_mask  ),      

               .pe48__std__lane20_strm1_ready         ( pe48__std__lane20_strm1_ready      ),      
               .std__pe48__lane20_strm1_cntl          ( std__pe48__lane20_strm1_cntl       ),      
               .std__pe48__lane20_strm1_data          ( std__pe48__lane20_strm1_data       ),      
               .std__pe48__lane20_strm1_data_valid    ( std__pe48__lane20_strm1_data_valid ),      
               .std__pe48__lane20_strm1_data_mask     ( std__pe48__lane20_strm1_data_mask  ),      

               // PE 48, Lane 21                 
               .pe48__std__lane21_strm0_ready         ( pe48__std__lane21_strm0_ready      ),      
               .std__pe48__lane21_strm0_cntl          ( std__pe48__lane21_strm0_cntl       ),      
               .std__pe48__lane21_strm0_data          ( std__pe48__lane21_strm0_data       ),      
               .std__pe48__lane21_strm0_data_valid    ( std__pe48__lane21_strm0_data_valid ),      
               .std__pe48__lane21_strm0_data_mask     ( std__pe48__lane21_strm0_data_mask  ),      

               .pe48__std__lane21_strm1_ready         ( pe48__std__lane21_strm1_ready      ),      
               .std__pe48__lane21_strm1_cntl          ( std__pe48__lane21_strm1_cntl       ),      
               .std__pe48__lane21_strm1_data          ( std__pe48__lane21_strm1_data       ),      
               .std__pe48__lane21_strm1_data_valid    ( std__pe48__lane21_strm1_data_valid ),      
               .std__pe48__lane21_strm1_data_mask     ( std__pe48__lane21_strm1_data_mask  ),      

               // PE 48, Lane 22                 
               .pe48__std__lane22_strm0_ready         ( pe48__std__lane22_strm0_ready      ),      
               .std__pe48__lane22_strm0_cntl          ( std__pe48__lane22_strm0_cntl       ),      
               .std__pe48__lane22_strm0_data          ( std__pe48__lane22_strm0_data       ),      
               .std__pe48__lane22_strm0_data_valid    ( std__pe48__lane22_strm0_data_valid ),      
               .std__pe48__lane22_strm0_data_mask     ( std__pe48__lane22_strm0_data_mask  ),      

               .pe48__std__lane22_strm1_ready         ( pe48__std__lane22_strm1_ready      ),      
               .std__pe48__lane22_strm1_cntl          ( std__pe48__lane22_strm1_cntl       ),      
               .std__pe48__lane22_strm1_data          ( std__pe48__lane22_strm1_data       ),      
               .std__pe48__lane22_strm1_data_valid    ( std__pe48__lane22_strm1_data_valid ),      
               .std__pe48__lane22_strm1_data_mask     ( std__pe48__lane22_strm1_data_mask  ),      

               // PE 48, Lane 23                 
               .pe48__std__lane23_strm0_ready         ( pe48__std__lane23_strm0_ready      ),      
               .std__pe48__lane23_strm0_cntl          ( std__pe48__lane23_strm0_cntl       ),      
               .std__pe48__lane23_strm0_data          ( std__pe48__lane23_strm0_data       ),      
               .std__pe48__lane23_strm0_data_valid    ( std__pe48__lane23_strm0_data_valid ),      
               .std__pe48__lane23_strm0_data_mask     ( std__pe48__lane23_strm0_data_mask  ),      

               .pe48__std__lane23_strm1_ready         ( pe48__std__lane23_strm1_ready      ),      
               .std__pe48__lane23_strm1_cntl          ( std__pe48__lane23_strm1_cntl       ),      
               .std__pe48__lane23_strm1_data          ( std__pe48__lane23_strm1_data       ),      
               .std__pe48__lane23_strm1_data_valid    ( std__pe48__lane23_strm1_data_valid ),      
               .std__pe48__lane23_strm1_data_mask     ( std__pe48__lane23_strm1_data_mask  ),      

               // PE 48, Lane 24                 
               .pe48__std__lane24_strm0_ready         ( pe48__std__lane24_strm0_ready      ),      
               .std__pe48__lane24_strm0_cntl          ( std__pe48__lane24_strm0_cntl       ),      
               .std__pe48__lane24_strm0_data          ( std__pe48__lane24_strm0_data       ),      
               .std__pe48__lane24_strm0_data_valid    ( std__pe48__lane24_strm0_data_valid ),      
               .std__pe48__lane24_strm0_data_mask     ( std__pe48__lane24_strm0_data_mask  ),      

               .pe48__std__lane24_strm1_ready         ( pe48__std__lane24_strm1_ready      ),      
               .std__pe48__lane24_strm1_cntl          ( std__pe48__lane24_strm1_cntl       ),      
               .std__pe48__lane24_strm1_data          ( std__pe48__lane24_strm1_data       ),      
               .std__pe48__lane24_strm1_data_valid    ( std__pe48__lane24_strm1_data_valid ),      
               .std__pe48__lane24_strm1_data_mask     ( std__pe48__lane24_strm1_data_mask  ),      

               // PE 48, Lane 25                 
               .pe48__std__lane25_strm0_ready         ( pe48__std__lane25_strm0_ready      ),      
               .std__pe48__lane25_strm0_cntl          ( std__pe48__lane25_strm0_cntl       ),      
               .std__pe48__lane25_strm0_data          ( std__pe48__lane25_strm0_data       ),      
               .std__pe48__lane25_strm0_data_valid    ( std__pe48__lane25_strm0_data_valid ),      
               .std__pe48__lane25_strm0_data_mask     ( std__pe48__lane25_strm0_data_mask  ),      

               .pe48__std__lane25_strm1_ready         ( pe48__std__lane25_strm1_ready      ),      
               .std__pe48__lane25_strm1_cntl          ( std__pe48__lane25_strm1_cntl       ),      
               .std__pe48__lane25_strm1_data          ( std__pe48__lane25_strm1_data       ),      
               .std__pe48__lane25_strm1_data_valid    ( std__pe48__lane25_strm1_data_valid ),      
               .std__pe48__lane25_strm1_data_mask     ( std__pe48__lane25_strm1_data_mask  ),      

               // PE 48, Lane 26                 
               .pe48__std__lane26_strm0_ready         ( pe48__std__lane26_strm0_ready      ),      
               .std__pe48__lane26_strm0_cntl          ( std__pe48__lane26_strm0_cntl       ),      
               .std__pe48__lane26_strm0_data          ( std__pe48__lane26_strm0_data       ),      
               .std__pe48__lane26_strm0_data_valid    ( std__pe48__lane26_strm0_data_valid ),      
               .std__pe48__lane26_strm0_data_mask     ( std__pe48__lane26_strm0_data_mask  ),      

               .pe48__std__lane26_strm1_ready         ( pe48__std__lane26_strm1_ready      ),      
               .std__pe48__lane26_strm1_cntl          ( std__pe48__lane26_strm1_cntl       ),      
               .std__pe48__lane26_strm1_data          ( std__pe48__lane26_strm1_data       ),      
               .std__pe48__lane26_strm1_data_valid    ( std__pe48__lane26_strm1_data_valid ),      
               .std__pe48__lane26_strm1_data_mask     ( std__pe48__lane26_strm1_data_mask  ),      

               // PE 48, Lane 27                 
               .pe48__std__lane27_strm0_ready         ( pe48__std__lane27_strm0_ready      ),      
               .std__pe48__lane27_strm0_cntl          ( std__pe48__lane27_strm0_cntl       ),      
               .std__pe48__lane27_strm0_data          ( std__pe48__lane27_strm0_data       ),      
               .std__pe48__lane27_strm0_data_valid    ( std__pe48__lane27_strm0_data_valid ),      
               .std__pe48__lane27_strm0_data_mask     ( std__pe48__lane27_strm0_data_mask  ),      

               .pe48__std__lane27_strm1_ready         ( pe48__std__lane27_strm1_ready      ),      
               .std__pe48__lane27_strm1_cntl          ( std__pe48__lane27_strm1_cntl       ),      
               .std__pe48__lane27_strm1_data          ( std__pe48__lane27_strm1_data       ),      
               .std__pe48__lane27_strm1_data_valid    ( std__pe48__lane27_strm1_data_valid ),      
               .std__pe48__lane27_strm1_data_mask     ( std__pe48__lane27_strm1_data_mask  ),      

               // PE 48, Lane 28                 
               .pe48__std__lane28_strm0_ready         ( pe48__std__lane28_strm0_ready      ),      
               .std__pe48__lane28_strm0_cntl          ( std__pe48__lane28_strm0_cntl       ),      
               .std__pe48__lane28_strm0_data          ( std__pe48__lane28_strm0_data       ),      
               .std__pe48__lane28_strm0_data_valid    ( std__pe48__lane28_strm0_data_valid ),      
               .std__pe48__lane28_strm0_data_mask     ( std__pe48__lane28_strm0_data_mask  ),      

               .pe48__std__lane28_strm1_ready         ( pe48__std__lane28_strm1_ready      ),      
               .std__pe48__lane28_strm1_cntl          ( std__pe48__lane28_strm1_cntl       ),      
               .std__pe48__lane28_strm1_data          ( std__pe48__lane28_strm1_data       ),      
               .std__pe48__lane28_strm1_data_valid    ( std__pe48__lane28_strm1_data_valid ),      
               .std__pe48__lane28_strm1_data_mask     ( std__pe48__lane28_strm1_data_mask  ),      

               // PE 48, Lane 29                 
               .pe48__std__lane29_strm0_ready         ( pe48__std__lane29_strm0_ready      ),      
               .std__pe48__lane29_strm0_cntl          ( std__pe48__lane29_strm0_cntl       ),      
               .std__pe48__lane29_strm0_data          ( std__pe48__lane29_strm0_data       ),      
               .std__pe48__lane29_strm0_data_valid    ( std__pe48__lane29_strm0_data_valid ),      
               .std__pe48__lane29_strm0_data_mask     ( std__pe48__lane29_strm0_data_mask  ),      

               .pe48__std__lane29_strm1_ready         ( pe48__std__lane29_strm1_ready      ),      
               .std__pe48__lane29_strm1_cntl          ( std__pe48__lane29_strm1_cntl       ),      
               .std__pe48__lane29_strm1_data          ( std__pe48__lane29_strm1_data       ),      
               .std__pe48__lane29_strm1_data_valid    ( std__pe48__lane29_strm1_data_valid ),      
               .std__pe48__lane29_strm1_data_mask     ( std__pe48__lane29_strm1_data_mask  ),      

               // PE 48, Lane 30                 
               .pe48__std__lane30_strm0_ready         ( pe48__std__lane30_strm0_ready      ),      
               .std__pe48__lane30_strm0_cntl          ( std__pe48__lane30_strm0_cntl       ),      
               .std__pe48__lane30_strm0_data          ( std__pe48__lane30_strm0_data       ),      
               .std__pe48__lane30_strm0_data_valid    ( std__pe48__lane30_strm0_data_valid ),      
               .std__pe48__lane30_strm0_data_mask     ( std__pe48__lane30_strm0_data_mask  ),      

               .pe48__std__lane30_strm1_ready         ( pe48__std__lane30_strm1_ready      ),      
               .std__pe48__lane30_strm1_cntl          ( std__pe48__lane30_strm1_cntl       ),      
               .std__pe48__lane30_strm1_data          ( std__pe48__lane30_strm1_data       ),      
               .std__pe48__lane30_strm1_data_valid    ( std__pe48__lane30_strm1_data_valid ),      
               .std__pe48__lane30_strm1_data_mask     ( std__pe48__lane30_strm1_data_mask  ),      

               // PE 48, Lane 31                 
               .pe48__std__lane31_strm0_ready         ( pe48__std__lane31_strm0_ready      ),      
               .std__pe48__lane31_strm0_cntl          ( std__pe48__lane31_strm0_cntl       ),      
               .std__pe48__lane31_strm0_data          ( std__pe48__lane31_strm0_data       ),      
               .std__pe48__lane31_strm0_data_valid    ( std__pe48__lane31_strm0_data_valid ),      
               .std__pe48__lane31_strm0_data_mask     ( std__pe48__lane31_strm0_data_mask  ),      

               .pe48__std__lane31_strm1_ready         ( pe48__std__lane31_strm1_ready      ),      
               .std__pe48__lane31_strm1_cntl          ( std__pe48__lane31_strm1_cntl       ),      
               .std__pe48__lane31_strm1_data          ( std__pe48__lane31_strm1_data       ),      
               .std__pe48__lane31_strm1_data_valid    ( std__pe48__lane31_strm1_data_valid ),      
               .std__pe48__lane31_strm1_data_mask     ( std__pe48__lane31_strm1_data_mask  ),      

               // PE 49, Lane 0                 
               .pe49__std__lane0_strm0_ready         ( pe49__std__lane0_strm0_ready      ),      
               .std__pe49__lane0_strm0_cntl          ( std__pe49__lane0_strm0_cntl       ),      
               .std__pe49__lane0_strm0_data          ( std__pe49__lane0_strm0_data       ),      
               .std__pe49__lane0_strm0_data_valid    ( std__pe49__lane0_strm0_data_valid ),      
               .std__pe49__lane0_strm0_data_mask     ( std__pe49__lane0_strm0_data_mask  ),      

               .pe49__std__lane0_strm1_ready         ( pe49__std__lane0_strm1_ready      ),      
               .std__pe49__lane0_strm1_cntl          ( std__pe49__lane0_strm1_cntl       ),      
               .std__pe49__lane0_strm1_data          ( std__pe49__lane0_strm1_data       ),      
               .std__pe49__lane0_strm1_data_valid    ( std__pe49__lane0_strm1_data_valid ),      
               .std__pe49__lane0_strm1_data_mask     ( std__pe49__lane0_strm1_data_mask  ),      

               // PE 49, Lane 1                 
               .pe49__std__lane1_strm0_ready         ( pe49__std__lane1_strm0_ready      ),      
               .std__pe49__lane1_strm0_cntl          ( std__pe49__lane1_strm0_cntl       ),      
               .std__pe49__lane1_strm0_data          ( std__pe49__lane1_strm0_data       ),      
               .std__pe49__lane1_strm0_data_valid    ( std__pe49__lane1_strm0_data_valid ),      
               .std__pe49__lane1_strm0_data_mask     ( std__pe49__lane1_strm0_data_mask  ),      

               .pe49__std__lane1_strm1_ready         ( pe49__std__lane1_strm1_ready      ),      
               .std__pe49__lane1_strm1_cntl          ( std__pe49__lane1_strm1_cntl       ),      
               .std__pe49__lane1_strm1_data          ( std__pe49__lane1_strm1_data       ),      
               .std__pe49__lane1_strm1_data_valid    ( std__pe49__lane1_strm1_data_valid ),      
               .std__pe49__lane1_strm1_data_mask     ( std__pe49__lane1_strm1_data_mask  ),      

               // PE 49, Lane 2                 
               .pe49__std__lane2_strm0_ready         ( pe49__std__lane2_strm0_ready      ),      
               .std__pe49__lane2_strm0_cntl          ( std__pe49__lane2_strm0_cntl       ),      
               .std__pe49__lane2_strm0_data          ( std__pe49__lane2_strm0_data       ),      
               .std__pe49__lane2_strm0_data_valid    ( std__pe49__lane2_strm0_data_valid ),      
               .std__pe49__lane2_strm0_data_mask     ( std__pe49__lane2_strm0_data_mask  ),      

               .pe49__std__lane2_strm1_ready         ( pe49__std__lane2_strm1_ready      ),      
               .std__pe49__lane2_strm1_cntl          ( std__pe49__lane2_strm1_cntl       ),      
               .std__pe49__lane2_strm1_data          ( std__pe49__lane2_strm1_data       ),      
               .std__pe49__lane2_strm1_data_valid    ( std__pe49__lane2_strm1_data_valid ),      
               .std__pe49__lane2_strm1_data_mask     ( std__pe49__lane2_strm1_data_mask  ),      

               // PE 49, Lane 3                 
               .pe49__std__lane3_strm0_ready         ( pe49__std__lane3_strm0_ready      ),      
               .std__pe49__lane3_strm0_cntl          ( std__pe49__lane3_strm0_cntl       ),      
               .std__pe49__lane3_strm0_data          ( std__pe49__lane3_strm0_data       ),      
               .std__pe49__lane3_strm0_data_valid    ( std__pe49__lane3_strm0_data_valid ),      
               .std__pe49__lane3_strm0_data_mask     ( std__pe49__lane3_strm0_data_mask  ),      

               .pe49__std__lane3_strm1_ready         ( pe49__std__lane3_strm1_ready      ),      
               .std__pe49__lane3_strm1_cntl          ( std__pe49__lane3_strm1_cntl       ),      
               .std__pe49__lane3_strm1_data          ( std__pe49__lane3_strm1_data       ),      
               .std__pe49__lane3_strm1_data_valid    ( std__pe49__lane3_strm1_data_valid ),      
               .std__pe49__lane3_strm1_data_mask     ( std__pe49__lane3_strm1_data_mask  ),      

               // PE 49, Lane 4                 
               .pe49__std__lane4_strm0_ready         ( pe49__std__lane4_strm0_ready      ),      
               .std__pe49__lane4_strm0_cntl          ( std__pe49__lane4_strm0_cntl       ),      
               .std__pe49__lane4_strm0_data          ( std__pe49__lane4_strm0_data       ),      
               .std__pe49__lane4_strm0_data_valid    ( std__pe49__lane4_strm0_data_valid ),      
               .std__pe49__lane4_strm0_data_mask     ( std__pe49__lane4_strm0_data_mask  ),      

               .pe49__std__lane4_strm1_ready         ( pe49__std__lane4_strm1_ready      ),      
               .std__pe49__lane4_strm1_cntl          ( std__pe49__lane4_strm1_cntl       ),      
               .std__pe49__lane4_strm1_data          ( std__pe49__lane4_strm1_data       ),      
               .std__pe49__lane4_strm1_data_valid    ( std__pe49__lane4_strm1_data_valid ),      
               .std__pe49__lane4_strm1_data_mask     ( std__pe49__lane4_strm1_data_mask  ),      

               // PE 49, Lane 5                 
               .pe49__std__lane5_strm0_ready         ( pe49__std__lane5_strm0_ready      ),      
               .std__pe49__lane5_strm0_cntl          ( std__pe49__lane5_strm0_cntl       ),      
               .std__pe49__lane5_strm0_data          ( std__pe49__lane5_strm0_data       ),      
               .std__pe49__lane5_strm0_data_valid    ( std__pe49__lane5_strm0_data_valid ),      
               .std__pe49__lane5_strm0_data_mask     ( std__pe49__lane5_strm0_data_mask  ),      

               .pe49__std__lane5_strm1_ready         ( pe49__std__lane5_strm1_ready      ),      
               .std__pe49__lane5_strm1_cntl          ( std__pe49__lane5_strm1_cntl       ),      
               .std__pe49__lane5_strm1_data          ( std__pe49__lane5_strm1_data       ),      
               .std__pe49__lane5_strm1_data_valid    ( std__pe49__lane5_strm1_data_valid ),      
               .std__pe49__lane5_strm1_data_mask     ( std__pe49__lane5_strm1_data_mask  ),      

               // PE 49, Lane 6                 
               .pe49__std__lane6_strm0_ready         ( pe49__std__lane6_strm0_ready      ),      
               .std__pe49__lane6_strm0_cntl          ( std__pe49__lane6_strm0_cntl       ),      
               .std__pe49__lane6_strm0_data          ( std__pe49__lane6_strm0_data       ),      
               .std__pe49__lane6_strm0_data_valid    ( std__pe49__lane6_strm0_data_valid ),      
               .std__pe49__lane6_strm0_data_mask     ( std__pe49__lane6_strm0_data_mask  ),      

               .pe49__std__lane6_strm1_ready         ( pe49__std__lane6_strm1_ready      ),      
               .std__pe49__lane6_strm1_cntl          ( std__pe49__lane6_strm1_cntl       ),      
               .std__pe49__lane6_strm1_data          ( std__pe49__lane6_strm1_data       ),      
               .std__pe49__lane6_strm1_data_valid    ( std__pe49__lane6_strm1_data_valid ),      
               .std__pe49__lane6_strm1_data_mask     ( std__pe49__lane6_strm1_data_mask  ),      

               // PE 49, Lane 7                 
               .pe49__std__lane7_strm0_ready         ( pe49__std__lane7_strm0_ready      ),      
               .std__pe49__lane7_strm0_cntl          ( std__pe49__lane7_strm0_cntl       ),      
               .std__pe49__lane7_strm0_data          ( std__pe49__lane7_strm0_data       ),      
               .std__pe49__lane7_strm0_data_valid    ( std__pe49__lane7_strm0_data_valid ),      
               .std__pe49__lane7_strm0_data_mask     ( std__pe49__lane7_strm0_data_mask  ),      

               .pe49__std__lane7_strm1_ready         ( pe49__std__lane7_strm1_ready      ),      
               .std__pe49__lane7_strm1_cntl          ( std__pe49__lane7_strm1_cntl       ),      
               .std__pe49__lane7_strm1_data          ( std__pe49__lane7_strm1_data       ),      
               .std__pe49__lane7_strm1_data_valid    ( std__pe49__lane7_strm1_data_valid ),      
               .std__pe49__lane7_strm1_data_mask     ( std__pe49__lane7_strm1_data_mask  ),      

               // PE 49, Lane 8                 
               .pe49__std__lane8_strm0_ready         ( pe49__std__lane8_strm0_ready      ),      
               .std__pe49__lane8_strm0_cntl          ( std__pe49__lane8_strm0_cntl       ),      
               .std__pe49__lane8_strm0_data          ( std__pe49__lane8_strm0_data       ),      
               .std__pe49__lane8_strm0_data_valid    ( std__pe49__lane8_strm0_data_valid ),      
               .std__pe49__lane8_strm0_data_mask     ( std__pe49__lane8_strm0_data_mask  ),      

               .pe49__std__lane8_strm1_ready         ( pe49__std__lane8_strm1_ready      ),      
               .std__pe49__lane8_strm1_cntl          ( std__pe49__lane8_strm1_cntl       ),      
               .std__pe49__lane8_strm1_data          ( std__pe49__lane8_strm1_data       ),      
               .std__pe49__lane8_strm1_data_valid    ( std__pe49__lane8_strm1_data_valid ),      
               .std__pe49__lane8_strm1_data_mask     ( std__pe49__lane8_strm1_data_mask  ),      

               // PE 49, Lane 9                 
               .pe49__std__lane9_strm0_ready         ( pe49__std__lane9_strm0_ready      ),      
               .std__pe49__lane9_strm0_cntl          ( std__pe49__lane9_strm0_cntl       ),      
               .std__pe49__lane9_strm0_data          ( std__pe49__lane9_strm0_data       ),      
               .std__pe49__lane9_strm0_data_valid    ( std__pe49__lane9_strm0_data_valid ),      
               .std__pe49__lane9_strm0_data_mask     ( std__pe49__lane9_strm0_data_mask  ),      

               .pe49__std__lane9_strm1_ready         ( pe49__std__lane9_strm1_ready      ),      
               .std__pe49__lane9_strm1_cntl          ( std__pe49__lane9_strm1_cntl       ),      
               .std__pe49__lane9_strm1_data          ( std__pe49__lane9_strm1_data       ),      
               .std__pe49__lane9_strm1_data_valid    ( std__pe49__lane9_strm1_data_valid ),      
               .std__pe49__lane9_strm1_data_mask     ( std__pe49__lane9_strm1_data_mask  ),      

               // PE 49, Lane 10                 
               .pe49__std__lane10_strm0_ready         ( pe49__std__lane10_strm0_ready      ),      
               .std__pe49__lane10_strm0_cntl          ( std__pe49__lane10_strm0_cntl       ),      
               .std__pe49__lane10_strm0_data          ( std__pe49__lane10_strm0_data       ),      
               .std__pe49__lane10_strm0_data_valid    ( std__pe49__lane10_strm0_data_valid ),      
               .std__pe49__lane10_strm0_data_mask     ( std__pe49__lane10_strm0_data_mask  ),      

               .pe49__std__lane10_strm1_ready         ( pe49__std__lane10_strm1_ready      ),      
               .std__pe49__lane10_strm1_cntl          ( std__pe49__lane10_strm1_cntl       ),      
               .std__pe49__lane10_strm1_data          ( std__pe49__lane10_strm1_data       ),      
               .std__pe49__lane10_strm1_data_valid    ( std__pe49__lane10_strm1_data_valid ),      
               .std__pe49__lane10_strm1_data_mask     ( std__pe49__lane10_strm1_data_mask  ),      

               // PE 49, Lane 11                 
               .pe49__std__lane11_strm0_ready         ( pe49__std__lane11_strm0_ready      ),      
               .std__pe49__lane11_strm0_cntl          ( std__pe49__lane11_strm0_cntl       ),      
               .std__pe49__lane11_strm0_data          ( std__pe49__lane11_strm0_data       ),      
               .std__pe49__lane11_strm0_data_valid    ( std__pe49__lane11_strm0_data_valid ),      
               .std__pe49__lane11_strm0_data_mask     ( std__pe49__lane11_strm0_data_mask  ),      

               .pe49__std__lane11_strm1_ready         ( pe49__std__lane11_strm1_ready      ),      
               .std__pe49__lane11_strm1_cntl          ( std__pe49__lane11_strm1_cntl       ),      
               .std__pe49__lane11_strm1_data          ( std__pe49__lane11_strm1_data       ),      
               .std__pe49__lane11_strm1_data_valid    ( std__pe49__lane11_strm1_data_valid ),      
               .std__pe49__lane11_strm1_data_mask     ( std__pe49__lane11_strm1_data_mask  ),      

               // PE 49, Lane 12                 
               .pe49__std__lane12_strm0_ready         ( pe49__std__lane12_strm0_ready      ),      
               .std__pe49__lane12_strm0_cntl          ( std__pe49__lane12_strm0_cntl       ),      
               .std__pe49__lane12_strm0_data          ( std__pe49__lane12_strm0_data       ),      
               .std__pe49__lane12_strm0_data_valid    ( std__pe49__lane12_strm0_data_valid ),      
               .std__pe49__lane12_strm0_data_mask     ( std__pe49__lane12_strm0_data_mask  ),      

               .pe49__std__lane12_strm1_ready         ( pe49__std__lane12_strm1_ready      ),      
               .std__pe49__lane12_strm1_cntl          ( std__pe49__lane12_strm1_cntl       ),      
               .std__pe49__lane12_strm1_data          ( std__pe49__lane12_strm1_data       ),      
               .std__pe49__lane12_strm1_data_valid    ( std__pe49__lane12_strm1_data_valid ),      
               .std__pe49__lane12_strm1_data_mask     ( std__pe49__lane12_strm1_data_mask  ),      

               // PE 49, Lane 13                 
               .pe49__std__lane13_strm0_ready         ( pe49__std__lane13_strm0_ready      ),      
               .std__pe49__lane13_strm0_cntl          ( std__pe49__lane13_strm0_cntl       ),      
               .std__pe49__lane13_strm0_data          ( std__pe49__lane13_strm0_data       ),      
               .std__pe49__lane13_strm0_data_valid    ( std__pe49__lane13_strm0_data_valid ),      
               .std__pe49__lane13_strm0_data_mask     ( std__pe49__lane13_strm0_data_mask  ),      

               .pe49__std__lane13_strm1_ready         ( pe49__std__lane13_strm1_ready      ),      
               .std__pe49__lane13_strm1_cntl          ( std__pe49__lane13_strm1_cntl       ),      
               .std__pe49__lane13_strm1_data          ( std__pe49__lane13_strm1_data       ),      
               .std__pe49__lane13_strm1_data_valid    ( std__pe49__lane13_strm1_data_valid ),      
               .std__pe49__lane13_strm1_data_mask     ( std__pe49__lane13_strm1_data_mask  ),      

               // PE 49, Lane 14                 
               .pe49__std__lane14_strm0_ready         ( pe49__std__lane14_strm0_ready      ),      
               .std__pe49__lane14_strm0_cntl          ( std__pe49__lane14_strm0_cntl       ),      
               .std__pe49__lane14_strm0_data          ( std__pe49__lane14_strm0_data       ),      
               .std__pe49__lane14_strm0_data_valid    ( std__pe49__lane14_strm0_data_valid ),      
               .std__pe49__lane14_strm0_data_mask     ( std__pe49__lane14_strm0_data_mask  ),      

               .pe49__std__lane14_strm1_ready         ( pe49__std__lane14_strm1_ready      ),      
               .std__pe49__lane14_strm1_cntl          ( std__pe49__lane14_strm1_cntl       ),      
               .std__pe49__lane14_strm1_data          ( std__pe49__lane14_strm1_data       ),      
               .std__pe49__lane14_strm1_data_valid    ( std__pe49__lane14_strm1_data_valid ),      
               .std__pe49__lane14_strm1_data_mask     ( std__pe49__lane14_strm1_data_mask  ),      

               // PE 49, Lane 15                 
               .pe49__std__lane15_strm0_ready         ( pe49__std__lane15_strm0_ready      ),      
               .std__pe49__lane15_strm0_cntl          ( std__pe49__lane15_strm0_cntl       ),      
               .std__pe49__lane15_strm0_data          ( std__pe49__lane15_strm0_data       ),      
               .std__pe49__lane15_strm0_data_valid    ( std__pe49__lane15_strm0_data_valid ),      
               .std__pe49__lane15_strm0_data_mask     ( std__pe49__lane15_strm0_data_mask  ),      

               .pe49__std__lane15_strm1_ready         ( pe49__std__lane15_strm1_ready      ),      
               .std__pe49__lane15_strm1_cntl          ( std__pe49__lane15_strm1_cntl       ),      
               .std__pe49__lane15_strm1_data          ( std__pe49__lane15_strm1_data       ),      
               .std__pe49__lane15_strm1_data_valid    ( std__pe49__lane15_strm1_data_valid ),      
               .std__pe49__lane15_strm1_data_mask     ( std__pe49__lane15_strm1_data_mask  ),      

               // PE 49, Lane 16                 
               .pe49__std__lane16_strm0_ready         ( pe49__std__lane16_strm0_ready      ),      
               .std__pe49__lane16_strm0_cntl          ( std__pe49__lane16_strm0_cntl       ),      
               .std__pe49__lane16_strm0_data          ( std__pe49__lane16_strm0_data       ),      
               .std__pe49__lane16_strm0_data_valid    ( std__pe49__lane16_strm0_data_valid ),      
               .std__pe49__lane16_strm0_data_mask     ( std__pe49__lane16_strm0_data_mask  ),      

               .pe49__std__lane16_strm1_ready         ( pe49__std__lane16_strm1_ready      ),      
               .std__pe49__lane16_strm1_cntl          ( std__pe49__lane16_strm1_cntl       ),      
               .std__pe49__lane16_strm1_data          ( std__pe49__lane16_strm1_data       ),      
               .std__pe49__lane16_strm1_data_valid    ( std__pe49__lane16_strm1_data_valid ),      
               .std__pe49__lane16_strm1_data_mask     ( std__pe49__lane16_strm1_data_mask  ),      

               // PE 49, Lane 17                 
               .pe49__std__lane17_strm0_ready         ( pe49__std__lane17_strm0_ready      ),      
               .std__pe49__lane17_strm0_cntl          ( std__pe49__lane17_strm0_cntl       ),      
               .std__pe49__lane17_strm0_data          ( std__pe49__lane17_strm0_data       ),      
               .std__pe49__lane17_strm0_data_valid    ( std__pe49__lane17_strm0_data_valid ),      
               .std__pe49__lane17_strm0_data_mask     ( std__pe49__lane17_strm0_data_mask  ),      

               .pe49__std__lane17_strm1_ready         ( pe49__std__lane17_strm1_ready      ),      
               .std__pe49__lane17_strm1_cntl          ( std__pe49__lane17_strm1_cntl       ),      
               .std__pe49__lane17_strm1_data          ( std__pe49__lane17_strm1_data       ),      
               .std__pe49__lane17_strm1_data_valid    ( std__pe49__lane17_strm1_data_valid ),      
               .std__pe49__lane17_strm1_data_mask     ( std__pe49__lane17_strm1_data_mask  ),      

               // PE 49, Lane 18                 
               .pe49__std__lane18_strm0_ready         ( pe49__std__lane18_strm0_ready      ),      
               .std__pe49__lane18_strm0_cntl          ( std__pe49__lane18_strm0_cntl       ),      
               .std__pe49__lane18_strm0_data          ( std__pe49__lane18_strm0_data       ),      
               .std__pe49__lane18_strm0_data_valid    ( std__pe49__lane18_strm0_data_valid ),      
               .std__pe49__lane18_strm0_data_mask     ( std__pe49__lane18_strm0_data_mask  ),      

               .pe49__std__lane18_strm1_ready         ( pe49__std__lane18_strm1_ready      ),      
               .std__pe49__lane18_strm1_cntl          ( std__pe49__lane18_strm1_cntl       ),      
               .std__pe49__lane18_strm1_data          ( std__pe49__lane18_strm1_data       ),      
               .std__pe49__lane18_strm1_data_valid    ( std__pe49__lane18_strm1_data_valid ),      
               .std__pe49__lane18_strm1_data_mask     ( std__pe49__lane18_strm1_data_mask  ),      

               // PE 49, Lane 19                 
               .pe49__std__lane19_strm0_ready         ( pe49__std__lane19_strm0_ready      ),      
               .std__pe49__lane19_strm0_cntl          ( std__pe49__lane19_strm0_cntl       ),      
               .std__pe49__lane19_strm0_data          ( std__pe49__lane19_strm0_data       ),      
               .std__pe49__lane19_strm0_data_valid    ( std__pe49__lane19_strm0_data_valid ),      
               .std__pe49__lane19_strm0_data_mask     ( std__pe49__lane19_strm0_data_mask  ),      

               .pe49__std__lane19_strm1_ready         ( pe49__std__lane19_strm1_ready      ),      
               .std__pe49__lane19_strm1_cntl          ( std__pe49__lane19_strm1_cntl       ),      
               .std__pe49__lane19_strm1_data          ( std__pe49__lane19_strm1_data       ),      
               .std__pe49__lane19_strm1_data_valid    ( std__pe49__lane19_strm1_data_valid ),      
               .std__pe49__lane19_strm1_data_mask     ( std__pe49__lane19_strm1_data_mask  ),      

               // PE 49, Lane 20                 
               .pe49__std__lane20_strm0_ready         ( pe49__std__lane20_strm0_ready      ),      
               .std__pe49__lane20_strm0_cntl          ( std__pe49__lane20_strm0_cntl       ),      
               .std__pe49__lane20_strm0_data          ( std__pe49__lane20_strm0_data       ),      
               .std__pe49__lane20_strm0_data_valid    ( std__pe49__lane20_strm0_data_valid ),      
               .std__pe49__lane20_strm0_data_mask     ( std__pe49__lane20_strm0_data_mask  ),      

               .pe49__std__lane20_strm1_ready         ( pe49__std__lane20_strm1_ready      ),      
               .std__pe49__lane20_strm1_cntl          ( std__pe49__lane20_strm1_cntl       ),      
               .std__pe49__lane20_strm1_data          ( std__pe49__lane20_strm1_data       ),      
               .std__pe49__lane20_strm1_data_valid    ( std__pe49__lane20_strm1_data_valid ),      
               .std__pe49__lane20_strm1_data_mask     ( std__pe49__lane20_strm1_data_mask  ),      

               // PE 49, Lane 21                 
               .pe49__std__lane21_strm0_ready         ( pe49__std__lane21_strm0_ready      ),      
               .std__pe49__lane21_strm0_cntl          ( std__pe49__lane21_strm0_cntl       ),      
               .std__pe49__lane21_strm0_data          ( std__pe49__lane21_strm0_data       ),      
               .std__pe49__lane21_strm0_data_valid    ( std__pe49__lane21_strm0_data_valid ),      
               .std__pe49__lane21_strm0_data_mask     ( std__pe49__lane21_strm0_data_mask  ),      

               .pe49__std__lane21_strm1_ready         ( pe49__std__lane21_strm1_ready      ),      
               .std__pe49__lane21_strm1_cntl          ( std__pe49__lane21_strm1_cntl       ),      
               .std__pe49__lane21_strm1_data          ( std__pe49__lane21_strm1_data       ),      
               .std__pe49__lane21_strm1_data_valid    ( std__pe49__lane21_strm1_data_valid ),      
               .std__pe49__lane21_strm1_data_mask     ( std__pe49__lane21_strm1_data_mask  ),      

               // PE 49, Lane 22                 
               .pe49__std__lane22_strm0_ready         ( pe49__std__lane22_strm0_ready      ),      
               .std__pe49__lane22_strm0_cntl          ( std__pe49__lane22_strm0_cntl       ),      
               .std__pe49__lane22_strm0_data          ( std__pe49__lane22_strm0_data       ),      
               .std__pe49__lane22_strm0_data_valid    ( std__pe49__lane22_strm0_data_valid ),      
               .std__pe49__lane22_strm0_data_mask     ( std__pe49__lane22_strm0_data_mask  ),      

               .pe49__std__lane22_strm1_ready         ( pe49__std__lane22_strm1_ready      ),      
               .std__pe49__lane22_strm1_cntl          ( std__pe49__lane22_strm1_cntl       ),      
               .std__pe49__lane22_strm1_data          ( std__pe49__lane22_strm1_data       ),      
               .std__pe49__lane22_strm1_data_valid    ( std__pe49__lane22_strm1_data_valid ),      
               .std__pe49__lane22_strm1_data_mask     ( std__pe49__lane22_strm1_data_mask  ),      

               // PE 49, Lane 23                 
               .pe49__std__lane23_strm0_ready         ( pe49__std__lane23_strm0_ready      ),      
               .std__pe49__lane23_strm0_cntl          ( std__pe49__lane23_strm0_cntl       ),      
               .std__pe49__lane23_strm0_data          ( std__pe49__lane23_strm0_data       ),      
               .std__pe49__lane23_strm0_data_valid    ( std__pe49__lane23_strm0_data_valid ),      
               .std__pe49__lane23_strm0_data_mask     ( std__pe49__lane23_strm0_data_mask  ),      

               .pe49__std__lane23_strm1_ready         ( pe49__std__lane23_strm1_ready      ),      
               .std__pe49__lane23_strm1_cntl          ( std__pe49__lane23_strm1_cntl       ),      
               .std__pe49__lane23_strm1_data          ( std__pe49__lane23_strm1_data       ),      
               .std__pe49__lane23_strm1_data_valid    ( std__pe49__lane23_strm1_data_valid ),      
               .std__pe49__lane23_strm1_data_mask     ( std__pe49__lane23_strm1_data_mask  ),      

               // PE 49, Lane 24                 
               .pe49__std__lane24_strm0_ready         ( pe49__std__lane24_strm0_ready      ),      
               .std__pe49__lane24_strm0_cntl          ( std__pe49__lane24_strm0_cntl       ),      
               .std__pe49__lane24_strm0_data          ( std__pe49__lane24_strm0_data       ),      
               .std__pe49__lane24_strm0_data_valid    ( std__pe49__lane24_strm0_data_valid ),      
               .std__pe49__lane24_strm0_data_mask     ( std__pe49__lane24_strm0_data_mask  ),      

               .pe49__std__lane24_strm1_ready         ( pe49__std__lane24_strm1_ready      ),      
               .std__pe49__lane24_strm1_cntl          ( std__pe49__lane24_strm1_cntl       ),      
               .std__pe49__lane24_strm1_data          ( std__pe49__lane24_strm1_data       ),      
               .std__pe49__lane24_strm1_data_valid    ( std__pe49__lane24_strm1_data_valid ),      
               .std__pe49__lane24_strm1_data_mask     ( std__pe49__lane24_strm1_data_mask  ),      

               // PE 49, Lane 25                 
               .pe49__std__lane25_strm0_ready         ( pe49__std__lane25_strm0_ready      ),      
               .std__pe49__lane25_strm0_cntl          ( std__pe49__lane25_strm0_cntl       ),      
               .std__pe49__lane25_strm0_data          ( std__pe49__lane25_strm0_data       ),      
               .std__pe49__lane25_strm0_data_valid    ( std__pe49__lane25_strm0_data_valid ),      
               .std__pe49__lane25_strm0_data_mask     ( std__pe49__lane25_strm0_data_mask  ),      

               .pe49__std__lane25_strm1_ready         ( pe49__std__lane25_strm1_ready      ),      
               .std__pe49__lane25_strm1_cntl          ( std__pe49__lane25_strm1_cntl       ),      
               .std__pe49__lane25_strm1_data          ( std__pe49__lane25_strm1_data       ),      
               .std__pe49__lane25_strm1_data_valid    ( std__pe49__lane25_strm1_data_valid ),      
               .std__pe49__lane25_strm1_data_mask     ( std__pe49__lane25_strm1_data_mask  ),      

               // PE 49, Lane 26                 
               .pe49__std__lane26_strm0_ready         ( pe49__std__lane26_strm0_ready      ),      
               .std__pe49__lane26_strm0_cntl          ( std__pe49__lane26_strm0_cntl       ),      
               .std__pe49__lane26_strm0_data          ( std__pe49__lane26_strm0_data       ),      
               .std__pe49__lane26_strm0_data_valid    ( std__pe49__lane26_strm0_data_valid ),      
               .std__pe49__lane26_strm0_data_mask     ( std__pe49__lane26_strm0_data_mask  ),      

               .pe49__std__lane26_strm1_ready         ( pe49__std__lane26_strm1_ready      ),      
               .std__pe49__lane26_strm1_cntl          ( std__pe49__lane26_strm1_cntl       ),      
               .std__pe49__lane26_strm1_data          ( std__pe49__lane26_strm1_data       ),      
               .std__pe49__lane26_strm1_data_valid    ( std__pe49__lane26_strm1_data_valid ),      
               .std__pe49__lane26_strm1_data_mask     ( std__pe49__lane26_strm1_data_mask  ),      

               // PE 49, Lane 27                 
               .pe49__std__lane27_strm0_ready         ( pe49__std__lane27_strm0_ready      ),      
               .std__pe49__lane27_strm0_cntl          ( std__pe49__lane27_strm0_cntl       ),      
               .std__pe49__lane27_strm0_data          ( std__pe49__lane27_strm0_data       ),      
               .std__pe49__lane27_strm0_data_valid    ( std__pe49__lane27_strm0_data_valid ),      
               .std__pe49__lane27_strm0_data_mask     ( std__pe49__lane27_strm0_data_mask  ),      

               .pe49__std__lane27_strm1_ready         ( pe49__std__lane27_strm1_ready      ),      
               .std__pe49__lane27_strm1_cntl          ( std__pe49__lane27_strm1_cntl       ),      
               .std__pe49__lane27_strm1_data          ( std__pe49__lane27_strm1_data       ),      
               .std__pe49__lane27_strm1_data_valid    ( std__pe49__lane27_strm1_data_valid ),      
               .std__pe49__lane27_strm1_data_mask     ( std__pe49__lane27_strm1_data_mask  ),      

               // PE 49, Lane 28                 
               .pe49__std__lane28_strm0_ready         ( pe49__std__lane28_strm0_ready      ),      
               .std__pe49__lane28_strm0_cntl          ( std__pe49__lane28_strm0_cntl       ),      
               .std__pe49__lane28_strm0_data          ( std__pe49__lane28_strm0_data       ),      
               .std__pe49__lane28_strm0_data_valid    ( std__pe49__lane28_strm0_data_valid ),      
               .std__pe49__lane28_strm0_data_mask     ( std__pe49__lane28_strm0_data_mask  ),      

               .pe49__std__lane28_strm1_ready         ( pe49__std__lane28_strm1_ready      ),      
               .std__pe49__lane28_strm1_cntl          ( std__pe49__lane28_strm1_cntl       ),      
               .std__pe49__lane28_strm1_data          ( std__pe49__lane28_strm1_data       ),      
               .std__pe49__lane28_strm1_data_valid    ( std__pe49__lane28_strm1_data_valid ),      
               .std__pe49__lane28_strm1_data_mask     ( std__pe49__lane28_strm1_data_mask  ),      

               // PE 49, Lane 29                 
               .pe49__std__lane29_strm0_ready         ( pe49__std__lane29_strm0_ready      ),      
               .std__pe49__lane29_strm0_cntl          ( std__pe49__lane29_strm0_cntl       ),      
               .std__pe49__lane29_strm0_data          ( std__pe49__lane29_strm0_data       ),      
               .std__pe49__lane29_strm0_data_valid    ( std__pe49__lane29_strm0_data_valid ),      
               .std__pe49__lane29_strm0_data_mask     ( std__pe49__lane29_strm0_data_mask  ),      

               .pe49__std__lane29_strm1_ready         ( pe49__std__lane29_strm1_ready      ),      
               .std__pe49__lane29_strm1_cntl          ( std__pe49__lane29_strm1_cntl       ),      
               .std__pe49__lane29_strm1_data          ( std__pe49__lane29_strm1_data       ),      
               .std__pe49__lane29_strm1_data_valid    ( std__pe49__lane29_strm1_data_valid ),      
               .std__pe49__lane29_strm1_data_mask     ( std__pe49__lane29_strm1_data_mask  ),      

               // PE 49, Lane 30                 
               .pe49__std__lane30_strm0_ready         ( pe49__std__lane30_strm0_ready      ),      
               .std__pe49__lane30_strm0_cntl          ( std__pe49__lane30_strm0_cntl       ),      
               .std__pe49__lane30_strm0_data          ( std__pe49__lane30_strm0_data       ),      
               .std__pe49__lane30_strm0_data_valid    ( std__pe49__lane30_strm0_data_valid ),      
               .std__pe49__lane30_strm0_data_mask     ( std__pe49__lane30_strm0_data_mask  ),      

               .pe49__std__lane30_strm1_ready         ( pe49__std__lane30_strm1_ready      ),      
               .std__pe49__lane30_strm1_cntl          ( std__pe49__lane30_strm1_cntl       ),      
               .std__pe49__lane30_strm1_data          ( std__pe49__lane30_strm1_data       ),      
               .std__pe49__lane30_strm1_data_valid    ( std__pe49__lane30_strm1_data_valid ),      
               .std__pe49__lane30_strm1_data_mask     ( std__pe49__lane30_strm1_data_mask  ),      

               // PE 49, Lane 31                 
               .pe49__std__lane31_strm0_ready         ( pe49__std__lane31_strm0_ready      ),      
               .std__pe49__lane31_strm0_cntl          ( std__pe49__lane31_strm0_cntl       ),      
               .std__pe49__lane31_strm0_data          ( std__pe49__lane31_strm0_data       ),      
               .std__pe49__lane31_strm0_data_valid    ( std__pe49__lane31_strm0_data_valid ),      
               .std__pe49__lane31_strm0_data_mask     ( std__pe49__lane31_strm0_data_mask  ),      

               .pe49__std__lane31_strm1_ready         ( pe49__std__lane31_strm1_ready      ),      
               .std__pe49__lane31_strm1_cntl          ( std__pe49__lane31_strm1_cntl       ),      
               .std__pe49__lane31_strm1_data          ( std__pe49__lane31_strm1_data       ),      
               .std__pe49__lane31_strm1_data_valid    ( std__pe49__lane31_strm1_data_valid ),      
               .std__pe49__lane31_strm1_data_mask     ( std__pe49__lane31_strm1_data_mask  ),      

               // PE 50, Lane 0                 
               .pe50__std__lane0_strm0_ready         ( pe50__std__lane0_strm0_ready      ),      
               .std__pe50__lane0_strm0_cntl          ( std__pe50__lane0_strm0_cntl       ),      
               .std__pe50__lane0_strm0_data          ( std__pe50__lane0_strm0_data       ),      
               .std__pe50__lane0_strm0_data_valid    ( std__pe50__lane0_strm0_data_valid ),      
               .std__pe50__lane0_strm0_data_mask     ( std__pe50__lane0_strm0_data_mask  ),      

               .pe50__std__lane0_strm1_ready         ( pe50__std__lane0_strm1_ready      ),      
               .std__pe50__lane0_strm1_cntl          ( std__pe50__lane0_strm1_cntl       ),      
               .std__pe50__lane0_strm1_data          ( std__pe50__lane0_strm1_data       ),      
               .std__pe50__lane0_strm1_data_valid    ( std__pe50__lane0_strm1_data_valid ),      
               .std__pe50__lane0_strm1_data_mask     ( std__pe50__lane0_strm1_data_mask  ),      

               // PE 50, Lane 1                 
               .pe50__std__lane1_strm0_ready         ( pe50__std__lane1_strm0_ready      ),      
               .std__pe50__lane1_strm0_cntl          ( std__pe50__lane1_strm0_cntl       ),      
               .std__pe50__lane1_strm0_data          ( std__pe50__lane1_strm0_data       ),      
               .std__pe50__lane1_strm0_data_valid    ( std__pe50__lane1_strm0_data_valid ),      
               .std__pe50__lane1_strm0_data_mask     ( std__pe50__lane1_strm0_data_mask  ),      

               .pe50__std__lane1_strm1_ready         ( pe50__std__lane1_strm1_ready      ),      
               .std__pe50__lane1_strm1_cntl          ( std__pe50__lane1_strm1_cntl       ),      
               .std__pe50__lane1_strm1_data          ( std__pe50__lane1_strm1_data       ),      
               .std__pe50__lane1_strm1_data_valid    ( std__pe50__lane1_strm1_data_valid ),      
               .std__pe50__lane1_strm1_data_mask     ( std__pe50__lane1_strm1_data_mask  ),      

               // PE 50, Lane 2                 
               .pe50__std__lane2_strm0_ready         ( pe50__std__lane2_strm0_ready      ),      
               .std__pe50__lane2_strm0_cntl          ( std__pe50__lane2_strm0_cntl       ),      
               .std__pe50__lane2_strm0_data          ( std__pe50__lane2_strm0_data       ),      
               .std__pe50__lane2_strm0_data_valid    ( std__pe50__lane2_strm0_data_valid ),      
               .std__pe50__lane2_strm0_data_mask     ( std__pe50__lane2_strm0_data_mask  ),      

               .pe50__std__lane2_strm1_ready         ( pe50__std__lane2_strm1_ready      ),      
               .std__pe50__lane2_strm1_cntl          ( std__pe50__lane2_strm1_cntl       ),      
               .std__pe50__lane2_strm1_data          ( std__pe50__lane2_strm1_data       ),      
               .std__pe50__lane2_strm1_data_valid    ( std__pe50__lane2_strm1_data_valid ),      
               .std__pe50__lane2_strm1_data_mask     ( std__pe50__lane2_strm1_data_mask  ),      

               // PE 50, Lane 3                 
               .pe50__std__lane3_strm0_ready         ( pe50__std__lane3_strm0_ready      ),      
               .std__pe50__lane3_strm0_cntl          ( std__pe50__lane3_strm0_cntl       ),      
               .std__pe50__lane3_strm0_data          ( std__pe50__lane3_strm0_data       ),      
               .std__pe50__lane3_strm0_data_valid    ( std__pe50__lane3_strm0_data_valid ),      
               .std__pe50__lane3_strm0_data_mask     ( std__pe50__lane3_strm0_data_mask  ),      

               .pe50__std__lane3_strm1_ready         ( pe50__std__lane3_strm1_ready      ),      
               .std__pe50__lane3_strm1_cntl          ( std__pe50__lane3_strm1_cntl       ),      
               .std__pe50__lane3_strm1_data          ( std__pe50__lane3_strm1_data       ),      
               .std__pe50__lane3_strm1_data_valid    ( std__pe50__lane3_strm1_data_valid ),      
               .std__pe50__lane3_strm1_data_mask     ( std__pe50__lane3_strm1_data_mask  ),      

               // PE 50, Lane 4                 
               .pe50__std__lane4_strm0_ready         ( pe50__std__lane4_strm0_ready      ),      
               .std__pe50__lane4_strm0_cntl          ( std__pe50__lane4_strm0_cntl       ),      
               .std__pe50__lane4_strm0_data          ( std__pe50__lane4_strm0_data       ),      
               .std__pe50__lane4_strm0_data_valid    ( std__pe50__lane4_strm0_data_valid ),      
               .std__pe50__lane4_strm0_data_mask     ( std__pe50__lane4_strm0_data_mask  ),      

               .pe50__std__lane4_strm1_ready         ( pe50__std__lane4_strm1_ready      ),      
               .std__pe50__lane4_strm1_cntl          ( std__pe50__lane4_strm1_cntl       ),      
               .std__pe50__lane4_strm1_data          ( std__pe50__lane4_strm1_data       ),      
               .std__pe50__lane4_strm1_data_valid    ( std__pe50__lane4_strm1_data_valid ),      
               .std__pe50__lane4_strm1_data_mask     ( std__pe50__lane4_strm1_data_mask  ),      

               // PE 50, Lane 5                 
               .pe50__std__lane5_strm0_ready         ( pe50__std__lane5_strm0_ready      ),      
               .std__pe50__lane5_strm0_cntl          ( std__pe50__lane5_strm0_cntl       ),      
               .std__pe50__lane5_strm0_data          ( std__pe50__lane5_strm0_data       ),      
               .std__pe50__lane5_strm0_data_valid    ( std__pe50__lane5_strm0_data_valid ),      
               .std__pe50__lane5_strm0_data_mask     ( std__pe50__lane5_strm0_data_mask  ),      

               .pe50__std__lane5_strm1_ready         ( pe50__std__lane5_strm1_ready      ),      
               .std__pe50__lane5_strm1_cntl          ( std__pe50__lane5_strm1_cntl       ),      
               .std__pe50__lane5_strm1_data          ( std__pe50__lane5_strm1_data       ),      
               .std__pe50__lane5_strm1_data_valid    ( std__pe50__lane5_strm1_data_valid ),      
               .std__pe50__lane5_strm1_data_mask     ( std__pe50__lane5_strm1_data_mask  ),      

               // PE 50, Lane 6                 
               .pe50__std__lane6_strm0_ready         ( pe50__std__lane6_strm0_ready      ),      
               .std__pe50__lane6_strm0_cntl          ( std__pe50__lane6_strm0_cntl       ),      
               .std__pe50__lane6_strm0_data          ( std__pe50__lane6_strm0_data       ),      
               .std__pe50__lane6_strm0_data_valid    ( std__pe50__lane6_strm0_data_valid ),      
               .std__pe50__lane6_strm0_data_mask     ( std__pe50__lane6_strm0_data_mask  ),      

               .pe50__std__lane6_strm1_ready         ( pe50__std__lane6_strm1_ready      ),      
               .std__pe50__lane6_strm1_cntl          ( std__pe50__lane6_strm1_cntl       ),      
               .std__pe50__lane6_strm1_data          ( std__pe50__lane6_strm1_data       ),      
               .std__pe50__lane6_strm1_data_valid    ( std__pe50__lane6_strm1_data_valid ),      
               .std__pe50__lane6_strm1_data_mask     ( std__pe50__lane6_strm1_data_mask  ),      

               // PE 50, Lane 7                 
               .pe50__std__lane7_strm0_ready         ( pe50__std__lane7_strm0_ready      ),      
               .std__pe50__lane7_strm0_cntl          ( std__pe50__lane7_strm0_cntl       ),      
               .std__pe50__lane7_strm0_data          ( std__pe50__lane7_strm0_data       ),      
               .std__pe50__lane7_strm0_data_valid    ( std__pe50__lane7_strm0_data_valid ),      
               .std__pe50__lane7_strm0_data_mask     ( std__pe50__lane7_strm0_data_mask  ),      

               .pe50__std__lane7_strm1_ready         ( pe50__std__lane7_strm1_ready      ),      
               .std__pe50__lane7_strm1_cntl          ( std__pe50__lane7_strm1_cntl       ),      
               .std__pe50__lane7_strm1_data          ( std__pe50__lane7_strm1_data       ),      
               .std__pe50__lane7_strm1_data_valid    ( std__pe50__lane7_strm1_data_valid ),      
               .std__pe50__lane7_strm1_data_mask     ( std__pe50__lane7_strm1_data_mask  ),      

               // PE 50, Lane 8                 
               .pe50__std__lane8_strm0_ready         ( pe50__std__lane8_strm0_ready      ),      
               .std__pe50__lane8_strm0_cntl          ( std__pe50__lane8_strm0_cntl       ),      
               .std__pe50__lane8_strm0_data          ( std__pe50__lane8_strm0_data       ),      
               .std__pe50__lane8_strm0_data_valid    ( std__pe50__lane8_strm0_data_valid ),      
               .std__pe50__lane8_strm0_data_mask     ( std__pe50__lane8_strm0_data_mask  ),      

               .pe50__std__lane8_strm1_ready         ( pe50__std__lane8_strm1_ready      ),      
               .std__pe50__lane8_strm1_cntl          ( std__pe50__lane8_strm1_cntl       ),      
               .std__pe50__lane8_strm1_data          ( std__pe50__lane8_strm1_data       ),      
               .std__pe50__lane8_strm1_data_valid    ( std__pe50__lane8_strm1_data_valid ),      
               .std__pe50__lane8_strm1_data_mask     ( std__pe50__lane8_strm1_data_mask  ),      

               // PE 50, Lane 9                 
               .pe50__std__lane9_strm0_ready         ( pe50__std__lane9_strm0_ready      ),      
               .std__pe50__lane9_strm0_cntl          ( std__pe50__lane9_strm0_cntl       ),      
               .std__pe50__lane9_strm0_data          ( std__pe50__lane9_strm0_data       ),      
               .std__pe50__lane9_strm0_data_valid    ( std__pe50__lane9_strm0_data_valid ),      
               .std__pe50__lane9_strm0_data_mask     ( std__pe50__lane9_strm0_data_mask  ),      

               .pe50__std__lane9_strm1_ready         ( pe50__std__lane9_strm1_ready      ),      
               .std__pe50__lane9_strm1_cntl          ( std__pe50__lane9_strm1_cntl       ),      
               .std__pe50__lane9_strm1_data          ( std__pe50__lane9_strm1_data       ),      
               .std__pe50__lane9_strm1_data_valid    ( std__pe50__lane9_strm1_data_valid ),      
               .std__pe50__lane9_strm1_data_mask     ( std__pe50__lane9_strm1_data_mask  ),      

               // PE 50, Lane 10                 
               .pe50__std__lane10_strm0_ready         ( pe50__std__lane10_strm0_ready      ),      
               .std__pe50__lane10_strm0_cntl          ( std__pe50__lane10_strm0_cntl       ),      
               .std__pe50__lane10_strm0_data          ( std__pe50__lane10_strm0_data       ),      
               .std__pe50__lane10_strm0_data_valid    ( std__pe50__lane10_strm0_data_valid ),      
               .std__pe50__lane10_strm0_data_mask     ( std__pe50__lane10_strm0_data_mask  ),      

               .pe50__std__lane10_strm1_ready         ( pe50__std__lane10_strm1_ready      ),      
               .std__pe50__lane10_strm1_cntl          ( std__pe50__lane10_strm1_cntl       ),      
               .std__pe50__lane10_strm1_data          ( std__pe50__lane10_strm1_data       ),      
               .std__pe50__lane10_strm1_data_valid    ( std__pe50__lane10_strm1_data_valid ),      
               .std__pe50__lane10_strm1_data_mask     ( std__pe50__lane10_strm1_data_mask  ),      

               // PE 50, Lane 11                 
               .pe50__std__lane11_strm0_ready         ( pe50__std__lane11_strm0_ready      ),      
               .std__pe50__lane11_strm0_cntl          ( std__pe50__lane11_strm0_cntl       ),      
               .std__pe50__lane11_strm0_data          ( std__pe50__lane11_strm0_data       ),      
               .std__pe50__lane11_strm0_data_valid    ( std__pe50__lane11_strm0_data_valid ),      
               .std__pe50__lane11_strm0_data_mask     ( std__pe50__lane11_strm0_data_mask  ),      

               .pe50__std__lane11_strm1_ready         ( pe50__std__lane11_strm1_ready      ),      
               .std__pe50__lane11_strm1_cntl          ( std__pe50__lane11_strm1_cntl       ),      
               .std__pe50__lane11_strm1_data          ( std__pe50__lane11_strm1_data       ),      
               .std__pe50__lane11_strm1_data_valid    ( std__pe50__lane11_strm1_data_valid ),      
               .std__pe50__lane11_strm1_data_mask     ( std__pe50__lane11_strm1_data_mask  ),      

               // PE 50, Lane 12                 
               .pe50__std__lane12_strm0_ready         ( pe50__std__lane12_strm0_ready      ),      
               .std__pe50__lane12_strm0_cntl          ( std__pe50__lane12_strm0_cntl       ),      
               .std__pe50__lane12_strm0_data          ( std__pe50__lane12_strm0_data       ),      
               .std__pe50__lane12_strm0_data_valid    ( std__pe50__lane12_strm0_data_valid ),      
               .std__pe50__lane12_strm0_data_mask     ( std__pe50__lane12_strm0_data_mask  ),      

               .pe50__std__lane12_strm1_ready         ( pe50__std__lane12_strm1_ready      ),      
               .std__pe50__lane12_strm1_cntl          ( std__pe50__lane12_strm1_cntl       ),      
               .std__pe50__lane12_strm1_data          ( std__pe50__lane12_strm1_data       ),      
               .std__pe50__lane12_strm1_data_valid    ( std__pe50__lane12_strm1_data_valid ),      
               .std__pe50__lane12_strm1_data_mask     ( std__pe50__lane12_strm1_data_mask  ),      

               // PE 50, Lane 13                 
               .pe50__std__lane13_strm0_ready         ( pe50__std__lane13_strm0_ready      ),      
               .std__pe50__lane13_strm0_cntl          ( std__pe50__lane13_strm0_cntl       ),      
               .std__pe50__lane13_strm0_data          ( std__pe50__lane13_strm0_data       ),      
               .std__pe50__lane13_strm0_data_valid    ( std__pe50__lane13_strm0_data_valid ),      
               .std__pe50__lane13_strm0_data_mask     ( std__pe50__lane13_strm0_data_mask  ),      

               .pe50__std__lane13_strm1_ready         ( pe50__std__lane13_strm1_ready      ),      
               .std__pe50__lane13_strm1_cntl          ( std__pe50__lane13_strm1_cntl       ),      
               .std__pe50__lane13_strm1_data          ( std__pe50__lane13_strm1_data       ),      
               .std__pe50__lane13_strm1_data_valid    ( std__pe50__lane13_strm1_data_valid ),      
               .std__pe50__lane13_strm1_data_mask     ( std__pe50__lane13_strm1_data_mask  ),      

               // PE 50, Lane 14                 
               .pe50__std__lane14_strm0_ready         ( pe50__std__lane14_strm0_ready      ),      
               .std__pe50__lane14_strm0_cntl          ( std__pe50__lane14_strm0_cntl       ),      
               .std__pe50__lane14_strm0_data          ( std__pe50__lane14_strm0_data       ),      
               .std__pe50__lane14_strm0_data_valid    ( std__pe50__lane14_strm0_data_valid ),      
               .std__pe50__lane14_strm0_data_mask     ( std__pe50__lane14_strm0_data_mask  ),      

               .pe50__std__lane14_strm1_ready         ( pe50__std__lane14_strm1_ready      ),      
               .std__pe50__lane14_strm1_cntl          ( std__pe50__lane14_strm1_cntl       ),      
               .std__pe50__lane14_strm1_data          ( std__pe50__lane14_strm1_data       ),      
               .std__pe50__lane14_strm1_data_valid    ( std__pe50__lane14_strm1_data_valid ),      
               .std__pe50__lane14_strm1_data_mask     ( std__pe50__lane14_strm1_data_mask  ),      

               // PE 50, Lane 15                 
               .pe50__std__lane15_strm0_ready         ( pe50__std__lane15_strm0_ready      ),      
               .std__pe50__lane15_strm0_cntl          ( std__pe50__lane15_strm0_cntl       ),      
               .std__pe50__lane15_strm0_data          ( std__pe50__lane15_strm0_data       ),      
               .std__pe50__lane15_strm0_data_valid    ( std__pe50__lane15_strm0_data_valid ),      
               .std__pe50__lane15_strm0_data_mask     ( std__pe50__lane15_strm0_data_mask  ),      

               .pe50__std__lane15_strm1_ready         ( pe50__std__lane15_strm1_ready      ),      
               .std__pe50__lane15_strm1_cntl          ( std__pe50__lane15_strm1_cntl       ),      
               .std__pe50__lane15_strm1_data          ( std__pe50__lane15_strm1_data       ),      
               .std__pe50__lane15_strm1_data_valid    ( std__pe50__lane15_strm1_data_valid ),      
               .std__pe50__lane15_strm1_data_mask     ( std__pe50__lane15_strm1_data_mask  ),      

               // PE 50, Lane 16                 
               .pe50__std__lane16_strm0_ready         ( pe50__std__lane16_strm0_ready      ),      
               .std__pe50__lane16_strm0_cntl          ( std__pe50__lane16_strm0_cntl       ),      
               .std__pe50__lane16_strm0_data          ( std__pe50__lane16_strm0_data       ),      
               .std__pe50__lane16_strm0_data_valid    ( std__pe50__lane16_strm0_data_valid ),      
               .std__pe50__lane16_strm0_data_mask     ( std__pe50__lane16_strm0_data_mask  ),      

               .pe50__std__lane16_strm1_ready         ( pe50__std__lane16_strm1_ready      ),      
               .std__pe50__lane16_strm1_cntl          ( std__pe50__lane16_strm1_cntl       ),      
               .std__pe50__lane16_strm1_data          ( std__pe50__lane16_strm1_data       ),      
               .std__pe50__lane16_strm1_data_valid    ( std__pe50__lane16_strm1_data_valid ),      
               .std__pe50__lane16_strm1_data_mask     ( std__pe50__lane16_strm1_data_mask  ),      

               // PE 50, Lane 17                 
               .pe50__std__lane17_strm0_ready         ( pe50__std__lane17_strm0_ready      ),      
               .std__pe50__lane17_strm0_cntl          ( std__pe50__lane17_strm0_cntl       ),      
               .std__pe50__lane17_strm0_data          ( std__pe50__lane17_strm0_data       ),      
               .std__pe50__lane17_strm0_data_valid    ( std__pe50__lane17_strm0_data_valid ),      
               .std__pe50__lane17_strm0_data_mask     ( std__pe50__lane17_strm0_data_mask  ),      

               .pe50__std__lane17_strm1_ready         ( pe50__std__lane17_strm1_ready      ),      
               .std__pe50__lane17_strm1_cntl          ( std__pe50__lane17_strm1_cntl       ),      
               .std__pe50__lane17_strm1_data          ( std__pe50__lane17_strm1_data       ),      
               .std__pe50__lane17_strm1_data_valid    ( std__pe50__lane17_strm1_data_valid ),      
               .std__pe50__lane17_strm1_data_mask     ( std__pe50__lane17_strm1_data_mask  ),      

               // PE 50, Lane 18                 
               .pe50__std__lane18_strm0_ready         ( pe50__std__lane18_strm0_ready      ),      
               .std__pe50__lane18_strm0_cntl          ( std__pe50__lane18_strm0_cntl       ),      
               .std__pe50__lane18_strm0_data          ( std__pe50__lane18_strm0_data       ),      
               .std__pe50__lane18_strm0_data_valid    ( std__pe50__lane18_strm0_data_valid ),      
               .std__pe50__lane18_strm0_data_mask     ( std__pe50__lane18_strm0_data_mask  ),      

               .pe50__std__lane18_strm1_ready         ( pe50__std__lane18_strm1_ready      ),      
               .std__pe50__lane18_strm1_cntl          ( std__pe50__lane18_strm1_cntl       ),      
               .std__pe50__lane18_strm1_data          ( std__pe50__lane18_strm1_data       ),      
               .std__pe50__lane18_strm1_data_valid    ( std__pe50__lane18_strm1_data_valid ),      
               .std__pe50__lane18_strm1_data_mask     ( std__pe50__lane18_strm1_data_mask  ),      

               // PE 50, Lane 19                 
               .pe50__std__lane19_strm0_ready         ( pe50__std__lane19_strm0_ready      ),      
               .std__pe50__lane19_strm0_cntl          ( std__pe50__lane19_strm0_cntl       ),      
               .std__pe50__lane19_strm0_data          ( std__pe50__lane19_strm0_data       ),      
               .std__pe50__lane19_strm0_data_valid    ( std__pe50__lane19_strm0_data_valid ),      
               .std__pe50__lane19_strm0_data_mask     ( std__pe50__lane19_strm0_data_mask  ),      

               .pe50__std__lane19_strm1_ready         ( pe50__std__lane19_strm1_ready      ),      
               .std__pe50__lane19_strm1_cntl          ( std__pe50__lane19_strm1_cntl       ),      
               .std__pe50__lane19_strm1_data          ( std__pe50__lane19_strm1_data       ),      
               .std__pe50__lane19_strm1_data_valid    ( std__pe50__lane19_strm1_data_valid ),      
               .std__pe50__lane19_strm1_data_mask     ( std__pe50__lane19_strm1_data_mask  ),      

               // PE 50, Lane 20                 
               .pe50__std__lane20_strm0_ready         ( pe50__std__lane20_strm0_ready      ),      
               .std__pe50__lane20_strm0_cntl          ( std__pe50__lane20_strm0_cntl       ),      
               .std__pe50__lane20_strm0_data          ( std__pe50__lane20_strm0_data       ),      
               .std__pe50__lane20_strm0_data_valid    ( std__pe50__lane20_strm0_data_valid ),      
               .std__pe50__lane20_strm0_data_mask     ( std__pe50__lane20_strm0_data_mask  ),      

               .pe50__std__lane20_strm1_ready         ( pe50__std__lane20_strm1_ready      ),      
               .std__pe50__lane20_strm1_cntl          ( std__pe50__lane20_strm1_cntl       ),      
               .std__pe50__lane20_strm1_data          ( std__pe50__lane20_strm1_data       ),      
               .std__pe50__lane20_strm1_data_valid    ( std__pe50__lane20_strm1_data_valid ),      
               .std__pe50__lane20_strm1_data_mask     ( std__pe50__lane20_strm1_data_mask  ),      

               // PE 50, Lane 21                 
               .pe50__std__lane21_strm0_ready         ( pe50__std__lane21_strm0_ready      ),      
               .std__pe50__lane21_strm0_cntl          ( std__pe50__lane21_strm0_cntl       ),      
               .std__pe50__lane21_strm0_data          ( std__pe50__lane21_strm0_data       ),      
               .std__pe50__lane21_strm0_data_valid    ( std__pe50__lane21_strm0_data_valid ),      
               .std__pe50__lane21_strm0_data_mask     ( std__pe50__lane21_strm0_data_mask  ),      

               .pe50__std__lane21_strm1_ready         ( pe50__std__lane21_strm1_ready      ),      
               .std__pe50__lane21_strm1_cntl          ( std__pe50__lane21_strm1_cntl       ),      
               .std__pe50__lane21_strm1_data          ( std__pe50__lane21_strm1_data       ),      
               .std__pe50__lane21_strm1_data_valid    ( std__pe50__lane21_strm1_data_valid ),      
               .std__pe50__lane21_strm1_data_mask     ( std__pe50__lane21_strm1_data_mask  ),      

               // PE 50, Lane 22                 
               .pe50__std__lane22_strm0_ready         ( pe50__std__lane22_strm0_ready      ),      
               .std__pe50__lane22_strm0_cntl          ( std__pe50__lane22_strm0_cntl       ),      
               .std__pe50__lane22_strm0_data          ( std__pe50__lane22_strm0_data       ),      
               .std__pe50__lane22_strm0_data_valid    ( std__pe50__lane22_strm0_data_valid ),      
               .std__pe50__lane22_strm0_data_mask     ( std__pe50__lane22_strm0_data_mask  ),      

               .pe50__std__lane22_strm1_ready         ( pe50__std__lane22_strm1_ready      ),      
               .std__pe50__lane22_strm1_cntl          ( std__pe50__lane22_strm1_cntl       ),      
               .std__pe50__lane22_strm1_data          ( std__pe50__lane22_strm1_data       ),      
               .std__pe50__lane22_strm1_data_valid    ( std__pe50__lane22_strm1_data_valid ),      
               .std__pe50__lane22_strm1_data_mask     ( std__pe50__lane22_strm1_data_mask  ),      

               // PE 50, Lane 23                 
               .pe50__std__lane23_strm0_ready         ( pe50__std__lane23_strm0_ready      ),      
               .std__pe50__lane23_strm0_cntl          ( std__pe50__lane23_strm0_cntl       ),      
               .std__pe50__lane23_strm0_data          ( std__pe50__lane23_strm0_data       ),      
               .std__pe50__lane23_strm0_data_valid    ( std__pe50__lane23_strm0_data_valid ),      
               .std__pe50__lane23_strm0_data_mask     ( std__pe50__lane23_strm0_data_mask  ),      

               .pe50__std__lane23_strm1_ready         ( pe50__std__lane23_strm1_ready      ),      
               .std__pe50__lane23_strm1_cntl          ( std__pe50__lane23_strm1_cntl       ),      
               .std__pe50__lane23_strm1_data          ( std__pe50__lane23_strm1_data       ),      
               .std__pe50__lane23_strm1_data_valid    ( std__pe50__lane23_strm1_data_valid ),      
               .std__pe50__lane23_strm1_data_mask     ( std__pe50__lane23_strm1_data_mask  ),      

               // PE 50, Lane 24                 
               .pe50__std__lane24_strm0_ready         ( pe50__std__lane24_strm0_ready      ),      
               .std__pe50__lane24_strm0_cntl          ( std__pe50__lane24_strm0_cntl       ),      
               .std__pe50__lane24_strm0_data          ( std__pe50__lane24_strm0_data       ),      
               .std__pe50__lane24_strm0_data_valid    ( std__pe50__lane24_strm0_data_valid ),      
               .std__pe50__lane24_strm0_data_mask     ( std__pe50__lane24_strm0_data_mask  ),      

               .pe50__std__lane24_strm1_ready         ( pe50__std__lane24_strm1_ready      ),      
               .std__pe50__lane24_strm1_cntl          ( std__pe50__lane24_strm1_cntl       ),      
               .std__pe50__lane24_strm1_data          ( std__pe50__lane24_strm1_data       ),      
               .std__pe50__lane24_strm1_data_valid    ( std__pe50__lane24_strm1_data_valid ),      
               .std__pe50__lane24_strm1_data_mask     ( std__pe50__lane24_strm1_data_mask  ),      

               // PE 50, Lane 25                 
               .pe50__std__lane25_strm0_ready         ( pe50__std__lane25_strm0_ready      ),      
               .std__pe50__lane25_strm0_cntl          ( std__pe50__lane25_strm0_cntl       ),      
               .std__pe50__lane25_strm0_data          ( std__pe50__lane25_strm0_data       ),      
               .std__pe50__lane25_strm0_data_valid    ( std__pe50__lane25_strm0_data_valid ),      
               .std__pe50__lane25_strm0_data_mask     ( std__pe50__lane25_strm0_data_mask  ),      

               .pe50__std__lane25_strm1_ready         ( pe50__std__lane25_strm1_ready      ),      
               .std__pe50__lane25_strm1_cntl          ( std__pe50__lane25_strm1_cntl       ),      
               .std__pe50__lane25_strm1_data          ( std__pe50__lane25_strm1_data       ),      
               .std__pe50__lane25_strm1_data_valid    ( std__pe50__lane25_strm1_data_valid ),      
               .std__pe50__lane25_strm1_data_mask     ( std__pe50__lane25_strm1_data_mask  ),      

               // PE 50, Lane 26                 
               .pe50__std__lane26_strm0_ready         ( pe50__std__lane26_strm0_ready      ),      
               .std__pe50__lane26_strm0_cntl          ( std__pe50__lane26_strm0_cntl       ),      
               .std__pe50__lane26_strm0_data          ( std__pe50__lane26_strm0_data       ),      
               .std__pe50__lane26_strm0_data_valid    ( std__pe50__lane26_strm0_data_valid ),      
               .std__pe50__lane26_strm0_data_mask     ( std__pe50__lane26_strm0_data_mask  ),      

               .pe50__std__lane26_strm1_ready         ( pe50__std__lane26_strm1_ready      ),      
               .std__pe50__lane26_strm1_cntl          ( std__pe50__lane26_strm1_cntl       ),      
               .std__pe50__lane26_strm1_data          ( std__pe50__lane26_strm1_data       ),      
               .std__pe50__lane26_strm1_data_valid    ( std__pe50__lane26_strm1_data_valid ),      
               .std__pe50__lane26_strm1_data_mask     ( std__pe50__lane26_strm1_data_mask  ),      

               // PE 50, Lane 27                 
               .pe50__std__lane27_strm0_ready         ( pe50__std__lane27_strm0_ready      ),      
               .std__pe50__lane27_strm0_cntl          ( std__pe50__lane27_strm0_cntl       ),      
               .std__pe50__lane27_strm0_data          ( std__pe50__lane27_strm0_data       ),      
               .std__pe50__lane27_strm0_data_valid    ( std__pe50__lane27_strm0_data_valid ),      
               .std__pe50__lane27_strm0_data_mask     ( std__pe50__lane27_strm0_data_mask  ),      

               .pe50__std__lane27_strm1_ready         ( pe50__std__lane27_strm1_ready      ),      
               .std__pe50__lane27_strm1_cntl          ( std__pe50__lane27_strm1_cntl       ),      
               .std__pe50__lane27_strm1_data          ( std__pe50__lane27_strm1_data       ),      
               .std__pe50__lane27_strm1_data_valid    ( std__pe50__lane27_strm1_data_valid ),      
               .std__pe50__lane27_strm1_data_mask     ( std__pe50__lane27_strm1_data_mask  ),      

               // PE 50, Lane 28                 
               .pe50__std__lane28_strm0_ready         ( pe50__std__lane28_strm0_ready      ),      
               .std__pe50__lane28_strm0_cntl          ( std__pe50__lane28_strm0_cntl       ),      
               .std__pe50__lane28_strm0_data          ( std__pe50__lane28_strm0_data       ),      
               .std__pe50__lane28_strm0_data_valid    ( std__pe50__lane28_strm0_data_valid ),      
               .std__pe50__lane28_strm0_data_mask     ( std__pe50__lane28_strm0_data_mask  ),      

               .pe50__std__lane28_strm1_ready         ( pe50__std__lane28_strm1_ready      ),      
               .std__pe50__lane28_strm1_cntl          ( std__pe50__lane28_strm1_cntl       ),      
               .std__pe50__lane28_strm1_data          ( std__pe50__lane28_strm1_data       ),      
               .std__pe50__lane28_strm1_data_valid    ( std__pe50__lane28_strm1_data_valid ),      
               .std__pe50__lane28_strm1_data_mask     ( std__pe50__lane28_strm1_data_mask  ),      

               // PE 50, Lane 29                 
               .pe50__std__lane29_strm0_ready         ( pe50__std__lane29_strm0_ready      ),      
               .std__pe50__lane29_strm0_cntl          ( std__pe50__lane29_strm0_cntl       ),      
               .std__pe50__lane29_strm0_data          ( std__pe50__lane29_strm0_data       ),      
               .std__pe50__lane29_strm0_data_valid    ( std__pe50__lane29_strm0_data_valid ),      
               .std__pe50__lane29_strm0_data_mask     ( std__pe50__lane29_strm0_data_mask  ),      

               .pe50__std__lane29_strm1_ready         ( pe50__std__lane29_strm1_ready      ),      
               .std__pe50__lane29_strm1_cntl          ( std__pe50__lane29_strm1_cntl       ),      
               .std__pe50__lane29_strm1_data          ( std__pe50__lane29_strm1_data       ),      
               .std__pe50__lane29_strm1_data_valid    ( std__pe50__lane29_strm1_data_valid ),      
               .std__pe50__lane29_strm1_data_mask     ( std__pe50__lane29_strm1_data_mask  ),      

               // PE 50, Lane 30                 
               .pe50__std__lane30_strm0_ready         ( pe50__std__lane30_strm0_ready      ),      
               .std__pe50__lane30_strm0_cntl          ( std__pe50__lane30_strm0_cntl       ),      
               .std__pe50__lane30_strm0_data          ( std__pe50__lane30_strm0_data       ),      
               .std__pe50__lane30_strm0_data_valid    ( std__pe50__lane30_strm0_data_valid ),      
               .std__pe50__lane30_strm0_data_mask     ( std__pe50__lane30_strm0_data_mask  ),      

               .pe50__std__lane30_strm1_ready         ( pe50__std__lane30_strm1_ready      ),      
               .std__pe50__lane30_strm1_cntl          ( std__pe50__lane30_strm1_cntl       ),      
               .std__pe50__lane30_strm1_data          ( std__pe50__lane30_strm1_data       ),      
               .std__pe50__lane30_strm1_data_valid    ( std__pe50__lane30_strm1_data_valid ),      
               .std__pe50__lane30_strm1_data_mask     ( std__pe50__lane30_strm1_data_mask  ),      

               // PE 50, Lane 31                 
               .pe50__std__lane31_strm0_ready         ( pe50__std__lane31_strm0_ready      ),      
               .std__pe50__lane31_strm0_cntl          ( std__pe50__lane31_strm0_cntl       ),      
               .std__pe50__lane31_strm0_data          ( std__pe50__lane31_strm0_data       ),      
               .std__pe50__lane31_strm0_data_valid    ( std__pe50__lane31_strm0_data_valid ),      
               .std__pe50__lane31_strm0_data_mask     ( std__pe50__lane31_strm0_data_mask  ),      

               .pe50__std__lane31_strm1_ready         ( pe50__std__lane31_strm1_ready      ),      
               .std__pe50__lane31_strm1_cntl          ( std__pe50__lane31_strm1_cntl       ),      
               .std__pe50__lane31_strm1_data          ( std__pe50__lane31_strm1_data       ),      
               .std__pe50__lane31_strm1_data_valid    ( std__pe50__lane31_strm1_data_valid ),      
               .std__pe50__lane31_strm1_data_mask     ( std__pe50__lane31_strm1_data_mask  ),      

               // PE 51, Lane 0                 
               .pe51__std__lane0_strm0_ready         ( pe51__std__lane0_strm0_ready      ),      
               .std__pe51__lane0_strm0_cntl          ( std__pe51__lane0_strm0_cntl       ),      
               .std__pe51__lane0_strm0_data          ( std__pe51__lane0_strm0_data       ),      
               .std__pe51__lane0_strm0_data_valid    ( std__pe51__lane0_strm0_data_valid ),      
               .std__pe51__lane0_strm0_data_mask     ( std__pe51__lane0_strm0_data_mask  ),      

               .pe51__std__lane0_strm1_ready         ( pe51__std__lane0_strm1_ready      ),      
               .std__pe51__lane0_strm1_cntl          ( std__pe51__lane0_strm1_cntl       ),      
               .std__pe51__lane0_strm1_data          ( std__pe51__lane0_strm1_data       ),      
               .std__pe51__lane0_strm1_data_valid    ( std__pe51__lane0_strm1_data_valid ),      
               .std__pe51__lane0_strm1_data_mask     ( std__pe51__lane0_strm1_data_mask  ),      

               // PE 51, Lane 1                 
               .pe51__std__lane1_strm0_ready         ( pe51__std__lane1_strm0_ready      ),      
               .std__pe51__lane1_strm0_cntl          ( std__pe51__lane1_strm0_cntl       ),      
               .std__pe51__lane1_strm0_data          ( std__pe51__lane1_strm0_data       ),      
               .std__pe51__lane1_strm0_data_valid    ( std__pe51__lane1_strm0_data_valid ),      
               .std__pe51__lane1_strm0_data_mask     ( std__pe51__lane1_strm0_data_mask  ),      

               .pe51__std__lane1_strm1_ready         ( pe51__std__lane1_strm1_ready      ),      
               .std__pe51__lane1_strm1_cntl          ( std__pe51__lane1_strm1_cntl       ),      
               .std__pe51__lane1_strm1_data          ( std__pe51__lane1_strm1_data       ),      
               .std__pe51__lane1_strm1_data_valid    ( std__pe51__lane1_strm1_data_valid ),      
               .std__pe51__lane1_strm1_data_mask     ( std__pe51__lane1_strm1_data_mask  ),      

               // PE 51, Lane 2                 
               .pe51__std__lane2_strm0_ready         ( pe51__std__lane2_strm0_ready      ),      
               .std__pe51__lane2_strm0_cntl          ( std__pe51__lane2_strm0_cntl       ),      
               .std__pe51__lane2_strm0_data          ( std__pe51__lane2_strm0_data       ),      
               .std__pe51__lane2_strm0_data_valid    ( std__pe51__lane2_strm0_data_valid ),      
               .std__pe51__lane2_strm0_data_mask     ( std__pe51__lane2_strm0_data_mask  ),      

               .pe51__std__lane2_strm1_ready         ( pe51__std__lane2_strm1_ready      ),      
               .std__pe51__lane2_strm1_cntl          ( std__pe51__lane2_strm1_cntl       ),      
               .std__pe51__lane2_strm1_data          ( std__pe51__lane2_strm1_data       ),      
               .std__pe51__lane2_strm1_data_valid    ( std__pe51__lane2_strm1_data_valid ),      
               .std__pe51__lane2_strm1_data_mask     ( std__pe51__lane2_strm1_data_mask  ),      

               // PE 51, Lane 3                 
               .pe51__std__lane3_strm0_ready         ( pe51__std__lane3_strm0_ready      ),      
               .std__pe51__lane3_strm0_cntl          ( std__pe51__lane3_strm0_cntl       ),      
               .std__pe51__lane3_strm0_data          ( std__pe51__lane3_strm0_data       ),      
               .std__pe51__lane3_strm0_data_valid    ( std__pe51__lane3_strm0_data_valid ),      
               .std__pe51__lane3_strm0_data_mask     ( std__pe51__lane3_strm0_data_mask  ),      

               .pe51__std__lane3_strm1_ready         ( pe51__std__lane3_strm1_ready      ),      
               .std__pe51__lane3_strm1_cntl          ( std__pe51__lane3_strm1_cntl       ),      
               .std__pe51__lane3_strm1_data          ( std__pe51__lane3_strm1_data       ),      
               .std__pe51__lane3_strm1_data_valid    ( std__pe51__lane3_strm1_data_valid ),      
               .std__pe51__lane3_strm1_data_mask     ( std__pe51__lane3_strm1_data_mask  ),      

               // PE 51, Lane 4                 
               .pe51__std__lane4_strm0_ready         ( pe51__std__lane4_strm0_ready      ),      
               .std__pe51__lane4_strm0_cntl          ( std__pe51__lane4_strm0_cntl       ),      
               .std__pe51__lane4_strm0_data          ( std__pe51__lane4_strm0_data       ),      
               .std__pe51__lane4_strm0_data_valid    ( std__pe51__lane4_strm0_data_valid ),      
               .std__pe51__lane4_strm0_data_mask     ( std__pe51__lane4_strm0_data_mask  ),      

               .pe51__std__lane4_strm1_ready         ( pe51__std__lane4_strm1_ready      ),      
               .std__pe51__lane4_strm1_cntl          ( std__pe51__lane4_strm1_cntl       ),      
               .std__pe51__lane4_strm1_data          ( std__pe51__lane4_strm1_data       ),      
               .std__pe51__lane4_strm1_data_valid    ( std__pe51__lane4_strm1_data_valid ),      
               .std__pe51__lane4_strm1_data_mask     ( std__pe51__lane4_strm1_data_mask  ),      

               // PE 51, Lane 5                 
               .pe51__std__lane5_strm0_ready         ( pe51__std__lane5_strm0_ready      ),      
               .std__pe51__lane5_strm0_cntl          ( std__pe51__lane5_strm0_cntl       ),      
               .std__pe51__lane5_strm0_data          ( std__pe51__lane5_strm0_data       ),      
               .std__pe51__lane5_strm0_data_valid    ( std__pe51__lane5_strm0_data_valid ),      
               .std__pe51__lane5_strm0_data_mask     ( std__pe51__lane5_strm0_data_mask  ),      

               .pe51__std__lane5_strm1_ready         ( pe51__std__lane5_strm1_ready      ),      
               .std__pe51__lane5_strm1_cntl          ( std__pe51__lane5_strm1_cntl       ),      
               .std__pe51__lane5_strm1_data          ( std__pe51__lane5_strm1_data       ),      
               .std__pe51__lane5_strm1_data_valid    ( std__pe51__lane5_strm1_data_valid ),      
               .std__pe51__lane5_strm1_data_mask     ( std__pe51__lane5_strm1_data_mask  ),      

               // PE 51, Lane 6                 
               .pe51__std__lane6_strm0_ready         ( pe51__std__lane6_strm0_ready      ),      
               .std__pe51__lane6_strm0_cntl          ( std__pe51__lane6_strm0_cntl       ),      
               .std__pe51__lane6_strm0_data          ( std__pe51__lane6_strm0_data       ),      
               .std__pe51__lane6_strm0_data_valid    ( std__pe51__lane6_strm0_data_valid ),      
               .std__pe51__lane6_strm0_data_mask     ( std__pe51__lane6_strm0_data_mask  ),      

               .pe51__std__lane6_strm1_ready         ( pe51__std__lane6_strm1_ready      ),      
               .std__pe51__lane6_strm1_cntl          ( std__pe51__lane6_strm1_cntl       ),      
               .std__pe51__lane6_strm1_data          ( std__pe51__lane6_strm1_data       ),      
               .std__pe51__lane6_strm1_data_valid    ( std__pe51__lane6_strm1_data_valid ),      
               .std__pe51__lane6_strm1_data_mask     ( std__pe51__lane6_strm1_data_mask  ),      

               // PE 51, Lane 7                 
               .pe51__std__lane7_strm0_ready         ( pe51__std__lane7_strm0_ready      ),      
               .std__pe51__lane7_strm0_cntl          ( std__pe51__lane7_strm0_cntl       ),      
               .std__pe51__lane7_strm0_data          ( std__pe51__lane7_strm0_data       ),      
               .std__pe51__lane7_strm0_data_valid    ( std__pe51__lane7_strm0_data_valid ),      
               .std__pe51__lane7_strm0_data_mask     ( std__pe51__lane7_strm0_data_mask  ),      

               .pe51__std__lane7_strm1_ready         ( pe51__std__lane7_strm1_ready      ),      
               .std__pe51__lane7_strm1_cntl          ( std__pe51__lane7_strm1_cntl       ),      
               .std__pe51__lane7_strm1_data          ( std__pe51__lane7_strm1_data       ),      
               .std__pe51__lane7_strm1_data_valid    ( std__pe51__lane7_strm1_data_valid ),      
               .std__pe51__lane7_strm1_data_mask     ( std__pe51__lane7_strm1_data_mask  ),      

               // PE 51, Lane 8                 
               .pe51__std__lane8_strm0_ready         ( pe51__std__lane8_strm0_ready      ),      
               .std__pe51__lane8_strm0_cntl          ( std__pe51__lane8_strm0_cntl       ),      
               .std__pe51__lane8_strm0_data          ( std__pe51__lane8_strm0_data       ),      
               .std__pe51__lane8_strm0_data_valid    ( std__pe51__lane8_strm0_data_valid ),      
               .std__pe51__lane8_strm0_data_mask     ( std__pe51__lane8_strm0_data_mask  ),      

               .pe51__std__lane8_strm1_ready         ( pe51__std__lane8_strm1_ready      ),      
               .std__pe51__lane8_strm1_cntl          ( std__pe51__lane8_strm1_cntl       ),      
               .std__pe51__lane8_strm1_data          ( std__pe51__lane8_strm1_data       ),      
               .std__pe51__lane8_strm1_data_valid    ( std__pe51__lane8_strm1_data_valid ),      
               .std__pe51__lane8_strm1_data_mask     ( std__pe51__lane8_strm1_data_mask  ),      

               // PE 51, Lane 9                 
               .pe51__std__lane9_strm0_ready         ( pe51__std__lane9_strm0_ready      ),      
               .std__pe51__lane9_strm0_cntl          ( std__pe51__lane9_strm0_cntl       ),      
               .std__pe51__lane9_strm0_data          ( std__pe51__lane9_strm0_data       ),      
               .std__pe51__lane9_strm0_data_valid    ( std__pe51__lane9_strm0_data_valid ),      
               .std__pe51__lane9_strm0_data_mask     ( std__pe51__lane9_strm0_data_mask  ),      

               .pe51__std__lane9_strm1_ready         ( pe51__std__lane9_strm1_ready      ),      
               .std__pe51__lane9_strm1_cntl          ( std__pe51__lane9_strm1_cntl       ),      
               .std__pe51__lane9_strm1_data          ( std__pe51__lane9_strm1_data       ),      
               .std__pe51__lane9_strm1_data_valid    ( std__pe51__lane9_strm1_data_valid ),      
               .std__pe51__lane9_strm1_data_mask     ( std__pe51__lane9_strm1_data_mask  ),      

               // PE 51, Lane 10                 
               .pe51__std__lane10_strm0_ready         ( pe51__std__lane10_strm0_ready      ),      
               .std__pe51__lane10_strm0_cntl          ( std__pe51__lane10_strm0_cntl       ),      
               .std__pe51__lane10_strm0_data          ( std__pe51__lane10_strm0_data       ),      
               .std__pe51__lane10_strm0_data_valid    ( std__pe51__lane10_strm0_data_valid ),      
               .std__pe51__lane10_strm0_data_mask     ( std__pe51__lane10_strm0_data_mask  ),      

               .pe51__std__lane10_strm1_ready         ( pe51__std__lane10_strm1_ready      ),      
               .std__pe51__lane10_strm1_cntl          ( std__pe51__lane10_strm1_cntl       ),      
               .std__pe51__lane10_strm1_data          ( std__pe51__lane10_strm1_data       ),      
               .std__pe51__lane10_strm1_data_valid    ( std__pe51__lane10_strm1_data_valid ),      
               .std__pe51__lane10_strm1_data_mask     ( std__pe51__lane10_strm1_data_mask  ),      

               // PE 51, Lane 11                 
               .pe51__std__lane11_strm0_ready         ( pe51__std__lane11_strm0_ready      ),      
               .std__pe51__lane11_strm0_cntl          ( std__pe51__lane11_strm0_cntl       ),      
               .std__pe51__lane11_strm0_data          ( std__pe51__lane11_strm0_data       ),      
               .std__pe51__lane11_strm0_data_valid    ( std__pe51__lane11_strm0_data_valid ),      
               .std__pe51__lane11_strm0_data_mask     ( std__pe51__lane11_strm0_data_mask  ),      

               .pe51__std__lane11_strm1_ready         ( pe51__std__lane11_strm1_ready      ),      
               .std__pe51__lane11_strm1_cntl          ( std__pe51__lane11_strm1_cntl       ),      
               .std__pe51__lane11_strm1_data          ( std__pe51__lane11_strm1_data       ),      
               .std__pe51__lane11_strm1_data_valid    ( std__pe51__lane11_strm1_data_valid ),      
               .std__pe51__lane11_strm1_data_mask     ( std__pe51__lane11_strm1_data_mask  ),      

               // PE 51, Lane 12                 
               .pe51__std__lane12_strm0_ready         ( pe51__std__lane12_strm0_ready      ),      
               .std__pe51__lane12_strm0_cntl          ( std__pe51__lane12_strm0_cntl       ),      
               .std__pe51__lane12_strm0_data          ( std__pe51__lane12_strm0_data       ),      
               .std__pe51__lane12_strm0_data_valid    ( std__pe51__lane12_strm0_data_valid ),      
               .std__pe51__lane12_strm0_data_mask     ( std__pe51__lane12_strm0_data_mask  ),      

               .pe51__std__lane12_strm1_ready         ( pe51__std__lane12_strm1_ready      ),      
               .std__pe51__lane12_strm1_cntl          ( std__pe51__lane12_strm1_cntl       ),      
               .std__pe51__lane12_strm1_data          ( std__pe51__lane12_strm1_data       ),      
               .std__pe51__lane12_strm1_data_valid    ( std__pe51__lane12_strm1_data_valid ),      
               .std__pe51__lane12_strm1_data_mask     ( std__pe51__lane12_strm1_data_mask  ),      

               // PE 51, Lane 13                 
               .pe51__std__lane13_strm0_ready         ( pe51__std__lane13_strm0_ready      ),      
               .std__pe51__lane13_strm0_cntl          ( std__pe51__lane13_strm0_cntl       ),      
               .std__pe51__lane13_strm0_data          ( std__pe51__lane13_strm0_data       ),      
               .std__pe51__lane13_strm0_data_valid    ( std__pe51__lane13_strm0_data_valid ),      
               .std__pe51__lane13_strm0_data_mask     ( std__pe51__lane13_strm0_data_mask  ),      

               .pe51__std__lane13_strm1_ready         ( pe51__std__lane13_strm1_ready      ),      
               .std__pe51__lane13_strm1_cntl          ( std__pe51__lane13_strm1_cntl       ),      
               .std__pe51__lane13_strm1_data          ( std__pe51__lane13_strm1_data       ),      
               .std__pe51__lane13_strm1_data_valid    ( std__pe51__lane13_strm1_data_valid ),      
               .std__pe51__lane13_strm1_data_mask     ( std__pe51__lane13_strm1_data_mask  ),      

               // PE 51, Lane 14                 
               .pe51__std__lane14_strm0_ready         ( pe51__std__lane14_strm0_ready      ),      
               .std__pe51__lane14_strm0_cntl          ( std__pe51__lane14_strm0_cntl       ),      
               .std__pe51__lane14_strm0_data          ( std__pe51__lane14_strm0_data       ),      
               .std__pe51__lane14_strm0_data_valid    ( std__pe51__lane14_strm0_data_valid ),      
               .std__pe51__lane14_strm0_data_mask     ( std__pe51__lane14_strm0_data_mask  ),      

               .pe51__std__lane14_strm1_ready         ( pe51__std__lane14_strm1_ready      ),      
               .std__pe51__lane14_strm1_cntl          ( std__pe51__lane14_strm1_cntl       ),      
               .std__pe51__lane14_strm1_data          ( std__pe51__lane14_strm1_data       ),      
               .std__pe51__lane14_strm1_data_valid    ( std__pe51__lane14_strm1_data_valid ),      
               .std__pe51__lane14_strm1_data_mask     ( std__pe51__lane14_strm1_data_mask  ),      

               // PE 51, Lane 15                 
               .pe51__std__lane15_strm0_ready         ( pe51__std__lane15_strm0_ready      ),      
               .std__pe51__lane15_strm0_cntl          ( std__pe51__lane15_strm0_cntl       ),      
               .std__pe51__lane15_strm0_data          ( std__pe51__lane15_strm0_data       ),      
               .std__pe51__lane15_strm0_data_valid    ( std__pe51__lane15_strm0_data_valid ),      
               .std__pe51__lane15_strm0_data_mask     ( std__pe51__lane15_strm0_data_mask  ),      

               .pe51__std__lane15_strm1_ready         ( pe51__std__lane15_strm1_ready      ),      
               .std__pe51__lane15_strm1_cntl          ( std__pe51__lane15_strm1_cntl       ),      
               .std__pe51__lane15_strm1_data          ( std__pe51__lane15_strm1_data       ),      
               .std__pe51__lane15_strm1_data_valid    ( std__pe51__lane15_strm1_data_valid ),      
               .std__pe51__lane15_strm1_data_mask     ( std__pe51__lane15_strm1_data_mask  ),      

               // PE 51, Lane 16                 
               .pe51__std__lane16_strm0_ready         ( pe51__std__lane16_strm0_ready      ),      
               .std__pe51__lane16_strm0_cntl          ( std__pe51__lane16_strm0_cntl       ),      
               .std__pe51__lane16_strm0_data          ( std__pe51__lane16_strm0_data       ),      
               .std__pe51__lane16_strm0_data_valid    ( std__pe51__lane16_strm0_data_valid ),      
               .std__pe51__lane16_strm0_data_mask     ( std__pe51__lane16_strm0_data_mask  ),      

               .pe51__std__lane16_strm1_ready         ( pe51__std__lane16_strm1_ready      ),      
               .std__pe51__lane16_strm1_cntl          ( std__pe51__lane16_strm1_cntl       ),      
               .std__pe51__lane16_strm1_data          ( std__pe51__lane16_strm1_data       ),      
               .std__pe51__lane16_strm1_data_valid    ( std__pe51__lane16_strm1_data_valid ),      
               .std__pe51__lane16_strm1_data_mask     ( std__pe51__lane16_strm1_data_mask  ),      

               // PE 51, Lane 17                 
               .pe51__std__lane17_strm0_ready         ( pe51__std__lane17_strm0_ready      ),      
               .std__pe51__lane17_strm0_cntl          ( std__pe51__lane17_strm0_cntl       ),      
               .std__pe51__lane17_strm0_data          ( std__pe51__lane17_strm0_data       ),      
               .std__pe51__lane17_strm0_data_valid    ( std__pe51__lane17_strm0_data_valid ),      
               .std__pe51__lane17_strm0_data_mask     ( std__pe51__lane17_strm0_data_mask  ),      

               .pe51__std__lane17_strm1_ready         ( pe51__std__lane17_strm1_ready      ),      
               .std__pe51__lane17_strm1_cntl          ( std__pe51__lane17_strm1_cntl       ),      
               .std__pe51__lane17_strm1_data          ( std__pe51__lane17_strm1_data       ),      
               .std__pe51__lane17_strm1_data_valid    ( std__pe51__lane17_strm1_data_valid ),      
               .std__pe51__lane17_strm1_data_mask     ( std__pe51__lane17_strm1_data_mask  ),      

               // PE 51, Lane 18                 
               .pe51__std__lane18_strm0_ready         ( pe51__std__lane18_strm0_ready      ),      
               .std__pe51__lane18_strm0_cntl          ( std__pe51__lane18_strm0_cntl       ),      
               .std__pe51__lane18_strm0_data          ( std__pe51__lane18_strm0_data       ),      
               .std__pe51__lane18_strm0_data_valid    ( std__pe51__lane18_strm0_data_valid ),      
               .std__pe51__lane18_strm0_data_mask     ( std__pe51__lane18_strm0_data_mask  ),      

               .pe51__std__lane18_strm1_ready         ( pe51__std__lane18_strm1_ready      ),      
               .std__pe51__lane18_strm1_cntl          ( std__pe51__lane18_strm1_cntl       ),      
               .std__pe51__lane18_strm1_data          ( std__pe51__lane18_strm1_data       ),      
               .std__pe51__lane18_strm1_data_valid    ( std__pe51__lane18_strm1_data_valid ),      
               .std__pe51__lane18_strm1_data_mask     ( std__pe51__lane18_strm1_data_mask  ),      

               // PE 51, Lane 19                 
               .pe51__std__lane19_strm0_ready         ( pe51__std__lane19_strm0_ready      ),      
               .std__pe51__lane19_strm0_cntl          ( std__pe51__lane19_strm0_cntl       ),      
               .std__pe51__lane19_strm0_data          ( std__pe51__lane19_strm0_data       ),      
               .std__pe51__lane19_strm0_data_valid    ( std__pe51__lane19_strm0_data_valid ),      
               .std__pe51__lane19_strm0_data_mask     ( std__pe51__lane19_strm0_data_mask  ),      

               .pe51__std__lane19_strm1_ready         ( pe51__std__lane19_strm1_ready      ),      
               .std__pe51__lane19_strm1_cntl          ( std__pe51__lane19_strm1_cntl       ),      
               .std__pe51__lane19_strm1_data          ( std__pe51__lane19_strm1_data       ),      
               .std__pe51__lane19_strm1_data_valid    ( std__pe51__lane19_strm1_data_valid ),      
               .std__pe51__lane19_strm1_data_mask     ( std__pe51__lane19_strm1_data_mask  ),      

               // PE 51, Lane 20                 
               .pe51__std__lane20_strm0_ready         ( pe51__std__lane20_strm0_ready      ),      
               .std__pe51__lane20_strm0_cntl          ( std__pe51__lane20_strm0_cntl       ),      
               .std__pe51__lane20_strm0_data          ( std__pe51__lane20_strm0_data       ),      
               .std__pe51__lane20_strm0_data_valid    ( std__pe51__lane20_strm0_data_valid ),      
               .std__pe51__lane20_strm0_data_mask     ( std__pe51__lane20_strm0_data_mask  ),      

               .pe51__std__lane20_strm1_ready         ( pe51__std__lane20_strm1_ready      ),      
               .std__pe51__lane20_strm1_cntl          ( std__pe51__lane20_strm1_cntl       ),      
               .std__pe51__lane20_strm1_data          ( std__pe51__lane20_strm1_data       ),      
               .std__pe51__lane20_strm1_data_valid    ( std__pe51__lane20_strm1_data_valid ),      
               .std__pe51__lane20_strm1_data_mask     ( std__pe51__lane20_strm1_data_mask  ),      

               // PE 51, Lane 21                 
               .pe51__std__lane21_strm0_ready         ( pe51__std__lane21_strm0_ready      ),      
               .std__pe51__lane21_strm0_cntl          ( std__pe51__lane21_strm0_cntl       ),      
               .std__pe51__lane21_strm0_data          ( std__pe51__lane21_strm0_data       ),      
               .std__pe51__lane21_strm0_data_valid    ( std__pe51__lane21_strm0_data_valid ),      
               .std__pe51__lane21_strm0_data_mask     ( std__pe51__lane21_strm0_data_mask  ),      

               .pe51__std__lane21_strm1_ready         ( pe51__std__lane21_strm1_ready      ),      
               .std__pe51__lane21_strm1_cntl          ( std__pe51__lane21_strm1_cntl       ),      
               .std__pe51__lane21_strm1_data          ( std__pe51__lane21_strm1_data       ),      
               .std__pe51__lane21_strm1_data_valid    ( std__pe51__lane21_strm1_data_valid ),      
               .std__pe51__lane21_strm1_data_mask     ( std__pe51__lane21_strm1_data_mask  ),      

               // PE 51, Lane 22                 
               .pe51__std__lane22_strm0_ready         ( pe51__std__lane22_strm0_ready      ),      
               .std__pe51__lane22_strm0_cntl          ( std__pe51__lane22_strm0_cntl       ),      
               .std__pe51__lane22_strm0_data          ( std__pe51__lane22_strm0_data       ),      
               .std__pe51__lane22_strm0_data_valid    ( std__pe51__lane22_strm0_data_valid ),      
               .std__pe51__lane22_strm0_data_mask     ( std__pe51__lane22_strm0_data_mask  ),      

               .pe51__std__lane22_strm1_ready         ( pe51__std__lane22_strm1_ready      ),      
               .std__pe51__lane22_strm1_cntl          ( std__pe51__lane22_strm1_cntl       ),      
               .std__pe51__lane22_strm1_data          ( std__pe51__lane22_strm1_data       ),      
               .std__pe51__lane22_strm1_data_valid    ( std__pe51__lane22_strm1_data_valid ),      
               .std__pe51__lane22_strm1_data_mask     ( std__pe51__lane22_strm1_data_mask  ),      

               // PE 51, Lane 23                 
               .pe51__std__lane23_strm0_ready         ( pe51__std__lane23_strm0_ready      ),      
               .std__pe51__lane23_strm0_cntl          ( std__pe51__lane23_strm0_cntl       ),      
               .std__pe51__lane23_strm0_data          ( std__pe51__lane23_strm0_data       ),      
               .std__pe51__lane23_strm0_data_valid    ( std__pe51__lane23_strm0_data_valid ),      
               .std__pe51__lane23_strm0_data_mask     ( std__pe51__lane23_strm0_data_mask  ),      

               .pe51__std__lane23_strm1_ready         ( pe51__std__lane23_strm1_ready      ),      
               .std__pe51__lane23_strm1_cntl          ( std__pe51__lane23_strm1_cntl       ),      
               .std__pe51__lane23_strm1_data          ( std__pe51__lane23_strm1_data       ),      
               .std__pe51__lane23_strm1_data_valid    ( std__pe51__lane23_strm1_data_valid ),      
               .std__pe51__lane23_strm1_data_mask     ( std__pe51__lane23_strm1_data_mask  ),      

               // PE 51, Lane 24                 
               .pe51__std__lane24_strm0_ready         ( pe51__std__lane24_strm0_ready      ),      
               .std__pe51__lane24_strm0_cntl          ( std__pe51__lane24_strm0_cntl       ),      
               .std__pe51__lane24_strm0_data          ( std__pe51__lane24_strm0_data       ),      
               .std__pe51__lane24_strm0_data_valid    ( std__pe51__lane24_strm0_data_valid ),      
               .std__pe51__lane24_strm0_data_mask     ( std__pe51__lane24_strm0_data_mask  ),      

               .pe51__std__lane24_strm1_ready         ( pe51__std__lane24_strm1_ready      ),      
               .std__pe51__lane24_strm1_cntl          ( std__pe51__lane24_strm1_cntl       ),      
               .std__pe51__lane24_strm1_data          ( std__pe51__lane24_strm1_data       ),      
               .std__pe51__lane24_strm1_data_valid    ( std__pe51__lane24_strm1_data_valid ),      
               .std__pe51__lane24_strm1_data_mask     ( std__pe51__lane24_strm1_data_mask  ),      

               // PE 51, Lane 25                 
               .pe51__std__lane25_strm0_ready         ( pe51__std__lane25_strm0_ready      ),      
               .std__pe51__lane25_strm0_cntl          ( std__pe51__lane25_strm0_cntl       ),      
               .std__pe51__lane25_strm0_data          ( std__pe51__lane25_strm0_data       ),      
               .std__pe51__lane25_strm0_data_valid    ( std__pe51__lane25_strm0_data_valid ),      
               .std__pe51__lane25_strm0_data_mask     ( std__pe51__lane25_strm0_data_mask  ),      

               .pe51__std__lane25_strm1_ready         ( pe51__std__lane25_strm1_ready      ),      
               .std__pe51__lane25_strm1_cntl          ( std__pe51__lane25_strm1_cntl       ),      
               .std__pe51__lane25_strm1_data          ( std__pe51__lane25_strm1_data       ),      
               .std__pe51__lane25_strm1_data_valid    ( std__pe51__lane25_strm1_data_valid ),      
               .std__pe51__lane25_strm1_data_mask     ( std__pe51__lane25_strm1_data_mask  ),      

               // PE 51, Lane 26                 
               .pe51__std__lane26_strm0_ready         ( pe51__std__lane26_strm0_ready      ),      
               .std__pe51__lane26_strm0_cntl          ( std__pe51__lane26_strm0_cntl       ),      
               .std__pe51__lane26_strm0_data          ( std__pe51__lane26_strm0_data       ),      
               .std__pe51__lane26_strm0_data_valid    ( std__pe51__lane26_strm0_data_valid ),      
               .std__pe51__lane26_strm0_data_mask     ( std__pe51__lane26_strm0_data_mask  ),      

               .pe51__std__lane26_strm1_ready         ( pe51__std__lane26_strm1_ready      ),      
               .std__pe51__lane26_strm1_cntl          ( std__pe51__lane26_strm1_cntl       ),      
               .std__pe51__lane26_strm1_data          ( std__pe51__lane26_strm1_data       ),      
               .std__pe51__lane26_strm1_data_valid    ( std__pe51__lane26_strm1_data_valid ),      
               .std__pe51__lane26_strm1_data_mask     ( std__pe51__lane26_strm1_data_mask  ),      

               // PE 51, Lane 27                 
               .pe51__std__lane27_strm0_ready         ( pe51__std__lane27_strm0_ready      ),      
               .std__pe51__lane27_strm0_cntl          ( std__pe51__lane27_strm0_cntl       ),      
               .std__pe51__lane27_strm0_data          ( std__pe51__lane27_strm0_data       ),      
               .std__pe51__lane27_strm0_data_valid    ( std__pe51__lane27_strm0_data_valid ),      
               .std__pe51__lane27_strm0_data_mask     ( std__pe51__lane27_strm0_data_mask  ),      

               .pe51__std__lane27_strm1_ready         ( pe51__std__lane27_strm1_ready      ),      
               .std__pe51__lane27_strm1_cntl          ( std__pe51__lane27_strm1_cntl       ),      
               .std__pe51__lane27_strm1_data          ( std__pe51__lane27_strm1_data       ),      
               .std__pe51__lane27_strm1_data_valid    ( std__pe51__lane27_strm1_data_valid ),      
               .std__pe51__lane27_strm1_data_mask     ( std__pe51__lane27_strm1_data_mask  ),      

               // PE 51, Lane 28                 
               .pe51__std__lane28_strm0_ready         ( pe51__std__lane28_strm0_ready      ),      
               .std__pe51__lane28_strm0_cntl          ( std__pe51__lane28_strm0_cntl       ),      
               .std__pe51__lane28_strm0_data          ( std__pe51__lane28_strm0_data       ),      
               .std__pe51__lane28_strm0_data_valid    ( std__pe51__lane28_strm0_data_valid ),      
               .std__pe51__lane28_strm0_data_mask     ( std__pe51__lane28_strm0_data_mask  ),      

               .pe51__std__lane28_strm1_ready         ( pe51__std__lane28_strm1_ready      ),      
               .std__pe51__lane28_strm1_cntl          ( std__pe51__lane28_strm1_cntl       ),      
               .std__pe51__lane28_strm1_data          ( std__pe51__lane28_strm1_data       ),      
               .std__pe51__lane28_strm1_data_valid    ( std__pe51__lane28_strm1_data_valid ),      
               .std__pe51__lane28_strm1_data_mask     ( std__pe51__lane28_strm1_data_mask  ),      

               // PE 51, Lane 29                 
               .pe51__std__lane29_strm0_ready         ( pe51__std__lane29_strm0_ready      ),      
               .std__pe51__lane29_strm0_cntl          ( std__pe51__lane29_strm0_cntl       ),      
               .std__pe51__lane29_strm0_data          ( std__pe51__lane29_strm0_data       ),      
               .std__pe51__lane29_strm0_data_valid    ( std__pe51__lane29_strm0_data_valid ),      
               .std__pe51__lane29_strm0_data_mask     ( std__pe51__lane29_strm0_data_mask  ),      

               .pe51__std__lane29_strm1_ready         ( pe51__std__lane29_strm1_ready      ),      
               .std__pe51__lane29_strm1_cntl          ( std__pe51__lane29_strm1_cntl       ),      
               .std__pe51__lane29_strm1_data          ( std__pe51__lane29_strm1_data       ),      
               .std__pe51__lane29_strm1_data_valid    ( std__pe51__lane29_strm1_data_valid ),      
               .std__pe51__lane29_strm1_data_mask     ( std__pe51__lane29_strm1_data_mask  ),      

               // PE 51, Lane 30                 
               .pe51__std__lane30_strm0_ready         ( pe51__std__lane30_strm0_ready      ),      
               .std__pe51__lane30_strm0_cntl          ( std__pe51__lane30_strm0_cntl       ),      
               .std__pe51__lane30_strm0_data          ( std__pe51__lane30_strm0_data       ),      
               .std__pe51__lane30_strm0_data_valid    ( std__pe51__lane30_strm0_data_valid ),      
               .std__pe51__lane30_strm0_data_mask     ( std__pe51__lane30_strm0_data_mask  ),      

               .pe51__std__lane30_strm1_ready         ( pe51__std__lane30_strm1_ready      ),      
               .std__pe51__lane30_strm1_cntl          ( std__pe51__lane30_strm1_cntl       ),      
               .std__pe51__lane30_strm1_data          ( std__pe51__lane30_strm1_data       ),      
               .std__pe51__lane30_strm1_data_valid    ( std__pe51__lane30_strm1_data_valid ),      
               .std__pe51__lane30_strm1_data_mask     ( std__pe51__lane30_strm1_data_mask  ),      

               // PE 51, Lane 31                 
               .pe51__std__lane31_strm0_ready         ( pe51__std__lane31_strm0_ready      ),      
               .std__pe51__lane31_strm0_cntl          ( std__pe51__lane31_strm0_cntl       ),      
               .std__pe51__lane31_strm0_data          ( std__pe51__lane31_strm0_data       ),      
               .std__pe51__lane31_strm0_data_valid    ( std__pe51__lane31_strm0_data_valid ),      
               .std__pe51__lane31_strm0_data_mask     ( std__pe51__lane31_strm0_data_mask  ),      

               .pe51__std__lane31_strm1_ready         ( pe51__std__lane31_strm1_ready      ),      
               .std__pe51__lane31_strm1_cntl          ( std__pe51__lane31_strm1_cntl       ),      
               .std__pe51__lane31_strm1_data          ( std__pe51__lane31_strm1_data       ),      
               .std__pe51__lane31_strm1_data_valid    ( std__pe51__lane31_strm1_data_valid ),      
               .std__pe51__lane31_strm1_data_mask     ( std__pe51__lane31_strm1_data_mask  ),      

               // PE 52, Lane 0                 
               .pe52__std__lane0_strm0_ready         ( pe52__std__lane0_strm0_ready      ),      
               .std__pe52__lane0_strm0_cntl          ( std__pe52__lane0_strm0_cntl       ),      
               .std__pe52__lane0_strm0_data          ( std__pe52__lane0_strm0_data       ),      
               .std__pe52__lane0_strm0_data_valid    ( std__pe52__lane0_strm0_data_valid ),      
               .std__pe52__lane0_strm0_data_mask     ( std__pe52__lane0_strm0_data_mask  ),      

               .pe52__std__lane0_strm1_ready         ( pe52__std__lane0_strm1_ready      ),      
               .std__pe52__lane0_strm1_cntl          ( std__pe52__lane0_strm1_cntl       ),      
               .std__pe52__lane0_strm1_data          ( std__pe52__lane0_strm1_data       ),      
               .std__pe52__lane0_strm1_data_valid    ( std__pe52__lane0_strm1_data_valid ),      
               .std__pe52__lane0_strm1_data_mask     ( std__pe52__lane0_strm1_data_mask  ),      

               // PE 52, Lane 1                 
               .pe52__std__lane1_strm0_ready         ( pe52__std__lane1_strm0_ready      ),      
               .std__pe52__lane1_strm0_cntl          ( std__pe52__lane1_strm0_cntl       ),      
               .std__pe52__lane1_strm0_data          ( std__pe52__lane1_strm0_data       ),      
               .std__pe52__lane1_strm0_data_valid    ( std__pe52__lane1_strm0_data_valid ),      
               .std__pe52__lane1_strm0_data_mask     ( std__pe52__lane1_strm0_data_mask  ),      

               .pe52__std__lane1_strm1_ready         ( pe52__std__lane1_strm1_ready      ),      
               .std__pe52__lane1_strm1_cntl          ( std__pe52__lane1_strm1_cntl       ),      
               .std__pe52__lane1_strm1_data          ( std__pe52__lane1_strm1_data       ),      
               .std__pe52__lane1_strm1_data_valid    ( std__pe52__lane1_strm1_data_valid ),      
               .std__pe52__lane1_strm1_data_mask     ( std__pe52__lane1_strm1_data_mask  ),      

               // PE 52, Lane 2                 
               .pe52__std__lane2_strm0_ready         ( pe52__std__lane2_strm0_ready      ),      
               .std__pe52__lane2_strm0_cntl          ( std__pe52__lane2_strm0_cntl       ),      
               .std__pe52__lane2_strm0_data          ( std__pe52__lane2_strm0_data       ),      
               .std__pe52__lane2_strm0_data_valid    ( std__pe52__lane2_strm0_data_valid ),      
               .std__pe52__lane2_strm0_data_mask     ( std__pe52__lane2_strm0_data_mask  ),      

               .pe52__std__lane2_strm1_ready         ( pe52__std__lane2_strm1_ready      ),      
               .std__pe52__lane2_strm1_cntl          ( std__pe52__lane2_strm1_cntl       ),      
               .std__pe52__lane2_strm1_data          ( std__pe52__lane2_strm1_data       ),      
               .std__pe52__lane2_strm1_data_valid    ( std__pe52__lane2_strm1_data_valid ),      
               .std__pe52__lane2_strm1_data_mask     ( std__pe52__lane2_strm1_data_mask  ),      

               // PE 52, Lane 3                 
               .pe52__std__lane3_strm0_ready         ( pe52__std__lane3_strm0_ready      ),      
               .std__pe52__lane3_strm0_cntl          ( std__pe52__lane3_strm0_cntl       ),      
               .std__pe52__lane3_strm0_data          ( std__pe52__lane3_strm0_data       ),      
               .std__pe52__lane3_strm0_data_valid    ( std__pe52__lane3_strm0_data_valid ),      
               .std__pe52__lane3_strm0_data_mask     ( std__pe52__lane3_strm0_data_mask  ),      

               .pe52__std__lane3_strm1_ready         ( pe52__std__lane3_strm1_ready      ),      
               .std__pe52__lane3_strm1_cntl          ( std__pe52__lane3_strm1_cntl       ),      
               .std__pe52__lane3_strm1_data          ( std__pe52__lane3_strm1_data       ),      
               .std__pe52__lane3_strm1_data_valid    ( std__pe52__lane3_strm1_data_valid ),      
               .std__pe52__lane3_strm1_data_mask     ( std__pe52__lane3_strm1_data_mask  ),      

               // PE 52, Lane 4                 
               .pe52__std__lane4_strm0_ready         ( pe52__std__lane4_strm0_ready      ),      
               .std__pe52__lane4_strm0_cntl          ( std__pe52__lane4_strm0_cntl       ),      
               .std__pe52__lane4_strm0_data          ( std__pe52__lane4_strm0_data       ),      
               .std__pe52__lane4_strm0_data_valid    ( std__pe52__lane4_strm0_data_valid ),      
               .std__pe52__lane4_strm0_data_mask     ( std__pe52__lane4_strm0_data_mask  ),      

               .pe52__std__lane4_strm1_ready         ( pe52__std__lane4_strm1_ready      ),      
               .std__pe52__lane4_strm1_cntl          ( std__pe52__lane4_strm1_cntl       ),      
               .std__pe52__lane4_strm1_data          ( std__pe52__lane4_strm1_data       ),      
               .std__pe52__lane4_strm1_data_valid    ( std__pe52__lane4_strm1_data_valid ),      
               .std__pe52__lane4_strm1_data_mask     ( std__pe52__lane4_strm1_data_mask  ),      

               // PE 52, Lane 5                 
               .pe52__std__lane5_strm0_ready         ( pe52__std__lane5_strm0_ready      ),      
               .std__pe52__lane5_strm0_cntl          ( std__pe52__lane5_strm0_cntl       ),      
               .std__pe52__lane5_strm0_data          ( std__pe52__lane5_strm0_data       ),      
               .std__pe52__lane5_strm0_data_valid    ( std__pe52__lane5_strm0_data_valid ),      
               .std__pe52__lane5_strm0_data_mask     ( std__pe52__lane5_strm0_data_mask  ),      

               .pe52__std__lane5_strm1_ready         ( pe52__std__lane5_strm1_ready      ),      
               .std__pe52__lane5_strm1_cntl          ( std__pe52__lane5_strm1_cntl       ),      
               .std__pe52__lane5_strm1_data          ( std__pe52__lane5_strm1_data       ),      
               .std__pe52__lane5_strm1_data_valid    ( std__pe52__lane5_strm1_data_valid ),      
               .std__pe52__lane5_strm1_data_mask     ( std__pe52__lane5_strm1_data_mask  ),      

               // PE 52, Lane 6                 
               .pe52__std__lane6_strm0_ready         ( pe52__std__lane6_strm0_ready      ),      
               .std__pe52__lane6_strm0_cntl          ( std__pe52__lane6_strm0_cntl       ),      
               .std__pe52__lane6_strm0_data          ( std__pe52__lane6_strm0_data       ),      
               .std__pe52__lane6_strm0_data_valid    ( std__pe52__lane6_strm0_data_valid ),      
               .std__pe52__lane6_strm0_data_mask     ( std__pe52__lane6_strm0_data_mask  ),      

               .pe52__std__lane6_strm1_ready         ( pe52__std__lane6_strm1_ready      ),      
               .std__pe52__lane6_strm1_cntl          ( std__pe52__lane6_strm1_cntl       ),      
               .std__pe52__lane6_strm1_data          ( std__pe52__lane6_strm1_data       ),      
               .std__pe52__lane6_strm1_data_valid    ( std__pe52__lane6_strm1_data_valid ),      
               .std__pe52__lane6_strm1_data_mask     ( std__pe52__lane6_strm1_data_mask  ),      

               // PE 52, Lane 7                 
               .pe52__std__lane7_strm0_ready         ( pe52__std__lane7_strm0_ready      ),      
               .std__pe52__lane7_strm0_cntl          ( std__pe52__lane7_strm0_cntl       ),      
               .std__pe52__lane7_strm0_data          ( std__pe52__lane7_strm0_data       ),      
               .std__pe52__lane7_strm0_data_valid    ( std__pe52__lane7_strm0_data_valid ),      
               .std__pe52__lane7_strm0_data_mask     ( std__pe52__lane7_strm0_data_mask  ),      

               .pe52__std__lane7_strm1_ready         ( pe52__std__lane7_strm1_ready      ),      
               .std__pe52__lane7_strm1_cntl          ( std__pe52__lane7_strm1_cntl       ),      
               .std__pe52__lane7_strm1_data          ( std__pe52__lane7_strm1_data       ),      
               .std__pe52__lane7_strm1_data_valid    ( std__pe52__lane7_strm1_data_valid ),      
               .std__pe52__lane7_strm1_data_mask     ( std__pe52__lane7_strm1_data_mask  ),      

               // PE 52, Lane 8                 
               .pe52__std__lane8_strm0_ready         ( pe52__std__lane8_strm0_ready      ),      
               .std__pe52__lane8_strm0_cntl          ( std__pe52__lane8_strm0_cntl       ),      
               .std__pe52__lane8_strm0_data          ( std__pe52__lane8_strm0_data       ),      
               .std__pe52__lane8_strm0_data_valid    ( std__pe52__lane8_strm0_data_valid ),      
               .std__pe52__lane8_strm0_data_mask     ( std__pe52__lane8_strm0_data_mask  ),      

               .pe52__std__lane8_strm1_ready         ( pe52__std__lane8_strm1_ready      ),      
               .std__pe52__lane8_strm1_cntl          ( std__pe52__lane8_strm1_cntl       ),      
               .std__pe52__lane8_strm1_data          ( std__pe52__lane8_strm1_data       ),      
               .std__pe52__lane8_strm1_data_valid    ( std__pe52__lane8_strm1_data_valid ),      
               .std__pe52__lane8_strm1_data_mask     ( std__pe52__lane8_strm1_data_mask  ),      

               // PE 52, Lane 9                 
               .pe52__std__lane9_strm0_ready         ( pe52__std__lane9_strm0_ready      ),      
               .std__pe52__lane9_strm0_cntl          ( std__pe52__lane9_strm0_cntl       ),      
               .std__pe52__lane9_strm0_data          ( std__pe52__lane9_strm0_data       ),      
               .std__pe52__lane9_strm0_data_valid    ( std__pe52__lane9_strm0_data_valid ),      
               .std__pe52__lane9_strm0_data_mask     ( std__pe52__lane9_strm0_data_mask  ),      

               .pe52__std__lane9_strm1_ready         ( pe52__std__lane9_strm1_ready      ),      
               .std__pe52__lane9_strm1_cntl          ( std__pe52__lane9_strm1_cntl       ),      
               .std__pe52__lane9_strm1_data          ( std__pe52__lane9_strm1_data       ),      
               .std__pe52__lane9_strm1_data_valid    ( std__pe52__lane9_strm1_data_valid ),      
               .std__pe52__lane9_strm1_data_mask     ( std__pe52__lane9_strm1_data_mask  ),      

               // PE 52, Lane 10                 
               .pe52__std__lane10_strm0_ready         ( pe52__std__lane10_strm0_ready      ),      
               .std__pe52__lane10_strm0_cntl          ( std__pe52__lane10_strm0_cntl       ),      
               .std__pe52__lane10_strm0_data          ( std__pe52__lane10_strm0_data       ),      
               .std__pe52__lane10_strm0_data_valid    ( std__pe52__lane10_strm0_data_valid ),      
               .std__pe52__lane10_strm0_data_mask     ( std__pe52__lane10_strm0_data_mask  ),      

               .pe52__std__lane10_strm1_ready         ( pe52__std__lane10_strm1_ready      ),      
               .std__pe52__lane10_strm1_cntl          ( std__pe52__lane10_strm1_cntl       ),      
               .std__pe52__lane10_strm1_data          ( std__pe52__lane10_strm1_data       ),      
               .std__pe52__lane10_strm1_data_valid    ( std__pe52__lane10_strm1_data_valid ),      
               .std__pe52__lane10_strm1_data_mask     ( std__pe52__lane10_strm1_data_mask  ),      

               // PE 52, Lane 11                 
               .pe52__std__lane11_strm0_ready         ( pe52__std__lane11_strm0_ready      ),      
               .std__pe52__lane11_strm0_cntl          ( std__pe52__lane11_strm0_cntl       ),      
               .std__pe52__lane11_strm0_data          ( std__pe52__lane11_strm0_data       ),      
               .std__pe52__lane11_strm0_data_valid    ( std__pe52__lane11_strm0_data_valid ),      
               .std__pe52__lane11_strm0_data_mask     ( std__pe52__lane11_strm0_data_mask  ),      

               .pe52__std__lane11_strm1_ready         ( pe52__std__lane11_strm1_ready      ),      
               .std__pe52__lane11_strm1_cntl          ( std__pe52__lane11_strm1_cntl       ),      
               .std__pe52__lane11_strm1_data          ( std__pe52__lane11_strm1_data       ),      
               .std__pe52__lane11_strm1_data_valid    ( std__pe52__lane11_strm1_data_valid ),      
               .std__pe52__lane11_strm1_data_mask     ( std__pe52__lane11_strm1_data_mask  ),      

               // PE 52, Lane 12                 
               .pe52__std__lane12_strm0_ready         ( pe52__std__lane12_strm0_ready      ),      
               .std__pe52__lane12_strm0_cntl          ( std__pe52__lane12_strm0_cntl       ),      
               .std__pe52__lane12_strm0_data          ( std__pe52__lane12_strm0_data       ),      
               .std__pe52__lane12_strm0_data_valid    ( std__pe52__lane12_strm0_data_valid ),      
               .std__pe52__lane12_strm0_data_mask     ( std__pe52__lane12_strm0_data_mask  ),      

               .pe52__std__lane12_strm1_ready         ( pe52__std__lane12_strm1_ready      ),      
               .std__pe52__lane12_strm1_cntl          ( std__pe52__lane12_strm1_cntl       ),      
               .std__pe52__lane12_strm1_data          ( std__pe52__lane12_strm1_data       ),      
               .std__pe52__lane12_strm1_data_valid    ( std__pe52__lane12_strm1_data_valid ),      
               .std__pe52__lane12_strm1_data_mask     ( std__pe52__lane12_strm1_data_mask  ),      

               // PE 52, Lane 13                 
               .pe52__std__lane13_strm0_ready         ( pe52__std__lane13_strm0_ready      ),      
               .std__pe52__lane13_strm0_cntl          ( std__pe52__lane13_strm0_cntl       ),      
               .std__pe52__lane13_strm0_data          ( std__pe52__lane13_strm0_data       ),      
               .std__pe52__lane13_strm0_data_valid    ( std__pe52__lane13_strm0_data_valid ),      
               .std__pe52__lane13_strm0_data_mask     ( std__pe52__lane13_strm0_data_mask  ),      

               .pe52__std__lane13_strm1_ready         ( pe52__std__lane13_strm1_ready      ),      
               .std__pe52__lane13_strm1_cntl          ( std__pe52__lane13_strm1_cntl       ),      
               .std__pe52__lane13_strm1_data          ( std__pe52__lane13_strm1_data       ),      
               .std__pe52__lane13_strm1_data_valid    ( std__pe52__lane13_strm1_data_valid ),      
               .std__pe52__lane13_strm1_data_mask     ( std__pe52__lane13_strm1_data_mask  ),      

               // PE 52, Lane 14                 
               .pe52__std__lane14_strm0_ready         ( pe52__std__lane14_strm0_ready      ),      
               .std__pe52__lane14_strm0_cntl          ( std__pe52__lane14_strm0_cntl       ),      
               .std__pe52__lane14_strm0_data          ( std__pe52__lane14_strm0_data       ),      
               .std__pe52__lane14_strm0_data_valid    ( std__pe52__lane14_strm0_data_valid ),      
               .std__pe52__lane14_strm0_data_mask     ( std__pe52__lane14_strm0_data_mask  ),      

               .pe52__std__lane14_strm1_ready         ( pe52__std__lane14_strm1_ready      ),      
               .std__pe52__lane14_strm1_cntl          ( std__pe52__lane14_strm1_cntl       ),      
               .std__pe52__lane14_strm1_data          ( std__pe52__lane14_strm1_data       ),      
               .std__pe52__lane14_strm1_data_valid    ( std__pe52__lane14_strm1_data_valid ),      
               .std__pe52__lane14_strm1_data_mask     ( std__pe52__lane14_strm1_data_mask  ),      

               // PE 52, Lane 15                 
               .pe52__std__lane15_strm0_ready         ( pe52__std__lane15_strm0_ready      ),      
               .std__pe52__lane15_strm0_cntl          ( std__pe52__lane15_strm0_cntl       ),      
               .std__pe52__lane15_strm0_data          ( std__pe52__lane15_strm0_data       ),      
               .std__pe52__lane15_strm0_data_valid    ( std__pe52__lane15_strm0_data_valid ),      
               .std__pe52__lane15_strm0_data_mask     ( std__pe52__lane15_strm0_data_mask  ),      

               .pe52__std__lane15_strm1_ready         ( pe52__std__lane15_strm1_ready      ),      
               .std__pe52__lane15_strm1_cntl          ( std__pe52__lane15_strm1_cntl       ),      
               .std__pe52__lane15_strm1_data          ( std__pe52__lane15_strm1_data       ),      
               .std__pe52__lane15_strm1_data_valid    ( std__pe52__lane15_strm1_data_valid ),      
               .std__pe52__lane15_strm1_data_mask     ( std__pe52__lane15_strm1_data_mask  ),      

               // PE 52, Lane 16                 
               .pe52__std__lane16_strm0_ready         ( pe52__std__lane16_strm0_ready      ),      
               .std__pe52__lane16_strm0_cntl          ( std__pe52__lane16_strm0_cntl       ),      
               .std__pe52__lane16_strm0_data          ( std__pe52__lane16_strm0_data       ),      
               .std__pe52__lane16_strm0_data_valid    ( std__pe52__lane16_strm0_data_valid ),      
               .std__pe52__lane16_strm0_data_mask     ( std__pe52__lane16_strm0_data_mask  ),      

               .pe52__std__lane16_strm1_ready         ( pe52__std__lane16_strm1_ready      ),      
               .std__pe52__lane16_strm1_cntl          ( std__pe52__lane16_strm1_cntl       ),      
               .std__pe52__lane16_strm1_data          ( std__pe52__lane16_strm1_data       ),      
               .std__pe52__lane16_strm1_data_valid    ( std__pe52__lane16_strm1_data_valid ),      
               .std__pe52__lane16_strm1_data_mask     ( std__pe52__lane16_strm1_data_mask  ),      

               // PE 52, Lane 17                 
               .pe52__std__lane17_strm0_ready         ( pe52__std__lane17_strm0_ready      ),      
               .std__pe52__lane17_strm0_cntl          ( std__pe52__lane17_strm0_cntl       ),      
               .std__pe52__lane17_strm0_data          ( std__pe52__lane17_strm0_data       ),      
               .std__pe52__lane17_strm0_data_valid    ( std__pe52__lane17_strm0_data_valid ),      
               .std__pe52__lane17_strm0_data_mask     ( std__pe52__lane17_strm0_data_mask  ),      

               .pe52__std__lane17_strm1_ready         ( pe52__std__lane17_strm1_ready      ),      
               .std__pe52__lane17_strm1_cntl          ( std__pe52__lane17_strm1_cntl       ),      
               .std__pe52__lane17_strm1_data          ( std__pe52__lane17_strm1_data       ),      
               .std__pe52__lane17_strm1_data_valid    ( std__pe52__lane17_strm1_data_valid ),      
               .std__pe52__lane17_strm1_data_mask     ( std__pe52__lane17_strm1_data_mask  ),      

               // PE 52, Lane 18                 
               .pe52__std__lane18_strm0_ready         ( pe52__std__lane18_strm0_ready      ),      
               .std__pe52__lane18_strm0_cntl          ( std__pe52__lane18_strm0_cntl       ),      
               .std__pe52__lane18_strm0_data          ( std__pe52__lane18_strm0_data       ),      
               .std__pe52__lane18_strm0_data_valid    ( std__pe52__lane18_strm0_data_valid ),      
               .std__pe52__lane18_strm0_data_mask     ( std__pe52__lane18_strm0_data_mask  ),      

               .pe52__std__lane18_strm1_ready         ( pe52__std__lane18_strm1_ready      ),      
               .std__pe52__lane18_strm1_cntl          ( std__pe52__lane18_strm1_cntl       ),      
               .std__pe52__lane18_strm1_data          ( std__pe52__lane18_strm1_data       ),      
               .std__pe52__lane18_strm1_data_valid    ( std__pe52__lane18_strm1_data_valid ),      
               .std__pe52__lane18_strm1_data_mask     ( std__pe52__lane18_strm1_data_mask  ),      

               // PE 52, Lane 19                 
               .pe52__std__lane19_strm0_ready         ( pe52__std__lane19_strm0_ready      ),      
               .std__pe52__lane19_strm0_cntl          ( std__pe52__lane19_strm0_cntl       ),      
               .std__pe52__lane19_strm0_data          ( std__pe52__lane19_strm0_data       ),      
               .std__pe52__lane19_strm0_data_valid    ( std__pe52__lane19_strm0_data_valid ),      
               .std__pe52__lane19_strm0_data_mask     ( std__pe52__lane19_strm0_data_mask  ),      

               .pe52__std__lane19_strm1_ready         ( pe52__std__lane19_strm1_ready      ),      
               .std__pe52__lane19_strm1_cntl          ( std__pe52__lane19_strm1_cntl       ),      
               .std__pe52__lane19_strm1_data          ( std__pe52__lane19_strm1_data       ),      
               .std__pe52__lane19_strm1_data_valid    ( std__pe52__lane19_strm1_data_valid ),      
               .std__pe52__lane19_strm1_data_mask     ( std__pe52__lane19_strm1_data_mask  ),      

               // PE 52, Lane 20                 
               .pe52__std__lane20_strm0_ready         ( pe52__std__lane20_strm0_ready      ),      
               .std__pe52__lane20_strm0_cntl          ( std__pe52__lane20_strm0_cntl       ),      
               .std__pe52__lane20_strm0_data          ( std__pe52__lane20_strm0_data       ),      
               .std__pe52__lane20_strm0_data_valid    ( std__pe52__lane20_strm0_data_valid ),      
               .std__pe52__lane20_strm0_data_mask     ( std__pe52__lane20_strm0_data_mask  ),      

               .pe52__std__lane20_strm1_ready         ( pe52__std__lane20_strm1_ready      ),      
               .std__pe52__lane20_strm1_cntl          ( std__pe52__lane20_strm1_cntl       ),      
               .std__pe52__lane20_strm1_data          ( std__pe52__lane20_strm1_data       ),      
               .std__pe52__lane20_strm1_data_valid    ( std__pe52__lane20_strm1_data_valid ),      
               .std__pe52__lane20_strm1_data_mask     ( std__pe52__lane20_strm1_data_mask  ),      

               // PE 52, Lane 21                 
               .pe52__std__lane21_strm0_ready         ( pe52__std__lane21_strm0_ready      ),      
               .std__pe52__lane21_strm0_cntl          ( std__pe52__lane21_strm0_cntl       ),      
               .std__pe52__lane21_strm0_data          ( std__pe52__lane21_strm0_data       ),      
               .std__pe52__lane21_strm0_data_valid    ( std__pe52__lane21_strm0_data_valid ),      
               .std__pe52__lane21_strm0_data_mask     ( std__pe52__lane21_strm0_data_mask  ),      

               .pe52__std__lane21_strm1_ready         ( pe52__std__lane21_strm1_ready      ),      
               .std__pe52__lane21_strm1_cntl          ( std__pe52__lane21_strm1_cntl       ),      
               .std__pe52__lane21_strm1_data          ( std__pe52__lane21_strm1_data       ),      
               .std__pe52__lane21_strm1_data_valid    ( std__pe52__lane21_strm1_data_valid ),      
               .std__pe52__lane21_strm1_data_mask     ( std__pe52__lane21_strm1_data_mask  ),      

               // PE 52, Lane 22                 
               .pe52__std__lane22_strm0_ready         ( pe52__std__lane22_strm0_ready      ),      
               .std__pe52__lane22_strm0_cntl          ( std__pe52__lane22_strm0_cntl       ),      
               .std__pe52__lane22_strm0_data          ( std__pe52__lane22_strm0_data       ),      
               .std__pe52__lane22_strm0_data_valid    ( std__pe52__lane22_strm0_data_valid ),      
               .std__pe52__lane22_strm0_data_mask     ( std__pe52__lane22_strm0_data_mask  ),      

               .pe52__std__lane22_strm1_ready         ( pe52__std__lane22_strm1_ready      ),      
               .std__pe52__lane22_strm1_cntl          ( std__pe52__lane22_strm1_cntl       ),      
               .std__pe52__lane22_strm1_data          ( std__pe52__lane22_strm1_data       ),      
               .std__pe52__lane22_strm1_data_valid    ( std__pe52__lane22_strm1_data_valid ),      
               .std__pe52__lane22_strm1_data_mask     ( std__pe52__lane22_strm1_data_mask  ),      

               // PE 52, Lane 23                 
               .pe52__std__lane23_strm0_ready         ( pe52__std__lane23_strm0_ready      ),      
               .std__pe52__lane23_strm0_cntl          ( std__pe52__lane23_strm0_cntl       ),      
               .std__pe52__lane23_strm0_data          ( std__pe52__lane23_strm0_data       ),      
               .std__pe52__lane23_strm0_data_valid    ( std__pe52__lane23_strm0_data_valid ),      
               .std__pe52__lane23_strm0_data_mask     ( std__pe52__lane23_strm0_data_mask  ),      

               .pe52__std__lane23_strm1_ready         ( pe52__std__lane23_strm1_ready      ),      
               .std__pe52__lane23_strm1_cntl          ( std__pe52__lane23_strm1_cntl       ),      
               .std__pe52__lane23_strm1_data          ( std__pe52__lane23_strm1_data       ),      
               .std__pe52__lane23_strm1_data_valid    ( std__pe52__lane23_strm1_data_valid ),      
               .std__pe52__lane23_strm1_data_mask     ( std__pe52__lane23_strm1_data_mask  ),      

               // PE 52, Lane 24                 
               .pe52__std__lane24_strm0_ready         ( pe52__std__lane24_strm0_ready      ),      
               .std__pe52__lane24_strm0_cntl          ( std__pe52__lane24_strm0_cntl       ),      
               .std__pe52__lane24_strm0_data          ( std__pe52__lane24_strm0_data       ),      
               .std__pe52__lane24_strm0_data_valid    ( std__pe52__lane24_strm0_data_valid ),      
               .std__pe52__lane24_strm0_data_mask     ( std__pe52__lane24_strm0_data_mask  ),      

               .pe52__std__lane24_strm1_ready         ( pe52__std__lane24_strm1_ready      ),      
               .std__pe52__lane24_strm1_cntl          ( std__pe52__lane24_strm1_cntl       ),      
               .std__pe52__lane24_strm1_data          ( std__pe52__lane24_strm1_data       ),      
               .std__pe52__lane24_strm1_data_valid    ( std__pe52__lane24_strm1_data_valid ),      
               .std__pe52__lane24_strm1_data_mask     ( std__pe52__lane24_strm1_data_mask  ),      

               // PE 52, Lane 25                 
               .pe52__std__lane25_strm0_ready         ( pe52__std__lane25_strm0_ready      ),      
               .std__pe52__lane25_strm0_cntl          ( std__pe52__lane25_strm0_cntl       ),      
               .std__pe52__lane25_strm0_data          ( std__pe52__lane25_strm0_data       ),      
               .std__pe52__lane25_strm0_data_valid    ( std__pe52__lane25_strm0_data_valid ),      
               .std__pe52__lane25_strm0_data_mask     ( std__pe52__lane25_strm0_data_mask  ),      

               .pe52__std__lane25_strm1_ready         ( pe52__std__lane25_strm1_ready      ),      
               .std__pe52__lane25_strm1_cntl          ( std__pe52__lane25_strm1_cntl       ),      
               .std__pe52__lane25_strm1_data          ( std__pe52__lane25_strm1_data       ),      
               .std__pe52__lane25_strm1_data_valid    ( std__pe52__lane25_strm1_data_valid ),      
               .std__pe52__lane25_strm1_data_mask     ( std__pe52__lane25_strm1_data_mask  ),      

               // PE 52, Lane 26                 
               .pe52__std__lane26_strm0_ready         ( pe52__std__lane26_strm0_ready      ),      
               .std__pe52__lane26_strm0_cntl          ( std__pe52__lane26_strm0_cntl       ),      
               .std__pe52__lane26_strm0_data          ( std__pe52__lane26_strm0_data       ),      
               .std__pe52__lane26_strm0_data_valid    ( std__pe52__lane26_strm0_data_valid ),      
               .std__pe52__lane26_strm0_data_mask     ( std__pe52__lane26_strm0_data_mask  ),      

               .pe52__std__lane26_strm1_ready         ( pe52__std__lane26_strm1_ready      ),      
               .std__pe52__lane26_strm1_cntl          ( std__pe52__lane26_strm1_cntl       ),      
               .std__pe52__lane26_strm1_data          ( std__pe52__lane26_strm1_data       ),      
               .std__pe52__lane26_strm1_data_valid    ( std__pe52__lane26_strm1_data_valid ),      
               .std__pe52__lane26_strm1_data_mask     ( std__pe52__lane26_strm1_data_mask  ),      

               // PE 52, Lane 27                 
               .pe52__std__lane27_strm0_ready         ( pe52__std__lane27_strm0_ready      ),      
               .std__pe52__lane27_strm0_cntl          ( std__pe52__lane27_strm0_cntl       ),      
               .std__pe52__lane27_strm0_data          ( std__pe52__lane27_strm0_data       ),      
               .std__pe52__lane27_strm0_data_valid    ( std__pe52__lane27_strm0_data_valid ),      
               .std__pe52__lane27_strm0_data_mask     ( std__pe52__lane27_strm0_data_mask  ),      

               .pe52__std__lane27_strm1_ready         ( pe52__std__lane27_strm1_ready      ),      
               .std__pe52__lane27_strm1_cntl          ( std__pe52__lane27_strm1_cntl       ),      
               .std__pe52__lane27_strm1_data          ( std__pe52__lane27_strm1_data       ),      
               .std__pe52__lane27_strm1_data_valid    ( std__pe52__lane27_strm1_data_valid ),      
               .std__pe52__lane27_strm1_data_mask     ( std__pe52__lane27_strm1_data_mask  ),      

               // PE 52, Lane 28                 
               .pe52__std__lane28_strm0_ready         ( pe52__std__lane28_strm0_ready      ),      
               .std__pe52__lane28_strm0_cntl          ( std__pe52__lane28_strm0_cntl       ),      
               .std__pe52__lane28_strm0_data          ( std__pe52__lane28_strm0_data       ),      
               .std__pe52__lane28_strm0_data_valid    ( std__pe52__lane28_strm0_data_valid ),      
               .std__pe52__lane28_strm0_data_mask     ( std__pe52__lane28_strm0_data_mask  ),      

               .pe52__std__lane28_strm1_ready         ( pe52__std__lane28_strm1_ready      ),      
               .std__pe52__lane28_strm1_cntl          ( std__pe52__lane28_strm1_cntl       ),      
               .std__pe52__lane28_strm1_data          ( std__pe52__lane28_strm1_data       ),      
               .std__pe52__lane28_strm1_data_valid    ( std__pe52__lane28_strm1_data_valid ),      
               .std__pe52__lane28_strm1_data_mask     ( std__pe52__lane28_strm1_data_mask  ),      

               // PE 52, Lane 29                 
               .pe52__std__lane29_strm0_ready         ( pe52__std__lane29_strm0_ready      ),      
               .std__pe52__lane29_strm0_cntl          ( std__pe52__lane29_strm0_cntl       ),      
               .std__pe52__lane29_strm0_data          ( std__pe52__lane29_strm0_data       ),      
               .std__pe52__lane29_strm0_data_valid    ( std__pe52__lane29_strm0_data_valid ),      
               .std__pe52__lane29_strm0_data_mask     ( std__pe52__lane29_strm0_data_mask  ),      

               .pe52__std__lane29_strm1_ready         ( pe52__std__lane29_strm1_ready      ),      
               .std__pe52__lane29_strm1_cntl          ( std__pe52__lane29_strm1_cntl       ),      
               .std__pe52__lane29_strm1_data          ( std__pe52__lane29_strm1_data       ),      
               .std__pe52__lane29_strm1_data_valid    ( std__pe52__lane29_strm1_data_valid ),      
               .std__pe52__lane29_strm1_data_mask     ( std__pe52__lane29_strm1_data_mask  ),      

               // PE 52, Lane 30                 
               .pe52__std__lane30_strm0_ready         ( pe52__std__lane30_strm0_ready      ),      
               .std__pe52__lane30_strm0_cntl          ( std__pe52__lane30_strm0_cntl       ),      
               .std__pe52__lane30_strm0_data          ( std__pe52__lane30_strm0_data       ),      
               .std__pe52__lane30_strm0_data_valid    ( std__pe52__lane30_strm0_data_valid ),      
               .std__pe52__lane30_strm0_data_mask     ( std__pe52__lane30_strm0_data_mask  ),      

               .pe52__std__lane30_strm1_ready         ( pe52__std__lane30_strm1_ready      ),      
               .std__pe52__lane30_strm1_cntl          ( std__pe52__lane30_strm1_cntl       ),      
               .std__pe52__lane30_strm1_data          ( std__pe52__lane30_strm1_data       ),      
               .std__pe52__lane30_strm1_data_valid    ( std__pe52__lane30_strm1_data_valid ),      
               .std__pe52__lane30_strm1_data_mask     ( std__pe52__lane30_strm1_data_mask  ),      

               // PE 52, Lane 31                 
               .pe52__std__lane31_strm0_ready         ( pe52__std__lane31_strm0_ready      ),      
               .std__pe52__lane31_strm0_cntl          ( std__pe52__lane31_strm0_cntl       ),      
               .std__pe52__lane31_strm0_data          ( std__pe52__lane31_strm0_data       ),      
               .std__pe52__lane31_strm0_data_valid    ( std__pe52__lane31_strm0_data_valid ),      
               .std__pe52__lane31_strm0_data_mask     ( std__pe52__lane31_strm0_data_mask  ),      

               .pe52__std__lane31_strm1_ready         ( pe52__std__lane31_strm1_ready      ),      
               .std__pe52__lane31_strm1_cntl          ( std__pe52__lane31_strm1_cntl       ),      
               .std__pe52__lane31_strm1_data          ( std__pe52__lane31_strm1_data       ),      
               .std__pe52__lane31_strm1_data_valid    ( std__pe52__lane31_strm1_data_valid ),      
               .std__pe52__lane31_strm1_data_mask     ( std__pe52__lane31_strm1_data_mask  ),      

               // PE 53, Lane 0                 
               .pe53__std__lane0_strm0_ready         ( pe53__std__lane0_strm0_ready      ),      
               .std__pe53__lane0_strm0_cntl          ( std__pe53__lane0_strm0_cntl       ),      
               .std__pe53__lane0_strm0_data          ( std__pe53__lane0_strm0_data       ),      
               .std__pe53__lane0_strm0_data_valid    ( std__pe53__lane0_strm0_data_valid ),      
               .std__pe53__lane0_strm0_data_mask     ( std__pe53__lane0_strm0_data_mask  ),      

               .pe53__std__lane0_strm1_ready         ( pe53__std__lane0_strm1_ready      ),      
               .std__pe53__lane0_strm1_cntl          ( std__pe53__lane0_strm1_cntl       ),      
               .std__pe53__lane0_strm1_data          ( std__pe53__lane0_strm1_data       ),      
               .std__pe53__lane0_strm1_data_valid    ( std__pe53__lane0_strm1_data_valid ),      
               .std__pe53__lane0_strm1_data_mask     ( std__pe53__lane0_strm1_data_mask  ),      

               // PE 53, Lane 1                 
               .pe53__std__lane1_strm0_ready         ( pe53__std__lane1_strm0_ready      ),      
               .std__pe53__lane1_strm0_cntl          ( std__pe53__lane1_strm0_cntl       ),      
               .std__pe53__lane1_strm0_data          ( std__pe53__lane1_strm0_data       ),      
               .std__pe53__lane1_strm0_data_valid    ( std__pe53__lane1_strm0_data_valid ),      
               .std__pe53__lane1_strm0_data_mask     ( std__pe53__lane1_strm0_data_mask  ),      

               .pe53__std__lane1_strm1_ready         ( pe53__std__lane1_strm1_ready      ),      
               .std__pe53__lane1_strm1_cntl          ( std__pe53__lane1_strm1_cntl       ),      
               .std__pe53__lane1_strm1_data          ( std__pe53__lane1_strm1_data       ),      
               .std__pe53__lane1_strm1_data_valid    ( std__pe53__lane1_strm1_data_valid ),      
               .std__pe53__lane1_strm1_data_mask     ( std__pe53__lane1_strm1_data_mask  ),      

               // PE 53, Lane 2                 
               .pe53__std__lane2_strm0_ready         ( pe53__std__lane2_strm0_ready      ),      
               .std__pe53__lane2_strm0_cntl          ( std__pe53__lane2_strm0_cntl       ),      
               .std__pe53__lane2_strm0_data          ( std__pe53__lane2_strm0_data       ),      
               .std__pe53__lane2_strm0_data_valid    ( std__pe53__lane2_strm0_data_valid ),      
               .std__pe53__lane2_strm0_data_mask     ( std__pe53__lane2_strm0_data_mask  ),      

               .pe53__std__lane2_strm1_ready         ( pe53__std__lane2_strm1_ready      ),      
               .std__pe53__lane2_strm1_cntl          ( std__pe53__lane2_strm1_cntl       ),      
               .std__pe53__lane2_strm1_data          ( std__pe53__lane2_strm1_data       ),      
               .std__pe53__lane2_strm1_data_valid    ( std__pe53__lane2_strm1_data_valid ),      
               .std__pe53__lane2_strm1_data_mask     ( std__pe53__lane2_strm1_data_mask  ),      

               // PE 53, Lane 3                 
               .pe53__std__lane3_strm0_ready         ( pe53__std__lane3_strm0_ready      ),      
               .std__pe53__lane3_strm0_cntl          ( std__pe53__lane3_strm0_cntl       ),      
               .std__pe53__lane3_strm0_data          ( std__pe53__lane3_strm0_data       ),      
               .std__pe53__lane3_strm0_data_valid    ( std__pe53__lane3_strm0_data_valid ),      
               .std__pe53__lane3_strm0_data_mask     ( std__pe53__lane3_strm0_data_mask  ),      

               .pe53__std__lane3_strm1_ready         ( pe53__std__lane3_strm1_ready      ),      
               .std__pe53__lane3_strm1_cntl          ( std__pe53__lane3_strm1_cntl       ),      
               .std__pe53__lane3_strm1_data          ( std__pe53__lane3_strm1_data       ),      
               .std__pe53__lane3_strm1_data_valid    ( std__pe53__lane3_strm1_data_valid ),      
               .std__pe53__lane3_strm1_data_mask     ( std__pe53__lane3_strm1_data_mask  ),      

               // PE 53, Lane 4                 
               .pe53__std__lane4_strm0_ready         ( pe53__std__lane4_strm0_ready      ),      
               .std__pe53__lane4_strm0_cntl          ( std__pe53__lane4_strm0_cntl       ),      
               .std__pe53__lane4_strm0_data          ( std__pe53__lane4_strm0_data       ),      
               .std__pe53__lane4_strm0_data_valid    ( std__pe53__lane4_strm0_data_valid ),      
               .std__pe53__lane4_strm0_data_mask     ( std__pe53__lane4_strm0_data_mask  ),      

               .pe53__std__lane4_strm1_ready         ( pe53__std__lane4_strm1_ready      ),      
               .std__pe53__lane4_strm1_cntl          ( std__pe53__lane4_strm1_cntl       ),      
               .std__pe53__lane4_strm1_data          ( std__pe53__lane4_strm1_data       ),      
               .std__pe53__lane4_strm1_data_valid    ( std__pe53__lane4_strm1_data_valid ),      
               .std__pe53__lane4_strm1_data_mask     ( std__pe53__lane4_strm1_data_mask  ),      

               // PE 53, Lane 5                 
               .pe53__std__lane5_strm0_ready         ( pe53__std__lane5_strm0_ready      ),      
               .std__pe53__lane5_strm0_cntl          ( std__pe53__lane5_strm0_cntl       ),      
               .std__pe53__lane5_strm0_data          ( std__pe53__lane5_strm0_data       ),      
               .std__pe53__lane5_strm0_data_valid    ( std__pe53__lane5_strm0_data_valid ),      
               .std__pe53__lane5_strm0_data_mask     ( std__pe53__lane5_strm0_data_mask  ),      

               .pe53__std__lane5_strm1_ready         ( pe53__std__lane5_strm1_ready      ),      
               .std__pe53__lane5_strm1_cntl          ( std__pe53__lane5_strm1_cntl       ),      
               .std__pe53__lane5_strm1_data          ( std__pe53__lane5_strm1_data       ),      
               .std__pe53__lane5_strm1_data_valid    ( std__pe53__lane5_strm1_data_valid ),      
               .std__pe53__lane5_strm1_data_mask     ( std__pe53__lane5_strm1_data_mask  ),      

               // PE 53, Lane 6                 
               .pe53__std__lane6_strm0_ready         ( pe53__std__lane6_strm0_ready      ),      
               .std__pe53__lane6_strm0_cntl          ( std__pe53__lane6_strm0_cntl       ),      
               .std__pe53__lane6_strm0_data          ( std__pe53__lane6_strm0_data       ),      
               .std__pe53__lane6_strm0_data_valid    ( std__pe53__lane6_strm0_data_valid ),      
               .std__pe53__lane6_strm0_data_mask     ( std__pe53__lane6_strm0_data_mask  ),      

               .pe53__std__lane6_strm1_ready         ( pe53__std__lane6_strm1_ready      ),      
               .std__pe53__lane6_strm1_cntl          ( std__pe53__lane6_strm1_cntl       ),      
               .std__pe53__lane6_strm1_data          ( std__pe53__lane6_strm1_data       ),      
               .std__pe53__lane6_strm1_data_valid    ( std__pe53__lane6_strm1_data_valid ),      
               .std__pe53__lane6_strm1_data_mask     ( std__pe53__lane6_strm1_data_mask  ),      

               // PE 53, Lane 7                 
               .pe53__std__lane7_strm0_ready         ( pe53__std__lane7_strm0_ready      ),      
               .std__pe53__lane7_strm0_cntl          ( std__pe53__lane7_strm0_cntl       ),      
               .std__pe53__lane7_strm0_data          ( std__pe53__lane7_strm0_data       ),      
               .std__pe53__lane7_strm0_data_valid    ( std__pe53__lane7_strm0_data_valid ),      
               .std__pe53__lane7_strm0_data_mask     ( std__pe53__lane7_strm0_data_mask  ),      

               .pe53__std__lane7_strm1_ready         ( pe53__std__lane7_strm1_ready      ),      
               .std__pe53__lane7_strm1_cntl          ( std__pe53__lane7_strm1_cntl       ),      
               .std__pe53__lane7_strm1_data          ( std__pe53__lane7_strm1_data       ),      
               .std__pe53__lane7_strm1_data_valid    ( std__pe53__lane7_strm1_data_valid ),      
               .std__pe53__lane7_strm1_data_mask     ( std__pe53__lane7_strm1_data_mask  ),      

               // PE 53, Lane 8                 
               .pe53__std__lane8_strm0_ready         ( pe53__std__lane8_strm0_ready      ),      
               .std__pe53__lane8_strm0_cntl          ( std__pe53__lane8_strm0_cntl       ),      
               .std__pe53__lane8_strm0_data          ( std__pe53__lane8_strm0_data       ),      
               .std__pe53__lane8_strm0_data_valid    ( std__pe53__lane8_strm0_data_valid ),      
               .std__pe53__lane8_strm0_data_mask     ( std__pe53__lane8_strm0_data_mask  ),      

               .pe53__std__lane8_strm1_ready         ( pe53__std__lane8_strm1_ready      ),      
               .std__pe53__lane8_strm1_cntl          ( std__pe53__lane8_strm1_cntl       ),      
               .std__pe53__lane8_strm1_data          ( std__pe53__lane8_strm1_data       ),      
               .std__pe53__lane8_strm1_data_valid    ( std__pe53__lane8_strm1_data_valid ),      
               .std__pe53__lane8_strm1_data_mask     ( std__pe53__lane8_strm1_data_mask  ),      

               // PE 53, Lane 9                 
               .pe53__std__lane9_strm0_ready         ( pe53__std__lane9_strm0_ready      ),      
               .std__pe53__lane9_strm0_cntl          ( std__pe53__lane9_strm0_cntl       ),      
               .std__pe53__lane9_strm0_data          ( std__pe53__lane9_strm0_data       ),      
               .std__pe53__lane9_strm0_data_valid    ( std__pe53__lane9_strm0_data_valid ),      
               .std__pe53__lane9_strm0_data_mask     ( std__pe53__lane9_strm0_data_mask  ),      

               .pe53__std__lane9_strm1_ready         ( pe53__std__lane9_strm1_ready      ),      
               .std__pe53__lane9_strm1_cntl          ( std__pe53__lane9_strm1_cntl       ),      
               .std__pe53__lane9_strm1_data          ( std__pe53__lane9_strm1_data       ),      
               .std__pe53__lane9_strm1_data_valid    ( std__pe53__lane9_strm1_data_valid ),      
               .std__pe53__lane9_strm1_data_mask     ( std__pe53__lane9_strm1_data_mask  ),      

               // PE 53, Lane 10                 
               .pe53__std__lane10_strm0_ready         ( pe53__std__lane10_strm0_ready      ),      
               .std__pe53__lane10_strm0_cntl          ( std__pe53__lane10_strm0_cntl       ),      
               .std__pe53__lane10_strm0_data          ( std__pe53__lane10_strm0_data       ),      
               .std__pe53__lane10_strm0_data_valid    ( std__pe53__lane10_strm0_data_valid ),      
               .std__pe53__lane10_strm0_data_mask     ( std__pe53__lane10_strm0_data_mask  ),      

               .pe53__std__lane10_strm1_ready         ( pe53__std__lane10_strm1_ready      ),      
               .std__pe53__lane10_strm1_cntl          ( std__pe53__lane10_strm1_cntl       ),      
               .std__pe53__lane10_strm1_data          ( std__pe53__lane10_strm1_data       ),      
               .std__pe53__lane10_strm1_data_valid    ( std__pe53__lane10_strm1_data_valid ),      
               .std__pe53__lane10_strm1_data_mask     ( std__pe53__lane10_strm1_data_mask  ),      

               // PE 53, Lane 11                 
               .pe53__std__lane11_strm0_ready         ( pe53__std__lane11_strm0_ready      ),      
               .std__pe53__lane11_strm0_cntl          ( std__pe53__lane11_strm0_cntl       ),      
               .std__pe53__lane11_strm0_data          ( std__pe53__lane11_strm0_data       ),      
               .std__pe53__lane11_strm0_data_valid    ( std__pe53__lane11_strm0_data_valid ),      
               .std__pe53__lane11_strm0_data_mask     ( std__pe53__lane11_strm0_data_mask  ),      

               .pe53__std__lane11_strm1_ready         ( pe53__std__lane11_strm1_ready      ),      
               .std__pe53__lane11_strm1_cntl          ( std__pe53__lane11_strm1_cntl       ),      
               .std__pe53__lane11_strm1_data          ( std__pe53__lane11_strm1_data       ),      
               .std__pe53__lane11_strm1_data_valid    ( std__pe53__lane11_strm1_data_valid ),      
               .std__pe53__lane11_strm1_data_mask     ( std__pe53__lane11_strm1_data_mask  ),      

               // PE 53, Lane 12                 
               .pe53__std__lane12_strm0_ready         ( pe53__std__lane12_strm0_ready      ),      
               .std__pe53__lane12_strm0_cntl          ( std__pe53__lane12_strm0_cntl       ),      
               .std__pe53__lane12_strm0_data          ( std__pe53__lane12_strm0_data       ),      
               .std__pe53__lane12_strm0_data_valid    ( std__pe53__lane12_strm0_data_valid ),      
               .std__pe53__lane12_strm0_data_mask     ( std__pe53__lane12_strm0_data_mask  ),      

               .pe53__std__lane12_strm1_ready         ( pe53__std__lane12_strm1_ready      ),      
               .std__pe53__lane12_strm1_cntl          ( std__pe53__lane12_strm1_cntl       ),      
               .std__pe53__lane12_strm1_data          ( std__pe53__lane12_strm1_data       ),      
               .std__pe53__lane12_strm1_data_valid    ( std__pe53__lane12_strm1_data_valid ),      
               .std__pe53__lane12_strm1_data_mask     ( std__pe53__lane12_strm1_data_mask  ),      

               // PE 53, Lane 13                 
               .pe53__std__lane13_strm0_ready         ( pe53__std__lane13_strm0_ready      ),      
               .std__pe53__lane13_strm0_cntl          ( std__pe53__lane13_strm0_cntl       ),      
               .std__pe53__lane13_strm0_data          ( std__pe53__lane13_strm0_data       ),      
               .std__pe53__lane13_strm0_data_valid    ( std__pe53__lane13_strm0_data_valid ),      
               .std__pe53__lane13_strm0_data_mask     ( std__pe53__lane13_strm0_data_mask  ),      

               .pe53__std__lane13_strm1_ready         ( pe53__std__lane13_strm1_ready      ),      
               .std__pe53__lane13_strm1_cntl          ( std__pe53__lane13_strm1_cntl       ),      
               .std__pe53__lane13_strm1_data          ( std__pe53__lane13_strm1_data       ),      
               .std__pe53__lane13_strm1_data_valid    ( std__pe53__lane13_strm1_data_valid ),      
               .std__pe53__lane13_strm1_data_mask     ( std__pe53__lane13_strm1_data_mask  ),      

               // PE 53, Lane 14                 
               .pe53__std__lane14_strm0_ready         ( pe53__std__lane14_strm0_ready      ),      
               .std__pe53__lane14_strm0_cntl          ( std__pe53__lane14_strm0_cntl       ),      
               .std__pe53__lane14_strm0_data          ( std__pe53__lane14_strm0_data       ),      
               .std__pe53__lane14_strm0_data_valid    ( std__pe53__lane14_strm0_data_valid ),      
               .std__pe53__lane14_strm0_data_mask     ( std__pe53__lane14_strm0_data_mask  ),      

               .pe53__std__lane14_strm1_ready         ( pe53__std__lane14_strm1_ready      ),      
               .std__pe53__lane14_strm1_cntl          ( std__pe53__lane14_strm1_cntl       ),      
               .std__pe53__lane14_strm1_data          ( std__pe53__lane14_strm1_data       ),      
               .std__pe53__lane14_strm1_data_valid    ( std__pe53__lane14_strm1_data_valid ),      
               .std__pe53__lane14_strm1_data_mask     ( std__pe53__lane14_strm1_data_mask  ),      

               // PE 53, Lane 15                 
               .pe53__std__lane15_strm0_ready         ( pe53__std__lane15_strm0_ready      ),      
               .std__pe53__lane15_strm0_cntl          ( std__pe53__lane15_strm0_cntl       ),      
               .std__pe53__lane15_strm0_data          ( std__pe53__lane15_strm0_data       ),      
               .std__pe53__lane15_strm0_data_valid    ( std__pe53__lane15_strm0_data_valid ),      
               .std__pe53__lane15_strm0_data_mask     ( std__pe53__lane15_strm0_data_mask  ),      

               .pe53__std__lane15_strm1_ready         ( pe53__std__lane15_strm1_ready      ),      
               .std__pe53__lane15_strm1_cntl          ( std__pe53__lane15_strm1_cntl       ),      
               .std__pe53__lane15_strm1_data          ( std__pe53__lane15_strm1_data       ),      
               .std__pe53__lane15_strm1_data_valid    ( std__pe53__lane15_strm1_data_valid ),      
               .std__pe53__lane15_strm1_data_mask     ( std__pe53__lane15_strm1_data_mask  ),      

               // PE 53, Lane 16                 
               .pe53__std__lane16_strm0_ready         ( pe53__std__lane16_strm0_ready      ),      
               .std__pe53__lane16_strm0_cntl          ( std__pe53__lane16_strm0_cntl       ),      
               .std__pe53__lane16_strm0_data          ( std__pe53__lane16_strm0_data       ),      
               .std__pe53__lane16_strm0_data_valid    ( std__pe53__lane16_strm0_data_valid ),      
               .std__pe53__lane16_strm0_data_mask     ( std__pe53__lane16_strm0_data_mask  ),      

               .pe53__std__lane16_strm1_ready         ( pe53__std__lane16_strm1_ready      ),      
               .std__pe53__lane16_strm1_cntl          ( std__pe53__lane16_strm1_cntl       ),      
               .std__pe53__lane16_strm1_data          ( std__pe53__lane16_strm1_data       ),      
               .std__pe53__lane16_strm1_data_valid    ( std__pe53__lane16_strm1_data_valid ),      
               .std__pe53__lane16_strm1_data_mask     ( std__pe53__lane16_strm1_data_mask  ),      

               // PE 53, Lane 17                 
               .pe53__std__lane17_strm0_ready         ( pe53__std__lane17_strm0_ready      ),      
               .std__pe53__lane17_strm0_cntl          ( std__pe53__lane17_strm0_cntl       ),      
               .std__pe53__lane17_strm0_data          ( std__pe53__lane17_strm0_data       ),      
               .std__pe53__lane17_strm0_data_valid    ( std__pe53__lane17_strm0_data_valid ),      
               .std__pe53__lane17_strm0_data_mask     ( std__pe53__lane17_strm0_data_mask  ),      

               .pe53__std__lane17_strm1_ready         ( pe53__std__lane17_strm1_ready      ),      
               .std__pe53__lane17_strm1_cntl          ( std__pe53__lane17_strm1_cntl       ),      
               .std__pe53__lane17_strm1_data          ( std__pe53__lane17_strm1_data       ),      
               .std__pe53__lane17_strm1_data_valid    ( std__pe53__lane17_strm1_data_valid ),      
               .std__pe53__lane17_strm1_data_mask     ( std__pe53__lane17_strm1_data_mask  ),      

               // PE 53, Lane 18                 
               .pe53__std__lane18_strm0_ready         ( pe53__std__lane18_strm0_ready      ),      
               .std__pe53__lane18_strm0_cntl          ( std__pe53__lane18_strm0_cntl       ),      
               .std__pe53__lane18_strm0_data          ( std__pe53__lane18_strm0_data       ),      
               .std__pe53__lane18_strm0_data_valid    ( std__pe53__lane18_strm0_data_valid ),      
               .std__pe53__lane18_strm0_data_mask     ( std__pe53__lane18_strm0_data_mask  ),      

               .pe53__std__lane18_strm1_ready         ( pe53__std__lane18_strm1_ready      ),      
               .std__pe53__lane18_strm1_cntl          ( std__pe53__lane18_strm1_cntl       ),      
               .std__pe53__lane18_strm1_data          ( std__pe53__lane18_strm1_data       ),      
               .std__pe53__lane18_strm1_data_valid    ( std__pe53__lane18_strm1_data_valid ),      
               .std__pe53__lane18_strm1_data_mask     ( std__pe53__lane18_strm1_data_mask  ),      

               // PE 53, Lane 19                 
               .pe53__std__lane19_strm0_ready         ( pe53__std__lane19_strm0_ready      ),      
               .std__pe53__lane19_strm0_cntl          ( std__pe53__lane19_strm0_cntl       ),      
               .std__pe53__lane19_strm0_data          ( std__pe53__lane19_strm0_data       ),      
               .std__pe53__lane19_strm0_data_valid    ( std__pe53__lane19_strm0_data_valid ),      
               .std__pe53__lane19_strm0_data_mask     ( std__pe53__lane19_strm0_data_mask  ),      

               .pe53__std__lane19_strm1_ready         ( pe53__std__lane19_strm1_ready      ),      
               .std__pe53__lane19_strm1_cntl          ( std__pe53__lane19_strm1_cntl       ),      
               .std__pe53__lane19_strm1_data          ( std__pe53__lane19_strm1_data       ),      
               .std__pe53__lane19_strm1_data_valid    ( std__pe53__lane19_strm1_data_valid ),      
               .std__pe53__lane19_strm1_data_mask     ( std__pe53__lane19_strm1_data_mask  ),      

               // PE 53, Lane 20                 
               .pe53__std__lane20_strm0_ready         ( pe53__std__lane20_strm0_ready      ),      
               .std__pe53__lane20_strm0_cntl          ( std__pe53__lane20_strm0_cntl       ),      
               .std__pe53__lane20_strm0_data          ( std__pe53__lane20_strm0_data       ),      
               .std__pe53__lane20_strm0_data_valid    ( std__pe53__lane20_strm0_data_valid ),      
               .std__pe53__lane20_strm0_data_mask     ( std__pe53__lane20_strm0_data_mask  ),      

               .pe53__std__lane20_strm1_ready         ( pe53__std__lane20_strm1_ready      ),      
               .std__pe53__lane20_strm1_cntl          ( std__pe53__lane20_strm1_cntl       ),      
               .std__pe53__lane20_strm1_data          ( std__pe53__lane20_strm1_data       ),      
               .std__pe53__lane20_strm1_data_valid    ( std__pe53__lane20_strm1_data_valid ),      
               .std__pe53__lane20_strm1_data_mask     ( std__pe53__lane20_strm1_data_mask  ),      

               // PE 53, Lane 21                 
               .pe53__std__lane21_strm0_ready         ( pe53__std__lane21_strm0_ready      ),      
               .std__pe53__lane21_strm0_cntl          ( std__pe53__lane21_strm0_cntl       ),      
               .std__pe53__lane21_strm0_data          ( std__pe53__lane21_strm0_data       ),      
               .std__pe53__lane21_strm0_data_valid    ( std__pe53__lane21_strm0_data_valid ),      
               .std__pe53__lane21_strm0_data_mask     ( std__pe53__lane21_strm0_data_mask  ),      

               .pe53__std__lane21_strm1_ready         ( pe53__std__lane21_strm1_ready      ),      
               .std__pe53__lane21_strm1_cntl          ( std__pe53__lane21_strm1_cntl       ),      
               .std__pe53__lane21_strm1_data          ( std__pe53__lane21_strm1_data       ),      
               .std__pe53__lane21_strm1_data_valid    ( std__pe53__lane21_strm1_data_valid ),      
               .std__pe53__lane21_strm1_data_mask     ( std__pe53__lane21_strm1_data_mask  ),      

               // PE 53, Lane 22                 
               .pe53__std__lane22_strm0_ready         ( pe53__std__lane22_strm0_ready      ),      
               .std__pe53__lane22_strm0_cntl          ( std__pe53__lane22_strm0_cntl       ),      
               .std__pe53__lane22_strm0_data          ( std__pe53__lane22_strm0_data       ),      
               .std__pe53__lane22_strm0_data_valid    ( std__pe53__lane22_strm0_data_valid ),      
               .std__pe53__lane22_strm0_data_mask     ( std__pe53__lane22_strm0_data_mask  ),      

               .pe53__std__lane22_strm1_ready         ( pe53__std__lane22_strm1_ready      ),      
               .std__pe53__lane22_strm1_cntl          ( std__pe53__lane22_strm1_cntl       ),      
               .std__pe53__lane22_strm1_data          ( std__pe53__lane22_strm1_data       ),      
               .std__pe53__lane22_strm1_data_valid    ( std__pe53__lane22_strm1_data_valid ),      
               .std__pe53__lane22_strm1_data_mask     ( std__pe53__lane22_strm1_data_mask  ),      

               // PE 53, Lane 23                 
               .pe53__std__lane23_strm0_ready         ( pe53__std__lane23_strm0_ready      ),      
               .std__pe53__lane23_strm0_cntl          ( std__pe53__lane23_strm0_cntl       ),      
               .std__pe53__lane23_strm0_data          ( std__pe53__lane23_strm0_data       ),      
               .std__pe53__lane23_strm0_data_valid    ( std__pe53__lane23_strm0_data_valid ),      
               .std__pe53__lane23_strm0_data_mask     ( std__pe53__lane23_strm0_data_mask  ),      

               .pe53__std__lane23_strm1_ready         ( pe53__std__lane23_strm1_ready      ),      
               .std__pe53__lane23_strm1_cntl          ( std__pe53__lane23_strm1_cntl       ),      
               .std__pe53__lane23_strm1_data          ( std__pe53__lane23_strm1_data       ),      
               .std__pe53__lane23_strm1_data_valid    ( std__pe53__lane23_strm1_data_valid ),      
               .std__pe53__lane23_strm1_data_mask     ( std__pe53__lane23_strm1_data_mask  ),      

               // PE 53, Lane 24                 
               .pe53__std__lane24_strm0_ready         ( pe53__std__lane24_strm0_ready      ),      
               .std__pe53__lane24_strm0_cntl          ( std__pe53__lane24_strm0_cntl       ),      
               .std__pe53__lane24_strm0_data          ( std__pe53__lane24_strm0_data       ),      
               .std__pe53__lane24_strm0_data_valid    ( std__pe53__lane24_strm0_data_valid ),      
               .std__pe53__lane24_strm0_data_mask     ( std__pe53__lane24_strm0_data_mask  ),      

               .pe53__std__lane24_strm1_ready         ( pe53__std__lane24_strm1_ready      ),      
               .std__pe53__lane24_strm1_cntl          ( std__pe53__lane24_strm1_cntl       ),      
               .std__pe53__lane24_strm1_data          ( std__pe53__lane24_strm1_data       ),      
               .std__pe53__lane24_strm1_data_valid    ( std__pe53__lane24_strm1_data_valid ),      
               .std__pe53__lane24_strm1_data_mask     ( std__pe53__lane24_strm1_data_mask  ),      

               // PE 53, Lane 25                 
               .pe53__std__lane25_strm0_ready         ( pe53__std__lane25_strm0_ready      ),      
               .std__pe53__lane25_strm0_cntl          ( std__pe53__lane25_strm0_cntl       ),      
               .std__pe53__lane25_strm0_data          ( std__pe53__lane25_strm0_data       ),      
               .std__pe53__lane25_strm0_data_valid    ( std__pe53__lane25_strm0_data_valid ),      
               .std__pe53__lane25_strm0_data_mask     ( std__pe53__lane25_strm0_data_mask  ),      

               .pe53__std__lane25_strm1_ready         ( pe53__std__lane25_strm1_ready      ),      
               .std__pe53__lane25_strm1_cntl          ( std__pe53__lane25_strm1_cntl       ),      
               .std__pe53__lane25_strm1_data          ( std__pe53__lane25_strm1_data       ),      
               .std__pe53__lane25_strm1_data_valid    ( std__pe53__lane25_strm1_data_valid ),      
               .std__pe53__lane25_strm1_data_mask     ( std__pe53__lane25_strm1_data_mask  ),      

               // PE 53, Lane 26                 
               .pe53__std__lane26_strm0_ready         ( pe53__std__lane26_strm0_ready      ),      
               .std__pe53__lane26_strm0_cntl          ( std__pe53__lane26_strm0_cntl       ),      
               .std__pe53__lane26_strm0_data          ( std__pe53__lane26_strm0_data       ),      
               .std__pe53__lane26_strm0_data_valid    ( std__pe53__lane26_strm0_data_valid ),      
               .std__pe53__lane26_strm0_data_mask     ( std__pe53__lane26_strm0_data_mask  ),      

               .pe53__std__lane26_strm1_ready         ( pe53__std__lane26_strm1_ready      ),      
               .std__pe53__lane26_strm1_cntl          ( std__pe53__lane26_strm1_cntl       ),      
               .std__pe53__lane26_strm1_data          ( std__pe53__lane26_strm1_data       ),      
               .std__pe53__lane26_strm1_data_valid    ( std__pe53__lane26_strm1_data_valid ),      
               .std__pe53__lane26_strm1_data_mask     ( std__pe53__lane26_strm1_data_mask  ),      

               // PE 53, Lane 27                 
               .pe53__std__lane27_strm0_ready         ( pe53__std__lane27_strm0_ready      ),      
               .std__pe53__lane27_strm0_cntl          ( std__pe53__lane27_strm0_cntl       ),      
               .std__pe53__lane27_strm0_data          ( std__pe53__lane27_strm0_data       ),      
               .std__pe53__lane27_strm0_data_valid    ( std__pe53__lane27_strm0_data_valid ),      
               .std__pe53__lane27_strm0_data_mask     ( std__pe53__lane27_strm0_data_mask  ),      

               .pe53__std__lane27_strm1_ready         ( pe53__std__lane27_strm1_ready      ),      
               .std__pe53__lane27_strm1_cntl          ( std__pe53__lane27_strm1_cntl       ),      
               .std__pe53__lane27_strm1_data          ( std__pe53__lane27_strm1_data       ),      
               .std__pe53__lane27_strm1_data_valid    ( std__pe53__lane27_strm1_data_valid ),      
               .std__pe53__lane27_strm1_data_mask     ( std__pe53__lane27_strm1_data_mask  ),      

               // PE 53, Lane 28                 
               .pe53__std__lane28_strm0_ready         ( pe53__std__lane28_strm0_ready      ),      
               .std__pe53__lane28_strm0_cntl          ( std__pe53__lane28_strm0_cntl       ),      
               .std__pe53__lane28_strm0_data          ( std__pe53__lane28_strm0_data       ),      
               .std__pe53__lane28_strm0_data_valid    ( std__pe53__lane28_strm0_data_valid ),      
               .std__pe53__lane28_strm0_data_mask     ( std__pe53__lane28_strm0_data_mask  ),      

               .pe53__std__lane28_strm1_ready         ( pe53__std__lane28_strm1_ready      ),      
               .std__pe53__lane28_strm1_cntl          ( std__pe53__lane28_strm1_cntl       ),      
               .std__pe53__lane28_strm1_data          ( std__pe53__lane28_strm1_data       ),      
               .std__pe53__lane28_strm1_data_valid    ( std__pe53__lane28_strm1_data_valid ),      
               .std__pe53__lane28_strm1_data_mask     ( std__pe53__lane28_strm1_data_mask  ),      

               // PE 53, Lane 29                 
               .pe53__std__lane29_strm0_ready         ( pe53__std__lane29_strm0_ready      ),      
               .std__pe53__lane29_strm0_cntl          ( std__pe53__lane29_strm0_cntl       ),      
               .std__pe53__lane29_strm0_data          ( std__pe53__lane29_strm0_data       ),      
               .std__pe53__lane29_strm0_data_valid    ( std__pe53__lane29_strm0_data_valid ),      
               .std__pe53__lane29_strm0_data_mask     ( std__pe53__lane29_strm0_data_mask  ),      

               .pe53__std__lane29_strm1_ready         ( pe53__std__lane29_strm1_ready      ),      
               .std__pe53__lane29_strm1_cntl          ( std__pe53__lane29_strm1_cntl       ),      
               .std__pe53__lane29_strm1_data          ( std__pe53__lane29_strm1_data       ),      
               .std__pe53__lane29_strm1_data_valid    ( std__pe53__lane29_strm1_data_valid ),      
               .std__pe53__lane29_strm1_data_mask     ( std__pe53__lane29_strm1_data_mask  ),      

               // PE 53, Lane 30                 
               .pe53__std__lane30_strm0_ready         ( pe53__std__lane30_strm0_ready      ),      
               .std__pe53__lane30_strm0_cntl          ( std__pe53__lane30_strm0_cntl       ),      
               .std__pe53__lane30_strm0_data          ( std__pe53__lane30_strm0_data       ),      
               .std__pe53__lane30_strm0_data_valid    ( std__pe53__lane30_strm0_data_valid ),      
               .std__pe53__lane30_strm0_data_mask     ( std__pe53__lane30_strm0_data_mask  ),      

               .pe53__std__lane30_strm1_ready         ( pe53__std__lane30_strm1_ready      ),      
               .std__pe53__lane30_strm1_cntl          ( std__pe53__lane30_strm1_cntl       ),      
               .std__pe53__lane30_strm1_data          ( std__pe53__lane30_strm1_data       ),      
               .std__pe53__lane30_strm1_data_valid    ( std__pe53__lane30_strm1_data_valid ),      
               .std__pe53__lane30_strm1_data_mask     ( std__pe53__lane30_strm1_data_mask  ),      

               // PE 53, Lane 31                 
               .pe53__std__lane31_strm0_ready         ( pe53__std__lane31_strm0_ready      ),      
               .std__pe53__lane31_strm0_cntl          ( std__pe53__lane31_strm0_cntl       ),      
               .std__pe53__lane31_strm0_data          ( std__pe53__lane31_strm0_data       ),      
               .std__pe53__lane31_strm0_data_valid    ( std__pe53__lane31_strm0_data_valid ),      
               .std__pe53__lane31_strm0_data_mask     ( std__pe53__lane31_strm0_data_mask  ),      

               .pe53__std__lane31_strm1_ready         ( pe53__std__lane31_strm1_ready      ),      
               .std__pe53__lane31_strm1_cntl          ( std__pe53__lane31_strm1_cntl       ),      
               .std__pe53__lane31_strm1_data          ( std__pe53__lane31_strm1_data       ),      
               .std__pe53__lane31_strm1_data_valid    ( std__pe53__lane31_strm1_data_valid ),      
               .std__pe53__lane31_strm1_data_mask     ( std__pe53__lane31_strm1_data_mask  ),      

               // PE 54, Lane 0                 
               .pe54__std__lane0_strm0_ready         ( pe54__std__lane0_strm0_ready      ),      
               .std__pe54__lane0_strm0_cntl          ( std__pe54__lane0_strm0_cntl       ),      
               .std__pe54__lane0_strm0_data          ( std__pe54__lane0_strm0_data       ),      
               .std__pe54__lane0_strm0_data_valid    ( std__pe54__lane0_strm0_data_valid ),      
               .std__pe54__lane0_strm0_data_mask     ( std__pe54__lane0_strm0_data_mask  ),      

               .pe54__std__lane0_strm1_ready         ( pe54__std__lane0_strm1_ready      ),      
               .std__pe54__lane0_strm1_cntl          ( std__pe54__lane0_strm1_cntl       ),      
               .std__pe54__lane0_strm1_data          ( std__pe54__lane0_strm1_data       ),      
               .std__pe54__lane0_strm1_data_valid    ( std__pe54__lane0_strm1_data_valid ),      
               .std__pe54__lane0_strm1_data_mask     ( std__pe54__lane0_strm1_data_mask  ),      

               // PE 54, Lane 1                 
               .pe54__std__lane1_strm0_ready         ( pe54__std__lane1_strm0_ready      ),      
               .std__pe54__lane1_strm0_cntl          ( std__pe54__lane1_strm0_cntl       ),      
               .std__pe54__lane1_strm0_data          ( std__pe54__lane1_strm0_data       ),      
               .std__pe54__lane1_strm0_data_valid    ( std__pe54__lane1_strm0_data_valid ),      
               .std__pe54__lane1_strm0_data_mask     ( std__pe54__lane1_strm0_data_mask  ),      

               .pe54__std__lane1_strm1_ready         ( pe54__std__lane1_strm1_ready      ),      
               .std__pe54__lane1_strm1_cntl          ( std__pe54__lane1_strm1_cntl       ),      
               .std__pe54__lane1_strm1_data          ( std__pe54__lane1_strm1_data       ),      
               .std__pe54__lane1_strm1_data_valid    ( std__pe54__lane1_strm1_data_valid ),      
               .std__pe54__lane1_strm1_data_mask     ( std__pe54__lane1_strm1_data_mask  ),      

               // PE 54, Lane 2                 
               .pe54__std__lane2_strm0_ready         ( pe54__std__lane2_strm0_ready      ),      
               .std__pe54__lane2_strm0_cntl          ( std__pe54__lane2_strm0_cntl       ),      
               .std__pe54__lane2_strm0_data          ( std__pe54__lane2_strm0_data       ),      
               .std__pe54__lane2_strm0_data_valid    ( std__pe54__lane2_strm0_data_valid ),      
               .std__pe54__lane2_strm0_data_mask     ( std__pe54__lane2_strm0_data_mask  ),      

               .pe54__std__lane2_strm1_ready         ( pe54__std__lane2_strm1_ready      ),      
               .std__pe54__lane2_strm1_cntl          ( std__pe54__lane2_strm1_cntl       ),      
               .std__pe54__lane2_strm1_data          ( std__pe54__lane2_strm1_data       ),      
               .std__pe54__lane2_strm1_data_valid    ( std__pe54__lane2_strm1_data_valid ),      
               .std__pe54__lane2_strm1_data_mask     ( std__pe54__lane2_strm1_data_mask  ),      

               // PE 54, Lane 3                 
               .pe54__std__lane3_strm0_ready         ( pe54__std__lane3_strm0_ready      ),      
               .std__pe54__lane3_strm0_cntl          ( std__pe54__lane3_strm0_cntl       ),      
               .std__pe54__lane3_strm0_data          ( std__pe54__lane3_strm0_data       ),      
               .std__pe54__lane3_strm0_data_valid    ( std__pe54__lane3_strm0_data_valid ),      
               .std__pe54__lane3_strm0_data_mask     ( std__pe54__lane3_strm0_data_mask  ),      

               .pe54__std__lane3_strm1_ready         ( pe54__std__lane3_strm1_ready      ),      
               .std__pe54__lane3_strm1_cntl          ( std__pe54__lane3_strm1_cntl       ),      
               .std__pe54__lane3_strm1_data          ( std__pe54__lane3_strm1_data       ),      
               .std__pe54__lane3_strm1_data_valid    ( std__pe54__lane3_strm1_data_valid ),      
               .std__pe54__lane3_strm1_data_mask     ( std__pe54__lane3_strm1_data_mask  ),      

               // PE 54, Lane 4                 
               .pe54__std__lane4_strm0_ready         ( pe54__std__lane4_strm0_ready      ),      
               .std__pe54__lane4_strm0_cntl          ( std__pe54__lane4_strm0_cntl       ),      
               .std__pe54__lane4_strm0_data          ( std__pe54__lane4_strm0_data       ),      
               .std__pe54__lane4_strm0_data_valid    ( std__pe54__lane4_strm0_data_valid ),      
               .std__pe54__lane4_strm0_data_mask     ( std__pe54__lane4_strm0_data_mask  ),      

               .pe54__std__lane4_strm1_ready         ( pe54__std__lane4_strm1_ready      ),      
               .std__pe54__lane4_strm1_cntl          ( std__pe54__lane4_strm1_cntl       ),      
               .std__pe54__lane4_strm1_data          ( std__pe54__lane4_strm1_data       ),      
               .std__pe54__lane4_strm1_data_valid    ( std__pe54__lane4_strm1_data_valid ),      
               .std__pe54__lane4_strm1_data_mask     ( std__pe54__lane4_strm1_data_mask  ),      

               // PE 54, Lane 5                 
               .pe54__std__lane5_strm0_ready         ( pe54__std__lane5_strm0_ready      ),      
               .std__pe54__lane5_strm0_cntl          ( std__pe54__lane5_strm0_cntl       ),      
               .std__pe54__lane5_strm0_data          ( std__pe54__lane5_strm0_data       ),      
               .std__pe54__lane5_strm0_data_valid    ( std__pe54__lane5_strm0_data_valid ),      
               .std__pe54__lane5_strm0_data_mask     ( std__pe54__lane5_strm0_data_mask  ),      

               .pe54__std__lane5_strm1_ready         ( pe54__std__lane5_strm1_ready      ),      
               .std__pe54__lane5_strm1_cntl          ( std__pe54__lane5_strm1_cntl       ),      
               .std__pe54__lane5_strm1_data          ( std__pe54__lane5_strm1_data       ),      
               .std__pe54__lane5_strm1_data_valid    ( std__pe54__lane5_strm1_data_valid ),      
               .std__pe54__lane5_strm1_data_mask     ( std__pe54__lane5_strm1_data_mask  ),      

               // PE 54, Lane 6                 
               .pe54__std__lane6_strm0_ready         ( pe54__std__lane6_strm0_ready      ),      
               .std__pe54__lane6_strm0_cntl          ( std__pe54__lane6_strm0_cntl       ),      
               .std__pe54__lane6_strm0_data          ( std__pe54__lane6_strm0_data       ),      
               .std__pe54__lane6_strm0_data_valid    ( std__pe54__lane6_strm0_data_valid ),      
               .std__pe54__lane6_strm0_data_mask     ( std__pe54__lane6_strm0_data_mask  ),      

               .pe54__std__lane6_strm1_ready         ( pe54__std__lane6_strm1_ready      ),      
               .std__pe54__lane6_strm1_cntl          ( std__pe54__lane6_strm1_cntl       ),      
               .std__pe54__lane6_strm1_data          ( std__pe54__lane6_strm1_data       ),      
               .std__pe54__lane6_strm1_data_valid    ( std__pe54__lane6_strm1_data_valid ),      
               .std__pe54__lane6_strm1_data_mask     ( std__pe54__lane6_strm1_data_mask  ),      

               // PE 54, Lane 7                 
               .pe54__std__lane7_strm0_ready         ( pe54__std__lane7_strm0_ready      ),      
               .std__pe54__lane7_strm0_cntl          ( std__pe54__lane7_strm0_cntl       ),      
               .std__pe54__lane7_strm0_data          ( std__pe54__lane7_strm0_data       ),      
               .std__pe54__lane7_strm0_data_valid    ( std__pe54__lane7_strm0_data_valid ),      
               .std__pe54__lane7_strm0_data_mask     ( std__pe54__lane7_strm0_data_mask  ),      

               .pe54__std__lane7_strm1_ready         ( pe54__std__lane7_strm1_ready      ),      
               .std__pe54__lane7_strm1_cntl          ( std__pe54__lane7_strm1_cntl       ),      
               .std__pe54__lane7_strm1_data          ( std__pe54__lane7_strm1_data       ),      
               .std__pe54__lane7_strm1_data_valid    ( std__pe54__lane7_strm1_data_valid ),      
               .std__pe54__lane7_strm1_data_mask     ( std__pe54__lane7_strm1_data_mask  ),      

               // PE 54, Lane 8                 
               .pe54__std__lane8_strm0_ready         ( pe54__std__lane8_strm0_ready      ),      
               .std__pe54__lane8_strm0_cntl          ( std__pe54__lane8_strm0_cntl       ),      
               .std__pe54__lane8_strm0_data          ( std__pe54__lane8_strm0_data       ),      
               .std__pe54__lane8_strm0_data_valid    ( std__pe54__lane8_strm0_data_valid ),      
               .std__pe54__lane8_strm0_data_mask     ( std__pe54__lane8_strm0_data_mask  ),      

               .pe54__std__lane8_strm1_ready         ( pe54__std__lane8_strm1_ready      ),      
               .std__pe54__lane8_strm1_cntl          ( std__pe54__lane8_strm1_cntl       ),      
               .std__pe54__lane8_strm1_data          ( std__pe54__lane8_strm1_data       ),      
               .std__pe54__lane8_strm1_data_valid    ( std__pe54__lane8_strm1_data_valid ),      
               .std__pe54__lane8_strm1_data_mask     ( std__pe54__lane8_strm1_data_mask  ),      

               // PE 54, Lane 9                 
               .pe54__std__lane9_strm0_ready         ( pe54__std__lane9_strm0_ready      ),      
               .std__pe54__lane9_strm0_cntl          ( std__pe54__lane9_strm0_cntl       ),      
               .std__pe54__lane9_strm0_data          ( std__pe54__lane9_strm0_data       ),      
               .std__pe54__lane9_strm0_data_valid    ( std__pe54__lane9_strm0_data_valid ),      
               .std__pe54__lane9_strm0_data_mask     ( std__pe54__lane9_strm0_data_mask  ),      

               .pe54__std__lane9_strm1_ready         ( pe54__std__lane9_strm1_ready      ),      
               .std__pe54__lane9_strm1_cntl          ( std__pe54__lane9_strm1_cntl       ),      
               .std__pe54__lane9_strm1_data          ( std__pe54__lane9_strm1_data       ),      
               .std__pe54__lane9_strm1_data_valid    ( std__pe54__lane9_strm1_data_valid ),      
               .std__pe54__lane9_strm1_data_mask     ( std__pe54__lane9_strm1_data_mask  ),      

               // PE 54, Lane 10                 
               .pe54__std__lane10_strm0_ready         ( pe54__std__lane10_strm0_ready      ),      
               .std__pe54__lane10_strm0_cntl          ( std__pe54__lane10_strm0_cntl       ),      
               .std__pe54__lane10_strm0_data          ( std__pe54__lane10_strm0_data       ),      
               .std__pe54__lane10_strm0_data_valid    ( std__pe54__lane10_strm0_data_valid ),      
               .std__pe54__lane10_strm0_data_mask     ( std__pe54__lane10_strm0_data_mask  ),      

               .pe54__std__lane10_strm1_ready         ( pe54__std__lane10_strm1_ready      ),      
               .std__pe54__lane10_strm1_cntl          ( std__pe54__lane10_strm1_cntl       ),      
               .std__pe54__lane10_strm1_data          ( std__pe54__lane10_strm1_data       ),      
               .std__pe54__lane10_strm1_data_valid    ( std__pe54__lane10_strm1_data_valid ),      
               .std__pe54__lane10_strm1_data_mask     ( std__pe54__lane10_strm1_data_mask  ),      

               // PE 54, Lane 11                 
               .pe54__std__lane11_strm0_ready         ( pe54__std__lane11_strm0_ready      ),      
               .std__pe54__lane11_strm0_cntl          ( std__pe54__lane11_strm0_cntl       ),      
               .std__pe54__lane11_strm0_data          ( std__pe54__lane11_strm0_data       ),      
               .std__pe54__lane11_strm0_data_valid    ( std__pe54__lane11_strm0_data_valid ),      
               .std__pe54__lane11_strm0_data_mask     ( std__pe54__lane11_strm0_data_mask  ),      

               .pe54__std__lane11_strm1_ready         ( pe54__std__lane11_strm1_ready      ),      
               .std__pe54__lane11_strm1_cntl          ( std__pe54__lane11_strm1_cntl       ),      
               .std__pe54__lane11_strm1_data          ( std__pe54__lane11_strm1_data       ),      
               .std__pe54__lane11_strm1_data_valid    ( std__pe54__lane11_strm1_data_valid ),      
               .std__pe54__lane11_strm1_data_mask     ( std__pe54__lane11_strm1_data_mask  ),      

               // PE 54, Lane 12                 
               .pe54__std__lane12_strm0_ready         ( pe54__std__lane12_strm0_ready      ),      
               .std__pe54__lane12_strm0_cntl          ( std__pe54__lane12_strm0_cntl       ),      
               .std__pe54__lane12_strm0_data          ( std__pe54__lane12_strm0_data       ),      
               .std__pe54__lane12_strm0_data_valid    ( std__pe54__lane12_strm0_data_valid ),      
               .std__pe54__lane12_strm0_data_mask     ( std__pe54__lane12_strm0_data_mask  ),      

               .pe54__std__lane12_strm1_ready         ( pe54__std__lane12_strm1_ready      ),      
               .std__pe54__lane12_strm1_cntl          ( std__pe54__lane12_strm1_cntl       ),      
               .std__pe54__lane12_strm1_data          ( std__pe54__lane12_strm1_data       ),      
               .std__pe54__lane12_strm1_data_valid    ( std__pe54__lane12_strm1_data_valid ),      
               .std__pe54__lane12_strm1_data_mask     ( std__pe54__lane12_strm1_data_mask  ),      

               // PE 54, Lane 13                 
               .pe54__std__lane13_strm0_ready         ( pe54__std__lane13_strm0_ready      ),      
               .std__pe54__lane13_strm0_cntl          ( std__pe54__lane13_strm0_cntl       ),      
               .std__pe54__lane13_strm0_data          ( std__pe54__lane13_strm0_data       ),      
               .std__pe54__lane13_strm0_data_valid    ( std__pe54__lane13_strm0_data_valid ),      
               .std__pe54__lane13_strm0_data_mask     ( std__pe54__lane13_strm0_data_mask  ),      

               .pe54__std__lane13_strm1_ready         ( pe54__std__lane13_strm1_ready      ),      
               .std__pe54__lane13_strm1_cntl          ( std__pe54__lane13_strm1_cntl       ),      
               .std__pe54__lane13_strm1_data          ( std__pe54__lane13_strm1_data       ),      
               .std__pe54__lane13_strm1_data_valid    ( std__pe54__lane13_strm1_data_valid ),      
               .std__pe54__lane13_strm1_data_mask     ( std__pe54__lane13_strm1_data_mask  ),      

               // PE 54, Lane 14                 
               .pe54__std__lane14_strm0_ready         ( pe54__std__lane14_strm0_ready      ),      
               .std__pe54__lane14_strm0_cntl          ( std__pe54__lane14_strm0_cntl       ),      
               .std__pe54__lane14_strm0_data          ( std__pe54__lane14_strm0_data       ),      
               .std__pe54__lane14_strm0_data_valid    ( std__pe54__lane14_strm0_data_valid ),      
               .std__pe54__lane14_strm0_data_mask     ( std__pe54__lane14_strm0_data_mask  ),      

               .pe54__std__lane14_strm1_ready         ( pe54__std__lane14_strm1_ready      ),      
               .std__pe54__lane14_strm1_cntl          ( std__pe54__lane14_strm1_cntl       ),      
               .std__pe54__lane14_strm1_data          ( std__pe54__lane14_strm1_data       ),      
               .std__pe54__lane14_strm1_data_valid    ( std__pe54__lane14_strm1_data_valid ),      
               .std__pe54__lane14_strm1_data_mask     ( std__pe54__lane14_strm1_data_mask  ),      

               // PE 54, Lane 15                 
               .pe54__std__lane15_strm0_ready         ( pe54__std__lane15_strm0_ready      ),      
               .std__pe54__lane15_strm0_cntl          ( std__pe54__lane15_strm0_cntl       ),      
               .std__pe54__lane15_strm0_data          ( std__pe54__lane15_strm0_data       ),      
               .std__pe54__lane15_strm0_data_valid    ( std__pe54__lane15_strm0_data_valid ),      
               .std__pe54__lane15_strm0_data_mask     ( std__pe54__lane15_strm0_data_mask  ),      

               .pe54__std__lane15_strm1_ready         ( pe54__std__lane15_strm1_ready      ),      
               .std__pe54__lane15_strm1_cntl          ( std__pe54__lane15_strm1_cntl       ),      
               .std__pe54__lane15_strm1_data          ( std__pe54__lane15_strm1_data       ),      
               .std__pe54__lane15_strm1_data_valid    ( std__pe54__lane15_strm1_data_valid ),      
               .std__pe54__lane15_strm1_data_mask     ( std__pe54__lane15_strm1_data_mask  ),      

               // PE 54, Lane 16                 
               .pe54__std__lane16_strm0_ready         ( pe54__std__lane16_strm0_ready      ),      
               .std__pe54__lane16_strm0_cntl          ( std__pe54__lane16_strm0_cntl       ),      
               .std__pe54__lane16_strm0_data          ( std__pe54__lane16_strm0_data       ),      
               .std__pe54__lane16_strm0_data_valid    ( std__pe54__lane16_strm0_data_valid ),      
               .std__pe54__lane16_strm0_data_mask     ( std__pe54__lane16_strm0_data_mask  ),      

               .pe54__std__lane16_strm1_ready         ( pe54__std__lane16_strm1_ready      ),      
               .std__pe54__lane16_strm1_cntl          ( std__pe54__lane16_strm1_cntl       ),      
               .std__pe54__lane16_strm1_data          ( std__pe54__lane16_strm1_data       ),      
               .std__pe54__lane16_strm1_data_valid    ( std__pe54__lane16_strm1_data_valid ),      
               .std__pe54__lane16_strm1_data_mask     ( std__pe54__lane16_strm1_data_mask  ),      

               // PE 54, Lane 17                 
               .pe54__std__lane17_strm0_ready         ( pe54__std__lane17_strm0_ready      ),      
               .std__pe54__lane17_strm0_cntl          ( std__pe54__lane17_strm0_cntl       ),      
               .std__pe54__lane17_strm0_data          ( std__pe54__lane17_strm0_data       ),      
               .std__pe54__lane17_strm0_data_valid    ( std__pe54__lane17_strm0_data_valid ),      
               .std__pe54__lane17_strm0_data_mask     ( std__pe54__lane17_strm0_data_mask  ),      

               .pe54__std__lane17_strm1_ready         ( pe54__std__lane17_strm1_ready      ),      
               .std__pe54__lane17_strm1_cntl          ( std__pe54__lane17_strm1_cntl       ),      
               .std__pe54__lane17_strm1_data          ( std__pe54__lane17_strm1_data       ),      
               .std__pe54__lane17_strm1_data_valid    ( std__pe54__lane17_strm1_data_valid ),      
               .std__pe54__lane17_strm1_data_mask     ( std__pe54__lane17_strm1_data_mask  ),      

               // PE 54, Lane 18                 
               .pe54__std__lane18_strm0_ready         ( pe54__std__lane18_strm0_ready      ),      
               .std__pe54__lane18_strm0_cntl          ( std__pe54__lane18_strm0_cntl       ),      
               .std__pe54__lane18_strm0_data          ( std__pe54__lane18_strm0_data       ),      
               .std__pe54__lane18_strm0_data_valid    ( std__pe54__lane18_strm0_data_valid ),      
               .std__pe54__lane18_strm0_data_mask     ( std__pe54__lane18_strm0_data_mask  ),      

               .pe54__std__lane18_strm1_ready         ( pe54__std__lane18_strm1_ready      ),      
               .std__pe54__lane18_strm1_cntl          ( std__pe54__lane18_strm1_cntl       ),      
               .std__pe54__lane18_strm1_data          ( std__pe54__lane18_strm1_data       ),      
               .std__pe54__lane18_strm1_data_valid    ( std__pe54__lane18_strm1_data_valid ),      
               .std__pe54__lane18_strm1_data_mask     ( std__pe54__lane18_strm1_data_mask  ),      

               // PE 54, Lane 19                 
               .pe54__std__lane19_strm0_ready         ( pe54__std__lane19_strm0_ready      ),      
               .std__pe54__lane19_strm0_cntl          ( std__pe54__lane19_strm0_cntl       ),      
               .std__pe54__lane19_strm0_data          ( std__pe54__lane19_strm0_data       ),      
               .std__pe54__lane19_strm0_data_valid    ( std__pe54__lane19_strm0_data_valid ),      
               .std__pe54__lane19_strm0_data_mask     ( std__pe54__lane19_strm0_data_mask  ),      

               .pe54__std__lane19_strm1_ready         ( pe54__std__lane19_strm1_ready      ),      
               .std__pe54__lane19_strm1_cntl          ( std__pe54__lane19_strm1_cntl       ),      
               .std__pe54__lane19_strm1_data          ( std__pe54__lane19_strm1_data       ),      
               .std__pe54__lane19_strm1_data_valid    ( std__pe54__lane19_strm1_data_valid ),      
               .std__pe54__lane19_strm1_data_mask     ( std__pe54__lane19_strm1_data_mask  ),      

               // PE 54, Lane 20                 
               .pe54__std__lane20_strm0_ready         ( pe54__std__lane20_strm0_ready      ),      
               .std__pe54__lane20_strm0_cntl          ( std__pe54__lane20_strm0_cntl       ),      
               .std__pe54__lane20_strm0_data          ( std__pe54__lane20_strm0_data       ),      
               .std__pe54__lane20_strm0_data_valid    ( std__pe54__lane20_strm0_data_valid ),      
               .std__pe54__lane20_strm0_data_mask     ( std__pe54__lane20_strm0_data_mask  ),      

               .pe54__std__lane20_strm1_ready         ( pe54__std__lane20_strm1_ready      ),      
               .std__pe54__lane20_strm1_cntl          ( std__pe54__lane20_strm1_cntl       ),      
               .std__pe54__lane20_strm1_data          ( std__pe54__lane20_strm1_data       ),      
               .std__pe54__lane20_strm1_data_valid    ( std__pe54__lane20_strm1_data_valid ),      
               .std__pe54__lane20_strm1_data_mask     ( std__pe54__lane20_strm1_data_mask  ),      

               // PE 54, Lane 21                 
               .pe54__std__lane21_strm0_ready         ( pe54__std__lane21_strm0_ready      ),      
               .std__pe54__lane21_strm0_cntl          ( std__pe54__lane21_strm0_cntl       ),      
               .std__pe54__lane21_strm0_data          ( std__pe54__lane21_strm0_data       ),      
               .std__pe54__lane21_strm0_data_valid    ( std__pe54__lane21_strm0_data_valid ),      
               .std__pe54__lane21_strm0_data_mask     ( std__pe54__lane21_strm0_data_mask  ),      

               .pe54__std__lane21_strm1_ready         ( pe54__std__lane21_strm1_ready      ),      
               .std__pe54__lane21_strm1_cntl          ( std__pe54__lane21_strm1_cntl       ),      
               .std__pe54__lane21_strm1_data          ( std__pe54__lane21_strm1_data       ),      
               .std__pe54__lane21_strm1_data_valid    ( std__pe54__lane21_strm1_data_valid ),      
               .std__pe54__lane21_strm1_data_mask     ( std__pe54__lane21_strm1_data_mask  ),      

               // PE 54, Lane 22                 
               .pe54__std__lane22_strm0_ready         ( pe54__std__lane22_strm0_ready      ),      
               .std__pe54__lane22_strm0_cntl          ( std__pe54__lane22_strm0_cntl       ),      
               .std__pe54__lane22_strm0_data          ( std__pe54__lane22_strm0_data       ),      
               .std__pe54__lane22_strm0_data_valid    ( std__pe54__lane22_strm0_data_valid ),      
               .std__pe54__lane22_strm0_data_mask     ( std__pe54__lane22_strm0_data_mask  ),      

               .pe54__std__lane22_strm1_ready         ( pe54__std__lane22_strm1_ready      ),      
               .std__pe54__lane22_strm1_cntl          ( std__pe54__lane22_strm1_cntl       ),      
               .std__pe54__lane22_strm1_data          ( std__pe54__lane22_strm1_data       ),      
               .std__pe54__lane22_strm1_data_valid    ( std__pe54__lane22_strm1_data_valid ),      
               .std__pe54__lane22_strm1_data_mask     ( std__pe54__lane22_strm1_data_mask  ),      

               // PE 54, Lane 23                 
               .pe54__std__lane23_strm0_ready         ( pe54__std__lane23_strm0_ready      ),      
               .std__pe54__lane23_strm0_cntl          ( std__pe54__lane23_strm0_cntl       ),      
               .std__pe54__lane23_strm0_data          ( std__pe54__lane23_strm0_data       ),      
               .std__pe54__lane23_strm0_data_valid    ( std__pe54__lane23_strm0_data_valid ),      
               .std__pe54__lane23_strm0_data_mask     ( std__pe54__lane23_strm0_data_mask  ),      

               .pe54__std__lane23_strm1_ready         ( pe54__std__lane23_strm1_ready      ),      
               .std__pe54__lane23_strm1_cntl          ( std__pe54__lane23_strm1_cntl       ),      
               .std__pe54__lane23_strm1_data          ( std__pe54__lane23_strm1_data       ),      
               .std__pe54__lane23_strm1_data_valid    ( std__pe54__lane23_strm1_data_valid ),      
               .std__pe54__lane23_strm1_data_mask     ( std__pe54__lane23_strm1_data_mask  ),      

               // PE 54, Lane 24                 
               .pe54__std__lane24_strm0_ready         ( pe54__std__lane24_strm0_ready      ),      
               .std__pe54__lane24_strm0_cntl          ( std__pe54__lane24_strm0_cntl       ),      
               .std__pe54__lane24_strm0_data          ( std__pe54__lane24_strm0_data       ),      
               .std__pe54__lane24_strm0_data_valid    ( std__pe54__lane24_strm0_data_valid ),      
               .std__pe54__lane24_strm0_data_mask     ( std__pe54__lane24_strm0_data_mask  ),      

               .pe54__std__lane24_strm1_ready         ( pe54__std__lane24_strm1_ready      ),      
               .std__pe54__lane24_strm1_cntl          ( std__pe54__lane24_strm1_cntl       ),      
               .std__pe54__lane24_strm1_data          ( std__pe54__lane24_strm1_data       ),      
               .std__pe54__lane24_strm1_data_valid    ( std__pe54__lane24_strm1_data_valid ),      
               .std__pe54__lane24_strm1_data_mask     ( std__pe54__lane24_strm1_data_mask  ),      

               // PE 54, Lane 25                 
               .pe54__std__lane25_strm0_ready         ( pe54__std__lane25_strm0_ready      ),      
               .std__pe54__lane25_strm0_cntl          ( std__pe54__lane25_strm0_cntl       ),      
               .std__pe54__lane25_strm0_data          ( std__pe54__lane25_strm0_data       ),      
               .std__pe54__lane25_strm0_data_valid    ( std__pe54__lane25_strm0_data_valid ),      
               .std__pe54__lane25_strm0_data_mask     ( std__pe54__lane25_strm0_data_mask  ),      

               .pe54__std__lane25_strm1_ready         ( pe54__std__lane25_strm1_ready      ),      
               .std__pe54__lane25_strm1_cntl          ( std__pe54__lane25_strm1_cntl       ),      
               .std__pe54__lane25_strm1_data          ( std__pe54__lane25_strm1_data       ),      
               .std__pe54__lane25_strm1_data_valid    ( std__pe54__lane25_strm1_data_valid ),      
               .std__pe54__lane25_strm1_data_mask     ( std__pe54__lane25_strm1_data_mask  ),      

               // PE 54, Lane 26                 
               .pe54__std__lane26_strm0_ready         ( pe54__std__lane26_strm0_ready      ),      
               .std__pe54__lane26_strm0_cntl          ( std__pe54__lane26_strm0_cntl       ),      
               .std__pe54__lane26_strm0_data          ( std__pe54__lane26_strm0_data       ),      
               .std__pe54__lane26_strm0_data_valid    ( std__pe54__lane26_strm0_data_valid ),      
               .std__pe54__lane26_strm0_data_mask     ( std__pe54__lane26_strm0_data_mask  ),      

               .pe54__std__lane26_strm1_ready         ( pe54__std__lane26_strm1_ready      ),      
               .std__pe54__lane26_strm1_cntl          ( std__pe54__lane26_strm1_cntl       ),      
               .std__pe54__lane26_strm1_data          ( std__pe54__lane26_strm1_data       ),      
               .std__pe54__lane26_strm1_data_valid    ( std__pe54__lane26_strm1_data_valid ),      
               .std__pe54__lane26_strm1_data_mask     ( std__pe54__lane26_strm1_data_mask  ),      

               // PE 54, Lane 27                 
               .pe54__std__lane27_strm0_ready         ( pe54__std__lane27_strm0_ready      ),      
               .std__pe54__lane27_strm0_cntl          ( std__pe54__lane27_strm0_cntl       ),      
               .std__pe54__lane27_strm0_data          ( std__pe54__lane27_strm0_data       ),      
               .std__pe54__lane27_strm0_data_valid    ( std__pe54__lane27_strm0_data_valid ),      
               .std__pe54__lane27_strm0_data_mask     ( std__pe54__lane27_strm0_data_mask  ),      

               .pe54__std__lane27_strm1_ready         ( pe54__std__lane27_strm1_ready      ),      
               .std__pe54__lane27_strm1_cntl          ( std__pe54__lane27_strm1_cntl       ),      
               .std__pe54__lane27_strm1_data          ( std__pe54__lane27_strm1_data       ),      
               .std__pe54__lane27_strm1_data_valid    ( std__pe54__lane27_strm1_data_valid ),      
               .std__pe54__lane27_strm1_data_mask     ( std__pe54__lane27_strm1_data_mask  ),      

               // PE 54, Lane 28                 
               .pe54__std__lane28_strm0_ready         ( pe54__std__lane28_strm0_ready      ),      
               .std__pe54__lane28_strm0_cntl          ( std__pe54__lane28_strm0_cntl       ),      
               .std__pe54__lane28_strm0_data          ( std__pe54__lane28_strm0_data       ),      
               .std__pe54__lane28_strm0_data_valid    ( std__pe54__lane28_strm0_data_valid ),      
               .std__pe54__lane28_strm0_data_mask     ( std__pe54__lane28_strm0_data_mask  ),      

               .pe54__std__lane28_strm1_ready         ( pe54__std__lane28_strm1_ready      ),      
               .std__pe54__lane28_strm1_cntl          ( std__pe54__lane28_strm1_cntl       ),      
               .std__pe54__lane28_strm1_data          ( std__pe54__lane28_strm1_data       ),      
               .std__pe54__lane28_strm1_data_valid    ( std__pe54__lane28_strm1_data_valid ),      
               .std__pe54__lane28_strm1_data_mask     ( std__pe54__lane28_strm1_data_mask  ),      

               // PE 54, Lane 29                 
               .pe54__std__lane29_strm0_ready         ( pe54__std__lane29_strm0_ready      ),      
               .std__pe54__lane29_strm0_cntl          ( std__pe54__lane29_strm0_cntl       ),      
               .std__pe54__lane29_strm0_data          ( std__pe54__lane29_strm0_data       ),      
               .std__pe54__lane29_strm0_data_valid    ( std__pe54__lane29_strm0_data_valid ),      
               .std__pe54__lane29_strm0_data_mask     ( std__pe54__lane29_strm0_data_mask  ),      

               .pe54__std__lane29_strm1_ready         ( pe54__std__lane29_strm1_ready      ),      
               .std__pe54__lane29_strm1_cntl          ( std__pe54__lane29_strm1_cntl       ),      
               .std__pe54__lane29_strm1_data          ( std__pe54__lane29_strm1_data       ),      
               .std__pe54__lane29_strm1_data_valid    ( std__pe54__lane29_strm1_data_valid ),      
               .std__pe54__lane29_strm1_data_mask     ( std__pe54__lane29_strm1_data_mask  ),      

               // PE 54, Lane 30                 
               .pe54__std__lane30_strm0_ready         ( pe54__std__lane30_strm0_ready      ),      
               .std__pe54__lane30_strm0_cntl          ( std__pe54__lane30_strm0_cntl       ),      
               .std__pe54__lane30_strm0_data          ( std__pe54__lane30_strm0_data       ),      
               .std__pe54__lane30_strm0_data_valid    ( std__pe54__lane30_strm0_data_valid ),      
               .std__pe54__lane30_strm0_data_mask     ( std__pe54__lane30_strm0_data_mask  ),      

               .pe54__std__lane30_strm1_ready         ( pe54__std__lane30_strm1_ready      ),      
               .std__pe54__lane30_strm1_cntl          ( std__pe54__lane30_strm1_cntl       ),      
               .std__pe54__lane30_strm1_data          ( std__pe54__lane30_strm1_data       ),      
               .std__pe54__lane30_strm1_data_valid    ( std__pe54__lane30_strm1_data_valid ),      
               .std__pe54__lane30_strm1_data_mask     ( std__pe54__lane30_strm1_data_mask  ),      

               // PE 54, Lane 31                 
               .pe54__std__lane31_strm0_ready         ( pe54__std__lane31_strm0_ready      ),      
               .std__pe54__lane31_strm0_cntl          ( std__pe54__lane31_strm0_cntl       ),      
               .std__pe54__lane31_strm0_data          ( std__pe54__lane31_strm0_data       ),      
               .std__pe54__lane31_strm0_data_valid    ( std__pe54__lane31_strm0_data_valid ),      
               .std__pe54__lane31_strm0_data_mask     ( std__pe54__lane31_strm0_data_mask  ),      

               .pe54__std__lane31_strm1_ready         ( pe54__std__lane31_strm1_ready      ),      
               .std__pe54__lane31_strm1_cntl          ( std__pe54__lane31_strm1_cntl       ),      
               .std__pe54__lane31_strm1_data          ( std__pe54__lane31_strm1_data       ),      
               .std__pe54__lane31_strm1_data_valid    ( std__pe54__lane31_strm1_data_valid ),      
               .std__pe54__lane31_strm1_data_mask     ( std__pe54__lane31_strm1_data_mask  ),      

               // PE 55, Lane 0                 
               .pe55__std__lane0_strm0_ready         ( pe55__std__lane0_strm0_ready      ),      
               .std__pe55__lane0_strm0_cntl          ( std__pe55__lane0_strm0_cntl       ),      
               .std__pe55__lane0_strm0_data          ( std__pe55__lane0_strm0_data       ),      
               .std__pe55__lane0_strm0_data_valid    ( std__pe55__lane0_strm0_data_valid ),      
               .std__pe55__lane0_strm0_data_mask     ( std__pe55__lane0_strm0_data_mask  ),      

               .pe55__std__lane0_strm1_ready         ( pe55__std__lane0_strm1_ready      ),      
               .std__pe55__lane0_strm1_cntl          ( std__pe55__lane0_strm1_cntl       ),      
               .std__pe55__lane0_strm1_data          ( std__pe55__lane0_strm1_data       ),      
               .std__pe55__lane0_strm1_data_valid    ( std__pe55__lane0_strm1_data_valid ),      
               .std__pe55__lane0_strm1_data_mask     ( std__pe55__lane0_strm1_data_mask  ),      

               // PE 55, Lane 1                 
               .pe55__std__lane1_strm0_ready         ( pe55__std__lane1_strm0_ready      ),      
               .std__pe55__lane1_strm0_cntl          ( std__pe55__lane1_strm0_cntl       ),      
               .std__pe55__lane1_strm0_data          ( std__pe55__lane1_strm0_data       ),      
               .std__pe55__lane1_strm0_data_valid    ( std__pe55__lane1_strm0_data_valid ),      
               .std__pe55__lane1_strm0_data_mask     ( std__pe55__lane1_strm0_data_mask  ),      

               .pe55__std__lane1_strm1_ready         ( pe55__std__lane1_strm1_ready      ),      
               .std__pe55__lane1_strm1_cntl          ( std__pe55__lane1_strm1_cntl       ),      
               .std__pe55__lane1_strm1_data          ( std__pe55__lane1_strm1_data       ),      
               .std__pe55__lane1_strm1_data_valid    ( std__pe55__lane1_strm1_data_valid ),      
               .std__pe55__lane1_strm1_data_mask     ( std__pe55__lane1_strm1_data_mask  ),      

               // PE 55, Lane 2                 
               .pe55__std__lane2_strm0_ready         ( pe55__std__lane2_strm0_ready      ),      
               .std__pe55__lane2_strm0_cntl          ( std__pe55__lane2_strm0_cntl       ),      
               .std__pe55__lane2_strm0_data          ( std__pe55__lane2_strm0_data       ),      
               .std__pe55__lane2_strm0_data_valid    ( std__pe55__lane2_strm0_data_valid ),      
               .std__pe55__lane2_strm0_data_mask     ( std__pe55__lane2_strm0_data_mask  ),      

               .pe55__std__lane2_strm1_ready         ( pe55__std__lane2_strm1_ready      ),      
               .std__pe55__lane2_strm1_cntl          ( std__pe55__lane2_strm1_cntl       ),      
               .std__pe55__lane2_strm1_data          ( std__pe55__lane2_strm1_data       ),      
               .std__pe55__lane2_strm1_data_valid    ( std__pe55__lane2_strm1_data_valid ),      
               .std__pe55__lane2_strm1_data_mask     ( std__pe55__lane2_strm1_data_mask  ),      

               // PE 55, Lane 3                 
               .pe55__std__lane3_strm0_ready         ( pe55__std__lane3_strm0_ready      ),      
               .std__pe55__lane3_strm0_cntl          ( std__pe55__lane3_strm0_cntl       ),      
               .std__pe55__lane3_strm0_data          ( std__pe55__lane3_strm0_data       ),      
               .std__pe55__lane3_strm0_data_valid    ( std__pe55__lane3_strm0_data_valid ),      
               .std__pe55__lane3_strm0_data_mask     ( std__pe55__lane3_strm0_data_mask  ),      

               .pe55__std__lane3_strm1_ready         ( pe55__std__lane3_strm1_ready      ),      
               .std__pe55__lane3_strm1_cntl          ( std__pe55__lane3_strm1_cntl       ),      
               .std__pe55__lane3_strm1_data          ( std__pe55__lane3_strm1_data       ),      
               .std__pe55__lane3_strm1_data_valid    ( std__pe55__lane3_strm1_data_valid ),      
               .std__pe55__lane3_strm1_data_mask     ( std__pe55__lane3_strm1_data_mask  ),      

               // PE 55, Lane 4                 
               .pe55__std__lane4_strm0_ready         ( pe55__std__lane4_strm0_ready      ),      
               .std__pe55__lane4_strm0_cntl          ( std__pe55__lane4_strm0_cntl       ),      
               .std__pe55__lane4_strm0_data          ( std__pe55__lane4_strm0_data       ),      
               .std__pe55__lane4_strm0_data_valid    ( std__pe55__lane4_strm0_data_valid ),      
               .std__pe55__lane4_strm0_data_mask     ( std__pe55__lane4_strm0_data_mask  ),      

               .pe55__std__lane4_strm1_ready         ( pe55__std__lane4_strm1_ready      ),      
               .std__pe55__lane4_strm1_cntl          ( std__pe55__lane4_strm1_cntl       ),      
               .std__pe55__lane4_strm1_data          ( std__pe55__lane4_strm1_data       ),      
               .std__pe55__lane4_strm1_data_valid    ( std__pe55__lane4_strm1_data_valid ),      
               .std__pe55__lane4_strm1_data_mask     ( std__pe55__lane4_strm1_data_mask  ),      

               // PE 55, Lane 5                 
               .pe55__std__lane5_strm0_ready         ( pe55__std__lane5_strm0_ready      ),      
               .std__pe55__lane5_strm0_cntl          ( std__pe55__lane5_strm0_cntl       ),      
               .std__pe55__lane5_strm0_data          ( std__pe55__lane5_strm0_data       ),      
               .std__pe55__lane5_strm0_data_valid    ( std__pe55__lane5_strm0_data_valid ),      
               .std__pe55__lane5_strm0_data_mask     ( std__pe55__lane5_strm0_data_mask  ),      

               .pe55__std__lane5_strm1_ready         ( pe55__std__lane5_strm1_ready      ),      
               .std__pe55__lane5_strm1_cntl          ( std__pe55__lane5_strm1_cntl       ),      
               .std__pe55__lane5_strm1_data          ( std__pe55__lane5_strm1_data       ),      
               .std__pe55__lane5_strm1_data_valid    ( std__pe55__lane5_strm1_data_valid ),      
               .std__pe55__lane5_strm1_data_mask     ( std__pe55__lane5_strm1_data_mask  ),      

               // PE 55, Lane 6                 
               .pe55__std__lane6_strm0_ready         ( pe55__std__lane6_strm0_ready      ),      
               .std__pe55__lane6_strm0_cntl          ( std__pe55__lane6_strm0_cntl       ),      
               .std__pe55__lane6_strm0_data          ( std__pe55__lane6_strm0_data       ),      
               .std__pe55__lane6_strm0_data_valid    ( std__pe55__lane6_strm0_data_valid ),      
               .std__pe55__lane6_strm0_data_mask     ( std__pe55__lane6_strm0_data_mask  ),      

               .pe55__std__lane6_strm1_ready         ( pe55__std__lane6_strm1_ready      ),      
               .std__pe55__lane6_strm1_cntl          ( std__pe55__lane6_strm1_cntl       ),      
               .std__pe55__lane6_strm1_data          ( std__pe55__lane6_strm1_data       ),      
               .std__pe55__lane6_strm1_data_valid    ( std__pe55__lane6_strm1_data_valid ),      
               .std__pe55__lane6_strm1_data_mask     ( std__pe55__lane6_strm1_data_mask  ),      

               // PE 55, Lane 7                 
               .pe55__std__lane7_strm0_ready         ( pe55__std__lane7_strm0_ready      ),      
               .std__pe55__lane7_strm0_cntl          ( std__pe55__lane7_strm0_cntl       ),      
               .std__pe55__lane7_strm0_data          ( std__pe55__lane7_strm0_data       ),      
               .std__pe55__lane7_strm0_data_valid    ( std__pe55__lane7_strm0_data_valid ),      
               .std__pe55__lane7_strm0_data_mask     ( std__pe55__lane7_strm0_data_mask  ),      

               .pe55__std__lane7_strm1_ready         ( pe55__std__lane7_strm1_ready      ),      
               .std__pe55__lane7_strm1_cntl          ( std__pe55__lane7_strm1_cntl       ),      
               .std__pe55__lane7_strm1_data          ( std__pe55__lane7_strm1_data       ),      
               .std__pe55__lane7_strm1_data_valid    ( std__pe55__lane7_strm1_data_valid ),      
               .std__pe55__lane7_strm1_data_mask     ( std__pe55__lane7_strm1_data_mask  ),      

               // PE 55, Lane 8                 
               .pe55__std__lane8_strm0_ready         ( pe55__std__lane8_strm0_ready      ),      
               .std__pe55__lane8_strm0_cntl          ( std__pe55__lane8_strm0_cntl       ),      
               .std__pe55__lane8_strm0_data          ( std__pe55__lane8_strm0_data       ),      
               .std__pe55__lane8_strm0_data_valid    ( std__pe55__lane8_strm0_data_valid ),      
               .std__pe55__lane8_strm0_data_mask     ( std__pe55__lane8_strm0_data_mask  ),      

               .pe55__std__lane8_strm1_ready         ( pe55__std__lane8_strm1_ready      ),      
               .std__pe55__lane8_strm1_cntl          ( std__pe55__lane8_strm1_cntl       ),      
               .std__pe55__lane8_strm1_data          ( std__pe55__lane8_strm1_data       ),      
               .std__pe55__lane8_strm1_data_valid    ( std__pe55__lane8_strm1_data_valid ),      
               .std__pe55__lane8_strm1_data_mask     ( std__pe55__lane8_strm1_data_mask  ),      

               // PE 55, Lane 9                 
               .pe55__std__lane9_strm0_ready         ( pe55__std__lane9_strm0_ready      ),      
               .std__pe55__lane9_strm0_cntl          ( std__pe55__lane9_strm0_cntl       ),      
               .std__pe55__lane9_strm0_data          ( std__pe55__lane9_strm0_data       ),      
               .std__pe55__lane9_strm0_data_valid    ( std__pe55__lane9_strm0_data_valid ),      
               .std__pe55__lane9_strm0_data_mask     ( std__pe55__lane9_strm0_data_mask  ),      

               .pe55__std__lane9_strm1_ready         ( pe55__std__lane9_strm1_ready      ),      
               .std__pe55__lane9_strm1_cntl          ( std__pe55__lane9_strm1_cntl       ),      
               .std__pe55__lane9_strm1_data          ( std__pe55__lane9_strm1_data       ),      
               .std__pe55__lane9_strm1_data_valid    ( std__pe55__lane9_strm1_data_valid ),      
               .std__pe55__lane9_strm1_data_mask     ( std__pe55__lane9_strm1_data_mask  ),      

               // PE 55, Lane 10                 
               .pe55__std__lane10_strm0_ready         ( pe55__std__lane10_strm0_ready      ),      
               .std__pe55__lane10_strm0_cntl          ( std__pe55__lane10_strm0_cntl       ),      
               .std__pe55__lane10_strm0_data          ( std__pe55__lane10_strm0_data       ),      
               .std__pe55__lane10_strm0_data_valid    ( std__pe55__lane10_strm0_data_valid ),      
               .std__pe55__lane10_strm0_data_mask     ( std__pe55__lane10_strm0_data_mask  ),      

               .pe55__std__lane10_strm1_ready         ( pe55__std__lane10_strm1_ready      ),      
               .std__pe55__lane10_strm1_cntl          ( std__pe55__lane10_strm1_cntl       ),      
               .std__pe55__lane10_strm1_data          ( std__pe55__lane10_strm1_data       ),      
               .std__pe55__lane10_strm1_data_valid    ( std__pe55__lane10_strm1_data_valid ),      
               .std__pe55__lane10_strm1_data_mask     ( std__pe55__lane10_strm1_data_mask  ),      

               // PE 55, Lane 11                 
               .pe55__std__lane11_strm0_ready         ( pe55__std__lane11_strm0_ready      ),      
               .std__pe55__lane11_strm0_cntl          ( std__pe55__lane11_strm0_cntl       ),      
               .std__pe55__lane11_strm0_data          ( std__pe55__lane11_strm0_data       ),      
               .std__pe55__lane11_strm0_data_valid    ( std__pe55__lane11_strm0_data_valid ),      
               .std__pe55__lane11_strm0_data_mask     ( std__pe55__lane11_strm0_data_mask  ),      

               .pe55__std__lane11_strm1_ready         ( pe55__std__lane11_strm1_ready      ),      
               .std__pe55__lane11_strm1_cntl          ( std__pe55__lane11_strm1_cntl       ),      
               .std__pe55__lane11_strm1_data          ( std__pe55__lane11_strm1_data       ),      
               .std__pe55__lane11_strm1_data_valid    ( std__pe55__lane11_strm1_data_valid ),      
               .std__pe55__lane11_strm1_data_mask     ( std__pe55__lane11_strm1_data_mask  ),      

               // PE 55, Lane 12                 
               .pe55__std__lane12_strm0_ready         ( pe55__std__lane12_strm0_ready      ),      
               .std__pe55__lane12_strm0_cntl          ( std__pe55__lane12_strm0_cntl       ),      
               .std__pe55__lane12_strm0_data          ( std__pe55__lane12_strm0_data       ),      
               .std__pe55__lane12_strm0_data_valid    ( std__pe55__lane12_strm0_data_valid ),      
               .std__pe55__lane12_strm0_data_mask     ( std__pe55__lane12_strm0_data_mask  ),      

               .pe55__std__lane12_strm1_ready         ( pe55__std__lane12_strm1_ready      ),      
               .std__pe55__lane12_strm1_cntl          ( std__pe55__lane12_strm1_cntl       ),      
               .std__pe55__lane12_strm1_data          ( std__pe55__lane12_strm1_data       ),      
               .std__pe55__lane12_strm1_data_valid    ( std__pe55__lane12_strm1_data_valid ),      
               .std__pe55__lane12_strm1_data_mask     ( std__pe55__lane12_strm1_data_mask  ),      

               // PE 55, Lane 13                 
               .pe55__std__lane13_strm0_ready         ( pe55__std__lane13_strm0_ready      ),      
               .std__pe55__lane13_strm0_cntl          ( std__pe55__lane13_strm0_cntl       ),      
               .std__pe55__lane13_strm0_data          ( std__pe55__lane13_strm0_data       ),      
               .std__pe55__lane13_strm0_data_valid    ( std__pe55__lane13_strm0_data_valid ),      
               .std__pe55__lane13_strm0_data_mask     ( std__pe55__lane13_strm0_data_mask  ),      

               .pe55__std__lane13_strm1_ready         ( pe55__std__lane13_strm1_ready      ),      
               .std__pe55__lane13_strm1_cntl          ( std__pe55__lane13_strm1_cntl       ),      
               .std__pe55__lane13_strm1_data          ( std__pe55__lane13_strm1_data       ),      
               .std__pe55__lane13_strm1_data_valid    ( std__pe55__lane13_strm1_data_valid ),      
               .std__pe55__lane13_strm1_data_mask     ( std__pe55__lane13_strm1_data_mask  ),      

               // PE 55, Lane 14                 
               .pe55__std__lane14_strm0_ready         ( pe55__std__lane14_strm0_ready      ),      
               .std__pe55__lane14_strm0_cntl          ( std__pe55__lane14_strm0_cntl       ),      
               .std__pe55__lane14_strm0_data          ( std__pe55__lane14_strm0_data       ),      
               .std__pe55__lane14_strm0_data_valid    ( std__pe55__lane14_strm0_data_valid ),      
               .std__pe55__lane14_strm0_data_mask     ( std__pe55__lane14_strm0_data_mask  ),      

               .pe55__std__lane14_strm1_ready         ( pe55__std__lane14_strm1_ready      ),      
               .std__pe55__lane14_strm1_cntl          ( std__pe55__lane14_strm1_cntl       ),      
               .std__pe55__lane14_strm1_data          ( std__pe55__lane14_strm1_data       ),      
               .std__pe55__lane14_strm1_data_valid    ( std__pe55__lane14_strm1_data_valid ),      
               .std__pe55__lane14_strm1_data_mask     ( std__pe55__lane14_strm1_data_mask  ),      

               // PE 55, Lane 15                 
               .pe55__std__lane15_strm0_ready         ( pe55__std__lane15_strm0_ready      ),      
               .std__pe55__lane15_strm0_cntl          ( std__pe55__lane15_strm0_cntl       ),      
               .std__pe55__lane15_strm0_data          ( std__pe55__lane15_strm0_data       ),      
               .std__pe55__lane15_strm0_data_valid    ( std__pe55__lane15_strm0_data_valid ),      
               .std__pe55__lane15_strm0_data_mask     ( std__pe55__lane15_strm0_data_mask  ),      

               .pe55__std__lane15_strm1_ready         ( pe55__std__lane15_strm1_ready      ),      
               .std__pe55__lane15_strm1_cntl          ( std__pe55__lane15_strm1_cntl       ),      
               .std__pe55__lane15_strm1_data          ( std__pe55__lane15_strm1_data       ),      
               .std__pe55__lane15_strm1_data_valid    ( std__pe55__lane15_strm1_data_valid ),      
               .std__pe55__lane15_strm1_data_mask     ( std__pe55__lane15_strm1_data_mask  ),      

               // PE 55, Lane 16                 
               .pe55__std__lane16_strm0_ready         ( pe55__std__lane16_strm0_ready      ),      
               .std__pe55__lane16_strm0_cntl          ( std__pe55__lane16_strm0_cntl       ),      
               .std__pe55__lane16_strm0_data          ( std__pe55__lane16_strm0_data       ),      
               .std__pe55__lane16_strm0_data_valid    ( std__pe55__lane16_strm0_data_valid ),      
               .std__pe55__lane16_strm0_data_mask     ( std__pe55__lane16_strm0_data_mask  ),      

               .pe55__std__lane16_strm1_ready         ( pe55__std__lane16_strm1_ready      ),      
               .std__pe55__lane16_strm1_cntl          ( std__pe55__lane16_strm1_cntl       ),      
               .std__pe55__lane16_strm1_data          ( std__pe55__lane16_strm1_data       ),      
               .std__pe55__lane16_strm1_data_valid    ( std__pe55__lane16_strm1_data_valid ),      
               .std__pe55__lane16_strm1_data_mask     ( std__pe55__lane16_strm1_data_mask  ),      

               // PE 55, Lane 17                 
               .pe55__std__lane17_strm0_ready         ( pe55__std__lane17_strm0_ready      ),      
               .std__pe55__lane17_strm0_cntl          ( std__pe55__lane17_strm0_cntl       ),      
               .std__pe55__lane17_strm0_data          ( std__pe55__lane17_strm0_data       ),      
               .std__pe55__lane17_strm0_data_valid    ( std__pe55__lane17_strm0_data_valid ),      
               .std__pe55__lane17_strm0_data_mask     ( std__pe55__lane17_strm0_data_mask  ),      

               .pe55__std__lane17_strm1_ready         ( pe55__std__lane17_strm1_ready      ),      
               .std__pe55__lane17_strm1_cntl          ( std__pe55__lane17_strm1_cntl       ),      
               .std__pe55__lane17_strm1_data          ( std__pe55__lane17_strm1_data       ),      
               .std__pe55__lane17_strm1_data_valid    ( std__pe55__lane17_strm1_data_valid ),      
               .std__pe55__lane17_strm1_data_mask     ( std__pe55__lane17_strm1_data_mask  ),      

               // PE 55, Lane 18                 
               .pe55__std__lane18_strm0_ready         ( pe55__std__lane18_strm0_ready      ),      
               .std__pe55__lane18_strm0_cntl          ( std__pe55__lane18_strm0_cntl       ),      
               .std__pe55__lane18_strm0_data          ( std__pe55__lane18_strm0_data       ),      
               .std__pe55__lane18_strm0_data_valid    ( std__pe55__lane18_strm0_data_valid ),      
               .std__pe55__lane18_strm0_data_mask     ( std__pe55__lane18_strm0_data_mask  ),      

               .pe55__std__lane18_strm1_ready         ( pe55__std__lane18_strm1_ready      ),      
               .std__pe55__lane18_strm1_cntl          ( std__pe55__lane18_strm1_cntl       ),      
               .std__pe55__lane18_strm1_data          ( std__pe55__lane18_strm1_data       ),      
               .std__pe55__lane18_strm1_data_valid    ( std__pe55__lane18_strm1_data_valid ),      
               .std__pe55__lane18_strm1_data_mask     ( std__pe55__lane18_strm1_data_mask  ),      

               // PE 55, Lane 19                 
               .pe55__std__lane19_strm0_ready         ( pe55__std__lane19_strm0_ready      ),      
               .std__pe55__lane19_strm0_cntl          ( std__pe55__lane19_strm0_cntl       ),      
               .std__pe55__lane19_strm0_data          ( std__pe55__lane19_strm0_data       ),      
               .std__pe55__lane19_strm0_data_valid    ( std__pe55__lane19_strm0_data_valid ),      
               .std__pe55__lane19_strm0_data_mask     ( std__pe55__lane19_strm0_data_mask  ),      

               .pe55__std__lane19_strm1_ready         ( pe55__std__lane19_strm1_ready      ),      
               .std__pe55__lane19_strm1_cntl          ( std__pe55__lane19_strm1_cntl       ),      
               .std__pe55__lane19_strm1_data          ( std__pe55__lane19_strm1_data       ),      
               .std__pe55__lane19_strm1_data_valid    ( std__pe55__lane19_strm1_data_valid ),      
               .std__pe55__lane19_strm1_data_mask     ( std__pe55__lane19_strm1_data_mask  ),      

               // PE 55, Lane 20                 
               .pe55__std__lane20_strm0_ready         ( pe55__std__lane20_strm0_ready      ),      
               .std__pe55__lane20_strm0_cntl          ( std__pe55__lane20_strm0_cntl       ),      
               .std__pe55__lane20_strm0_data          ( std__pe55__lane20_strm0_data       ),      
               .std__pe55__lane20_strm0_data_valid    ( std__pe55__lane20_strm0_data_valid ),      
               .std__pe55__lane20_strm0_data_mask     ( std__pe55__lane20_strm0_data_mask  ),      

               .pe55__std__lane20_strm1_ready         ( pe55__std__lane20_strm1_ready      ),      
               .std__pe55__lane20_strm1_cntl          ( std__pe55__lane20_strm1_cntl       ),      
               .std__pe55__lane20_strm1_data          ( std__pe55__lane20_strm1_data       ),      
               .std__pe55__lane20_strm1_data_valid    ( std__pe55__lane20_strm1_data_valid ),      
               .std__pe55__lane20_strm1_data_mask     ( std__pe55__lane20_strm1_data_mask  ),      

               // PE 55, Lane 21                 
               .pe55__std__lane21_strm0_ready         ( pe55__std__lane21_strm0_ready      ),      
               .std__pe55__lane21_strm0_cntl          ( std__pe55__lane21_strm0_cntl       ),      
               .std__pe55__lane21_strm0_data          ( std__pe55__lane21_strm0_data       ),      
               .std__pe55__lane21_strm0_data_valid    ( std__pe55__lane21_strm0_data_valid ),      
               .std__pe55__lane21_strm0_data_mask     ( std__pe55__lane21_strm0_data_mask  ),      

               .pe55__std__lane21_strm1_ready         ( pe55__std__lane21_strm1_ready      ),      
               .std__pe55__lane21_strm1_cntl          ( std__pe55__lane21_strm1_cntl       ),      
               .std__pe55__lane21_strm1_data          ( std__pe55__lane21_strm1_data       ),      
               .std__pe55__lane21_strm1_data_valid    ( std__pe55__lane21_strm1_data_valid ),      
               .std__pe55__lane21_strm1_data_mask     ( std__pe55__lane21_strm1_data_mask  ),      

               // PE 55, Lane 22                 
               .pe55__std__lane22_strm0_ready         ( pe55__std__lane22_strm0_ready      ),      
               .std__pe55__lane22_strm0_cntl          ( std__pe55__lane22_strm0_cntl       ),      
               .std__pe55__lane22_strm0_data          ( std__pe55__lane22_strm0_data       ),      
               .std__pe55__lane22_strm0_data_valid    ( std__pe55__lane22_strm0_data_valid ),      
               .std__pe55__lane22_strm0_data_mask     ( std__pe55__lane22_strm0_data_mask  ),      

               .pe55__std__lane22_strm1_ready         ( pe55__std__lane22_strm1_ready      ),      
               .std__pe55__lane22_strm1_cntl          ( std__pe55__lane22_strm1_cntl       ),      
               .std__pe55__lane22_strm1_data          ( std__pe55__lane22_strm1_data       ),      
               .std__pe55__lane22_strm1_data_valid    ( std__pe55__lane22_strm1_data_valid ),      
               .std__pe55__lane22_strm1_data_mask     ( std__pe55__lane22_strm1_data_mask  ),      

               // PE 55, Lane 23                 
               .pe55__std__lane23_strm0_ready         ( pe55__std__lane23_strm0_ready      ),      
               .std__pe55__lane23_strm0_cntl          ( std__pe55__lane23_strm0_cntl       ),      
               .std__pe55__lane23_strm0_data          ( std__pe55__lane23_strm0_data       ),      
               .std__pe55__lane23_strm0_data_valid    ( std__pe55__lane23_strm0_data_valid ),      
               .std__pe55__lane23_strm0_data_mask     ( std__pe55__lane23_strm0_data_mask  ),      

               .pe55__std__lane23_strm1_ready         ( pe55__std__lane23_strm1_ready      ),      
               .std__pe55__lane23_strm1_cntl          ( std__pe55__lane23_strm1_cntl       ),      
               .std__pe55__lane23_strm1_data          ( std__pe55__lane23_strm1_data       ),      
               .std__pe55__lane23_strm1_data_valid    ( std__pe55__lane23_strm1_data_valid ),      
               .std__pe55__lane23_strm1_data_mask     ( std__pe55__lane23_strm1_data_mask  ),      

               // PE 55, Lane 24                 
               .pe55__std__lane24_strm0_ready         ( pe55__std__lane24_strm0_ready      ),      
               .std__pe55__lane24_strm0_cntl          ( std__pe55__lane24_strm0_cntl       ),      
               .std__pe55__lane24_strm0_data          ( std__pe55__lane24_strm0_data       ),      
               .std__pe55__lane24_strm0_data_valid    ( std__pe55__lane24_strm0_data_valid ),      
               .std__pe55__lane24_strm0_data_mask     ( std__pe55__lane24_strm0_data_mask  ),      

               .pe55__std__lane24_strm1_ready         ( pe55__std__lane24_strm1_ready      ),      
               .std__pe55__lane24_strm1_cntl          ( std__pe55__lane24_strm1_cntl       ),      
               .std__pe55__lane24_strm1_data          ( std__pe55__lane24_strm1_data       ),      
               .std__pe55__lane24_strm1_data_valid    ( std__pe55__lane24_strm1_data_valid ),      
               .std__pe55__lane24_strm1_data_mask     ( std__pe55__lane24_strm1_data_mask  ),      

               // PE 55, Lane 25                 
               .pe55__std__lane25_strm0_ready         ( pe55__std__lane25_strm0_ready      ),      
               .std__pe55__lane25_strm0_cntl          ( std__pe55__lane25_strm0_cntl       ),      
               .std__pe55__lane25_strm0_data          ( std__pe55__lane25_strm0_data       ),      
               .std__pe55__lane25_strm0_data_valid    ( std__pe55__lane25_strm0_data_valid ),      
               .std__pe55__lane25_strm0_data_mask     ( std__pe55__lane25_strm0_data_mask  ),      

               .pe55__std__lane25_strm1_ready         ( pe55__std__lane25_strm1_ready      ),      
               .std__pe55__lane25_strm1_cntl          ( std__pe55__lane25_strm1_cntl       ),      
               .std__pe55__lane25_strm1_data          ( std__pe55__lane25_strm1_data       ),      
               .std__pe55__lane25_strm1_data_valid    ( std__pe55__lane25_strm1_data_valid ),      
               .std__pe55__lane25_strm1_data_mask     ( std__pe55__lane25_strm1_data_mask  ),      

               // PE 55, Lane 26                 
               .pe55__std__lane26_strm0_ready         ( pe55__std__lane26_strm0_ready      ),      
               .std__pe55__lane26_strm0_cntl          ( std__pe55__lane26_strm0_cntl       ),      
               .std__pe55__lane26_strm0_data          ( std__pe55__lane26_strm0_data       ),      
               .std__pe55__lane26_strm0_data_valid    ( std__pe55__lane26_strm0_data_valid ),      
               .std__pe55__lane26_strm0_data_mask     ( std__pe55__lane26_strm0_data_mask  ),      

               .pe55__std__lane26_strm1_ready         ( pe55__std__lane26_strm1_ready      ),      
               .std__pe55__lane26_strm1_cntl          ( std__pe55__lane26_strm1_cntl       ),      
               .std__pe55__lane26_strm1_data          ( std__pe55__lane26_strm1_data       ),      
               .std__pe55__lane26_strm1_data_valid    ( std__pe55__lane26_strm1_data_valid ),      
               .std__pe55__lane26_strm1_data_mask     ( std__pe55__lane26_strm1_data_mask  ),      

               // PE 55, Lane 27                 
               .pe55__std__lane27_strm0_ready         ( pe55__std__lane27_strm0_ready      ),      
               .std__pe55__lane27_strm0_cntl          ( std__pe55__lane27_strm0_cntl       ),      
               .std__pe55__lane27_strm0_data          ( std__pe55__lane27_strm0_data       ),      
               .std__pe55__lane27_strm0_data_valid    ( std__pe55__lane27_strm0_data_valid ),      
               .std__pe55__lane27_strm0_data_mask     ( std__pe55__lane27_strm0_data_mask  ),      

               .pe55__std__lane27_strm1_ready         ( pe55__std__lane27_strm1_ready      ),      
               .std__pe55__lane27_strm1_cntl          ( std__pe55__lane27_strm1_cntl       ),      
               .std__pe55__lane27_strm1_data          ( std__pe55__lane27_strm1_data       ),      
               .std__pe55__lane27_strm1_data_valid    ( std__pe55__lane27_strm1_data_valid ),      
               .std__pe55__lane27_strm1_data_mask     ( std__pe55__lane27_strm1_data_mask  ),      

               // PE 55, Lane 28                 
               .pe55__std__lane28_strm0_ready         ( pe55__std__lane28_strm0_ready      ),      
               .std__pe55__lane28_strm0_cntl          ( std__pe55__lane28_strm0_cntl       ),      
               .std__pe55__lane28_strm0_data          ( std__pe55__lane28_strm0_data       ),      
               .std__pe55__lane28_strm0_data_valid    ( std__pe55__lane28_strm0_data_valid ),      
               .std__pe55__lane28_strm0_data_mask     ( std__pe55__lane28_strm0_data_mask  ),      

               .pe55__std__lane28_strm1_ready         ( pe55__std__lane28_strm1_ready      ),      
               .std__pe55__lane28_strm1_cntl          ( std__pe55__lane28_strm1_cntl       ),      
               .std__pe55__lane28_strm1_data          ( std__pe55__lane28_strm1_data       ),      
               .std__pe55__lane28_strm1_data_valid    ( std__pe55__lane28_strm1_data_valid ),      
               .std__pe55__lane28_strm1_data_mask     ( std__pe55__lane28_strm1_data_mask  ),      

               // PE 55, Lane 29                 
               .pe55__std__lane29_strm0_ready         ( pe55__std__lane29_strm0_ready      ),      
               .std__pe55__lane29_strm0_cntl          ( std__pe55__lane29_strm0_cntl       ),      
               .std__pe55__lane29_strm0_data          ( std__pe55__lane29_strm0_data       ),      
               .std__pe55__lane29_strm0_data_valid    ( std__pe55__lane29_strm0_data_valid ),      
               .std__pe55__lane29_strm0_data_mask     ( std__pe55__lane29_strm0_data_mask  ),      

               .pe55__std__lane29_strm1_ready         ( pe55__std__lane29_strm1_ready      ),      
               .std__pe55__lane29_strm1_cntl          ( std__pe55__lane29_strm1_cntl       ),      
               .std__pe55__lane29_strm1_data          ( std__pe55__lane29_strm1_data       ),      
               .std__pe55__lane29_strm1_data_valid    ( std__pe55__lane29_strm1_data_valid ),      
               .std__pe55__lane29_strm1_data_mask     ( std__pe55__lane29_strm1_data_mask  ),      

               // PE 55, Lane 30                 
               .pe55__std__lane30_strm0_ready         ( pe55__std__lane30_strm0_ready      ),      
               .std__pe55__lane30_strm0_cntl          ( std__pe55__lane30_strm0_cntl       ),      
               .std__pe55__lane30_strm0_data          ( std__pe55__lane30_strm0_data       ),      
               .std__pe55__lane30_strm0_data_valid    ( std__pe55__lane30_strm0_data_valid ),      
               .std__pe55__lane30_strm0_data_mask     ( std__pe55__lane30_strm0_data_mask  ),      

               .pe55__std__lane30_strm1_ready         ( pe55__std__lane30_strm1_ready      ),      
               .std__pe55__lane30_strm1_cntl          ( std__pe55__lane30_strm1_cntl       ),      
               .std__pe55__lane30_strm1_data          ( std__pe55__lane30_strm1_data       ),      
               .std__pe55__lane30_strm1_data_valid    ( std__pe55__lane30_strm1_data_valid ),      
               .std__pe55__lane30_strm1_data_mask     ( std__pe55__lane30_strm1_data_mask  ),      

               // PE 55, Lane 31                 
               .pe55__std__lane31_strm0_ready         ( pe55__std__lane31_strm0_ready      ),      
               .std__pe55__lane31_strm0_cntl          ( std__pe55__lane31_strm0_cntl       ),      
               .std__pe55__lane31_strm0_data          ( std__pe55__lane31_strm0_data       ),      
               .std__pe55__lane31_strm0_data_valid    ( std__pe55__lane31_strm0_data_valid ),      
               .std__pe55__lane31_strm0_data_mask     ( std__pe55__lane31_strm0_data_mask  ),      

               .pe55__std__lane31_strm1_ready         ( pe55__std__lane31_strm1_ready      ),      
               .std__pe55__lane31_strm1_cntl          ( std__pe55__lane31_strm1_cntl       ),      
               .std__pe55__lane31_strm1_data          ( std__pe55__lane31_strm1_data       ),      
               .std__pe55__lane31_strm1_data_valid    ( std__pe55__lane31_strm1_data_valid ),      
               .std__pe55__lane31_strm1_data_mask     ( std__pe55__lane31_strm1_data_mask  ),      

               // PE 56, Lane 0                 
               .pe56__std__lane0_strm0_ready         ( pe56__std__lane0_strm0_ready      ),      
               .std__pe56__lane0_strm0_cntl          ( std__pe56__lane0_strm0_cntl       ),      
               .std__pe56__lane0_strm0_data          ( std__pe56__lane0_strm0_data       ),      
               .std__pe56__lane0_strm0_data_valid    ( std__pe56__lane0_strm0_data_valid ),      
               .std__pe56__lane0_strm0_data_mask     ( std__pe56__lane0_strm0_data_mask  ),      

               .pe56__std__lane0_strm1_ready         ( pe56__std__lane0_strm1_ready      ),      
               .std__pe56__lane0_strm1_cntl          ( std__pe56__lane0_strm1_cntl       ),      
               .std__pe56__lane0_strm1_data          ( std__pe56__lane0_strm1_data       ),      
               .std__pe56__lane0_strm1_data_valid    ( std__pe56__lane0_strm1_data_valid ),      
               .std__pe56__lane0_strm1_data_mask     ( std__pe56__lane0_strm1_data_mask  ),      

               // PE 56, Lane 1                 
               .pe56__std__lane1_strm0_ready         ( pe56__std__lane1_strm0_ready      ),      
               .std__pe56__lane1_strm0_cntl          ( std__pe56__lane1_strm0_cntl       ),      
               .std__pe56__lane1_strm0_data          ( std__pe56__lane1_strm0_data       ),      
               .std__pe56__lane1_strm0_data_valid    ( std__pe56__lane1_strm0_data_valid ),      
               .std__pe56__lane1_strm0_data_mask     ( std__pe56__lane1_strm0_data_mask  ),      

               .pe56__std__lane1_strm1_ready         ( pe56__std__lane1_strm1_ready      ),      
               .std__pe56__lane1_strm1_cntl          ( std__pe56__lane1_strm1_cntl       ),      
               .std__pe56__lane1_strm1_data          ( std__pe56__lane1_strm1_data       ),      
               .std__pe56__lane1_strm1_data_valid    ( std__pe56__lane1_strm1_data_valid ),      
               .std__pe56__lane1_strm1_data_mask     ( std__pe56__lane1_strm1_data_mask  ),      

               // PE 56, Lane 2                 
               .pe56__std__lane2_strm0_ready         ( pe56__std__lane2_strm0_ready      ),      
               .std__pe56__lane2_strm0_cntl          ( std__pe56__lane2_strm0_cntl       ),      
               .std__pe56__lane2_strm0_data          ( std__pe56__lane2_strm0_data       ),      
               .std__pe56__lane2_strm0_data_valid    ( std__pe56__lane2_strm0_data_valid ),      
               .std__pe56__lane2_strm0_data_mask     ( std__pe56__lane2_strm0_data_mask  ),      

               .pe56__std__lane2_strm1_ready         ( pe56__std__lane2_strm1_ready      ),      
               .std__pe56__lane2_strm1_cntl          ( std__pe56__lane2_strm1_cntl       ),      
               .std__pe56__lane2_strm1_data          ( std__pe56__lane2_strm1_data       ),      
               .std__pe56__lane2_strm1_data_valid    ( std__pe56__lane2_strm1_data_valid ),      
               .std__pe56__lane2_strm1_data_mask     ( std__pe56__lane2_strm1_data_mask  ),      

               // PE 56, Lane 3                 
               .pe56__std__lane3_strm0_ready         ( pe56__std__lane3_strm0_ready      ),      
               .std__pe56__lane3_strm0_cntl          ( std__pe56__lane3_strm0_cntl       ),      
               .std__pe56__lane3_strm0_data          ( std__pe56__lane3_strm0_data       ),      
               .std__pe56__lane3_strm0_data_valid    ( std__pe56__lane3_strm0_data_valid ),      
               .std__pe56__lane3_strm0_data_mask     ( std__pe56__lane3_strm0_data_mask  ),      

               .pe56__std__lane3_strm1_ready         ( pe56__std__lane3_strm1_ready      ),      
               .std__pe56__lane3_strm1_cntl          ( std__pe56__lane3_strm1_cntl       ),      
               .std__pe56__lane3_strm1_data          ( std__pe56__lane3_strm1_data       ),      
               .std__pe56__lane3_strm1_data_valid    ( std__pe56__lane3_strm1_data_valid ),      
               .std__pe56__lane3_strm1_data_mask     ( std__pe56__lane3_strm1_data_mask  ),      

               // PE 56, Lane 4                 
               .pe56__std__lane4_strm0_ready         ( pe56__std__lane4_strm0_ready      ),      
               .std__pe56__lane4_strm0_cntl          ( std__pe56__lane4_strm0_cntl       ),      
               .std__pe56__lane4_strm0_data          ( std__pe56__lane4_strm0_data       ),      
               .std__pe56__lane4_strm0_data_valid    ( std__pe56__lane4_strm0_data_valid ),      
               .std__pe56__lane4_strm0_data_mask     ( std__pe56__lane4_strm0_data_mask  ),      

               .pe56__std__lane4_strm1_ready         ( pe56__std__lane4_strm1_ready      ),      
               .std__pe56__lane4_strm1_cntl          ( std__pe56__lane4_strm1_cntl       ),      
               .std__pe56__lane4_strm1_data          ( std__pe56__lane4_strm1_data       ),      
               .std__pe56__lane4_strm1_data_valid    ( std__pe56__lane4_strm1_data_valid ),      
               .std__pe56__lane4_strm1_data_mask     ( std__pe56__lane4_strm1_data_mask  ),      

               // PE 56, Lane 5                 
               .pe56__std__lane5_strm0_ready         ( pe56__std__lane5_strm0_ready      ),      
               .std__pe56__lane5_strm0_cntl          ( std__pe56__lane5_strm0_cntl       ),      
               .std__pe56__lane5_strm0_data          ( std__pe56__lane5_strm0_data       ),      
               .std__pe56__lane5_strm0_data_valid    ( std__pe56__lane5_strm0_data_valid ),      
               .std__pe56__lane5_strm0_data_mask     ( std__pe56__lane5_strm0_data_mask  ),      

               .pe56__std__lane5_strm1_ready         ( pe56__std__lane5_strm1_ready      ),      
               .std__pe56__lane5_strm1_cntl          ( std__pe56__lane5_strm1_cntl       ),      
               .std__pe56__lane5_strm1_data          ( std__pe56__lane5_strm1_data       ),      
               .std__pe56__lane5_strm1_data_valid    ( std__pe56__lane5_strm1_data_valid ),      
               .std__pe56__lane5_strm1_data_mask     ( std__pe56__lane5_strm1_data_mask  ),      

               // PE 56, Lane 6                 
               .pe56__std__lane6_strm0_ready         ( pe56__std__lane6_strm0_ready      ),      
               .std__pe56__lane6_strm0_cntl          ( std__pe56__lane6_strm0_cntl       ),      
               .std__pe56__lane6_strm0_data          ( std__pe56__lane6_strm0_data       ),      
               .std__pe56__lane6_strm0_data_valid    ( std__pe56__lane6_strm0_data_valid ),      
               .std__pe56__lane6_strm0_data_mask     ( std__pe56__lane6_strm0_data_mask  ),      

               .pe56__std__lane6_strm1_ready         ( pe56__std__lane6_strm1_ready      ),      
               .std__pe56__lane6_strm1_cntl          ( std__pe56__lane6_strm1_cntl       ),      
               .std__pe56__lane6_strm1_data          ( std__pe56__lane6_strm1_data       ),      
               .std__pe56__lane6_strm1_data_valid    ( std__pe56__lane6_strm1_data_valid ),      
               .std__pe56__lane6_strm1_data_mask     ( std__pe56__lane6_strm1_data_mask  ),      

               // PE 56, Lane 7                 
               .pe56__std__lane7_strm0_ready         ( pe56__std__lane7_strm0_ready      ),      
               .std__pe56__lane7_strm0_cntl          ( std__pe56__lane7_strm0_cntl       ),      
               .std__pe56__lane7_strm0_data          ( std__pe56__lane7_strm0_data       ),      
               .std__pe56__lane7_strm0_data_valid    ( std__pe56__lane7_strm0_data_valid ),      
               .std__pe56__lane7_strm0_data_mask     ( std__pe56__lane7_strm0_data_mask  ),      

               .pe56__std__lane7_strm1_ready         ( pe56__std__lane7_strm1_ready      ),      
               .std__pe56__lane7_strm1_cntl          ( std__pe56__lane7_strm1_cntl       ),      
               .std__pe56__lane7_strm1_data          ( std__pe56__lane7_strm1_data       ),      
               .std__pe56__lane7_strm1_data_valid    ( std__pe56__lane7_strm1_data_valid ),      
               .std__pe56__lane7_strm1_data_mask     ( std__pe56__lane7_strm1_data_mask  ),      

               // PE 56, Lane 8                 
               .pe56__std__lane8_strm0_ready         ( pe56__std__lane8_strm0_ready      ),      
               .std__pe56__lane8_strm0_cntl          ( std__pe56__lane8_strm0_cntl       ),      
               .std__pe56__lane8_strm0_data          ( std__pe56__lane8_strm0_data       ),      
               .std__pe56__lane8_strm0_data_valid    ( std__pe56__lane8_strm0_data_valid ),      
               .std__pe56__lane8_strm0_data_mask     ( std__pe56__lane8_strm0_data_mask  ),      

               .pe56__std__lane8_strm1_ready         ( pe56__std__lane8_strm1_ready      ),      
               .std__pe56__lane8_strm1_cntl          ( std__pe56__lane8_strm1_cntl       ),      
               .std__pe56__lane8_strm1_data          ( std__pe56__lane8_strm1_data       ),      
               .std__pe56__lane8_strm1_data_valid    ( std__pe56__lane8_strm1_data_valid ),      
               .std__pe56__lane8_strm1_data_mask     ( std__pe56__lane8_strm1_data_mask  ),      

               // PE 56, Lane 9                 
               .pe56__std__lane9_strm0_ready         ( pe56__std__lane9_strm0_ready      ),      
               .std__pe56__lane9_strm0_cntl          ( std__pe56__lane9_strm0_cntl       ),      
               .std__pe56__lane9_strm0_data          ( std__pe56__lane9_strm0_data       ),      
               .std__pe56__lane9_strm0_data_valid    ( std__pe56__lane9_strm0_data_valid ),      
               .std__pe56__lane9_strm0_data_mask     ( std__pe56__lane9_strm0_data_mask  ),      

               .pe56__std__lane9_strm1_ready         ( pe56__std__lane9_strm1_ready      ),      
               .std__pe56__lane9_strm1_cntl          ( std__pe56__lane9_strm1_cntl       ),      
               .std__pe56__lane9_strm1_data          ( std__pe56__lane9_strm1_data       ),      
               .std__pe56__lane9_strm1_data_valid    ( std__pe56__lane9_strm1_data_valid ),      
               .std__pe56__lane9_strm1_data_mask     ( std__pe56__lane9_strm1_data_mask  ),      

               // PE 56, Lane 10                 
               .pe56__std__lane10_strm0_ready         ( pe56__std__lane10_strm0_ready      ),      
               .std__pe56__lane10_strm0_cntl          ( std__pe56__lane10_strm0_cntl       ),      
               .std__pe56__lane10_strm0_data          ( std__pe56__lane10_strm0_data       ),      
               .std__pe56__lane10_strm0_data_valid    ( std__pe56__lane10_strm0_data_valid ),      
               .std__pe56__lane10_strm0_data_mask     ( std__pe56__lane10_strm0_data_mask  ),      

               .pe56__std__lane10_strm1_ready         ( pe56__std__lane10_strm1_ready      ),      
               .std__pe56__lane10_strm1_cntl          ( std__pe56__lane10_strm1_cntl       ),      
               .std__pe56__lane10_strm1_data          ( std__pe56__lane10_strm1_data       ),      
               .std__pe56__lane10_strm1_data_valid    ( std__pe56__lane10_strm1_data_valid ),      
               .std__pe56__lane10_strm1_data_mask     ( std__pe56__lane10_strm1_data_mask  ),      

               // PE 56, Lane 11                 
               .pe56__std__lane11_strm0_ready         ( pe56__std__lane11_strm0_ready      ),      
               .std__pe56__lane11_strm0_cntl          ( std__pe56__lane11_strm0_cntl       ),      
               .std__pe56__lane11_strm0_data          ( std__pe56__lane11_strm0_data       ),      
               .std__pe56__lane11_strm0_data_valid    ( std__pe56__lane11_strm0_data_valid ),      
               .std__pe56__lane11_strm0_data_mask     ( std__pe56__lane11_strm0_data_mask  ),      

               .pe56__std__lane11_strm1_ready         ( pe56__std__lane11_strm1_ready      ),      
               .std__pe56__lane11_strm1_cntl          ( std__pe56__lane11_strm1_cntl       ),      
               .std__pe56__lane11_strm1_data          ( std__pe56__lane11_strm1_data       ),      
               .std__pe56__lane11_strm1_data_valid    ( std__pe56__lane11_strm1_data_valid ),      
               .std__pe56__lane11_strm1_data_mask     ( std__pe56__lane11_strm1_data_mask  ),      

               // PE 56, Lane 12                 
               .pe56__std__lane12_strm0_ready         ( pe56__std__lane12_strm0_ready      ),      
               .std__pe56__lane12_strm0_cntl          ( std__pe56__lane12_strm0_cntl       ),      
               .std__pe56__lane12_strm0_data          ( std__pe56__lane12_strm0_data       ),      
               .std__pe56__lane12_strm0_data_valid    ( std__pe56__lane12_strm0_data_valid ),      
               .std__pe56__lane12_strm0_data_mask     ( std__pe56__lane12_strm0_data_mask  ),      

               .pe56__std__lane12_strm1_ready         ( pe56__std__lane12_strm1_ready      ),      
               .std__pe56__lane12_strm1_cntl          ( std__pe56__lane12_strm1_cntl       ),      
               .std__pe56__lane12_strm1_data          ( std__pe56__lane12_strm1_data       ),      
               .std__pe56__lane12_strm1_data_valid    ( std__pe56__lane12_strm1_data_valid ),      
               .std__pe56__lane12_strm1_data_mask     ( std__pe56__lane12_strm1_data_mask  ),      

               // PE 56, Lane 13                 
               .pe56__std__lane13_strm0_ready         ( pe56__std__lane13_strm0_ready      ),      
               .std__pe56__lane13_strm0_cntl          ( std__pe56__lane13_strm0_cntl       ),      
               .std__pe56__lane13_strm0_data          ( std__pe56__lane13_strm0_data       ),      
               .std__pe56__lane13_strm0_data_valid    ( std__pe56__lane13_strm0_data_valid ),      
               .std__pe56__lane13_strm0_data_mask     ( std__pe56__lane13_strm0_data_mask  ),      

               .pe56__std__lane13_strm1_ready         ( pe56__std__lane13_strm1_ready      ),      
               .std__pe56__lane13_strm1_cntl          ( std__pe56__lane13_strm1_cntl       ),      
               .std__pe56__lane13_strm1_data          ( std__pe56__lane13_strm1_data       ),      
               .std__pe56__lane13_strm1_data_valid    ( std__pe56__lane13_strm1_data_valid ),      
               .std__pe56__lane13_strm1_data_mask     ( std__pe56__lane13_strm1_data_mask  ),      

               // PE 56, Lane 14                 
               .pe56__std__lane14_strm0_ready         ( pe56__std__lane14_strm0_ready      ),      
               .std__pe56__lane14_strm0_cntl          ( std__pe56__lane14_strm0_cntl       ),      
               .std__pe56__lane14_strm0_data          ( std__pe56__lane14_strm0_data       ),      
               .std__pe56__lane14_strm0_data_valid    ( std__pe56__lane14_strm0_data_valid ),      
               .std__pe56__lane14_strm0_data_mask     ( std__pe56__lane14_strm0_data_mask  ),      

               .pe56__std__lane14_strm1_ready         ( pe56__std__lane14_strm1_ready      ),      
               .std__pe56__lane14_strm1_cntl          ( std__pe56__lane14_strm1_cntl       ),      
               .std__pe56__lane14_strm1_data          ( std__pe56__lane14_strm1_data       ),      
               .std__pe56__lane14_strm1_data_valid    ( std__pe56__lane14_strm1_data_valid ),      
               .std__pe56__lane14_strm1_data_mask     ( std__pe56__lane14_strm1_data_mask  ),      

               // PE 56, Lane 15                 
               .pe56__std__lane15_strm0_ready         ( pe56__std__lane15_strm0_ready      ),      
               .std__pe56__lane15_strm0_cntl          ( std__pe56__lane15_strm0_cntl       ),      
               .std__pe56__lane15_strm0_data          ( std__pe56__lane15_strm0_data       ),      
               .std__pe56__lane15_strm0_data_valid    ( std__pe56__lane15_strm0_data_valid ),      
               .std__pe56__lane15_strm0_data_mask     ( std__pe56__lane15_strm0_data_mask  ),      

               .pe56__std__lane15_strm1_ready         ( pe56__std__lane15_strm1_ready      ),      
               .std__pe56__lane15_strm1_cntl          ( std__pe56__lane15_strm1_cntl       ),      
               .std__pe56__lane15_strm1_data          ( std__pe56__lane15_strm1_data       ),      
               .std__pe56__lane15_strm1_data_valid    ( std__pe56__lane15_strm1_data_valid ),      
               .std__pe56__lane15_strm1_data_mask     ( std__pe56__lane15_strm1_data_mask  ),      

               // PE 56, Lane 16                 
               .pe56__std__lane16_strm0_ready         ( pe56__std__lane16_strm0_ready      ),      
               .std__pe56__lane16_strm0_cntl          ( std__pe56__lane16_strm0_cntl       ),      
               .std__pe56__lane16_strm0_data          ( std__pe56__lane16_strm0_data       ),      
               .std__pe56__lane16_strm0_data_valid    ( std__pe56__lane16_strm0_data_valid ),      
               .std__pe56__lane16_strm0_data_mask     ( std__pe56__lane16_strm0_data_mask  ),      

               .pe56__std__lane16_strm1_ready         ( pe56__std__lane16_strm1_ready      ),      
               .std__pe56__lane16_strm1_cntl          ( std__pe56__lane16_strm1_cntl       ),      
               .std__pe56__lane16_strm1_data          ( std__pe56__lane16_strm1_data       ),      
               .std__pe56__lane16_strm1_data_valid    ( std__pe56__lane16_strm1_data_valid ),      
               .std__pe56__lane16_strm1_data_mask     ( std__pe56__lane16_strm1_data_mask  ),      

               // PE 56, Lane 17                 
               .pe56__std__lane17_strm0_ready         ( pe56__std__lane17_strm0_ready      ),      
               .std__pe56__lane17_strm0_cntl          ( std__pe56__lane17_strm0_cntl       ),      
               .std__pe56__lane17_strm0_data          ( std__pe56__lane17_strm0_data       ),      
               .std__pe56__lane17_strm0_data_valid    ( std__pe56__lane17_strm0_data_valid ),      
               .std__pe56__lane17_strm0_data_mask     ( std__pe56__lane17_strm0_data_mask  ),      

               .pe56__std__lane17_strm1_ready         ( pe56__std__lane17_strm1_ready      ),      
               .std__pe56__lane17_strm1_cntl          ( std__pe56__lane17_strm1_cntl       ),      
               .std__pe56__lane17_strm1_data          ( std__pe56__lane17_strm1_data       ),      
               .std__pe56__lane17_strm1_data_valid    ( std__pe56__lane17_strm1_data_valid ),      
               .std__pe56__lane17_strm1_data_mask     ( std__pe56__lane17_strm1_data_mask  ),      

               // PE 56, Lane 18                 
               .pe56__std__lane18_strm0_ready         ( pe56__std__lane18_strm0_ready      ),      
               .std__pe56__lane18_strm0_cntl          ( std__pe56__lane18_strm0_cntl       ),      
               .std__pe56__lane18_strm0_data          ( std__pe56__lane18_strm0_data       ),      
               .std__pe56__lane18_strm0_data_valid    ( std__pe56__lane18_strm0_data_valid ),      
               .std__pe56__lane18_strm0_data_mask     ( std__pe56__lane18_strm0_data_mask  ),      

               .pe56__std__lane18_strm1_ready         ( pe56__std__lane18_strm1_ready      ),      
               .std__pe56__lane18_strm1_cntl          ( std__pe56__lane18_strm1_cntl       ),      
               .std__pe56__lane18_strm1_data          ( std__pe56__lane18_strm1_data       ),      
               .std__pe56__lane18_strm1_data_valid    ( std__pe56__lane18_strm1_data_valid ),      
               .std__pe56__lane18_strm1_data_mask     ( std__pe56__lane18_strm1_data_mask  ),      

               // PE 56, Lane 19                 
               .pe56__std__lane19_strm0_ready         ( pe56__std__lane19_strm0_ready      ),      
               .std__pe56__lane19_strm0_cntl          ( std__pe56__lane19_strm0_cntl       ),      
               .std__pe56__lane19_strm0_data          ( std__pe56__lane19_strm0_data       ),      
               .std__pe56__lane19_strm0_data_valid    ( std__pe56__lane19_strm0_data_valid ),      
               .std__pe56__lane19_strm0_data_mask     ( std__pe56__lane19_strm0_data_mask  ),      

               .pe56__std__lane19_strm1_ready         ( pe56__std__lane19_strm1_ready      ),      
               .std__pe56__lane19_strm1_cntl          ( std__pe56__lane19_strm1_cntl       ),      
               .std__pe56__lane19_strm1_data          ( std__pe56__lane19_strm1_data       ),      
               .std__pe56__lane19_strm1_data_valid    ( std__pe56__lane19_strm1_data_valid ),      
               .std__pe56__lane19_strm1_data_mask     ( std__pe56__lane19_strm1_data_mask  ),      

               // PE 56, Lane 20                 
               .pe56__std__lane20_strm0_ready         ( pe56__std__lane20_strm0_ready      ),      
               .std__pe56__lane20_strm0_cntl          ( std__pe56__lane20_strm0_cntl       ),      
               .std__pe56__lane20_strm0_data          ( std__pe56__lane20_strm0_data       ),      
               .std__pe56__lane20_strm0_data_valid    ( std__pe56__lane20_strm0_data_valid ),      
               .std__pe56__lane20_strm0_data_mask     ( std__pe56__lane20_strm0_data_mask  ),      

               .pe56__std__lane20_strm1_ready         ( pe56__std__lane20_strm1_ready      ),      
               .std__pe56__lane20_strm1_cntl          ( std__pe56__lane20_strm1_cntl       ),      
               .std__pe56__lane20_strm1_data          ( std__pe56__lane20_strm1_data       ),      
               .std__pe56__lane20_strm1_data_valid    ( std__pe56__lane20_strm1_data_valid ),      
               .std__pe56__lane20_strm1_data_mask     ( std__pe56__lane20_strm1_data_mask  ),      

               // PE 56, Lane 21                 
               .pe56__std__lane21_strm0_ready         ( pe56__std__lane21_strm0_ready      ),      
               .std__pe56__lane21_strm0_cntl          ( std__pe56__lane21_strm0_cntl       ),      
               .std__pe56__lane21_strm0_data          ( std__pe56__lane21_strm0_data       ),      
               .std__pe56__lane21_strm0_data_valid    ( std__pe56__lane21_strm0_data_valid ),      
               .std__pe56__lane21_strm0_data_mask     ( std__pe56__lane21_strm0_data_mask  ),      

               .pe56__std__lane21_strm1_ready         ( pe56__std__lane21_strm1_ready      ),      
               .std__pe56__lane21_strm1_cntl          ( std__pe56__lane21_strm1_cntl       ),      
               .std__pe56__lane21_strm1_data          ( std__pe56__lane21_strm1_data       ),      
               .std__pe56__lane21_strm1_data_valid    ( std__pe56__lane21_strm1_data_valid ),      
               .std__pe56__lane21_strm1_data_mask     ( std__pe56__lane21_strm1_data_mask  ),      

               // PE 56, Lane 22                 
               .pe56__std__lane22_strm0_ready         ( pe56__std__lane22_strm0_ready      ),      
               .std__pe56__lane22_strm0_cntl          ( std__pe56__lane22_strm0_cntl       ),      
               .std__pe56__lane22_strm0_data          ( std__pe56__lane22_strm0_data       ),      
               .std__pe56__lane22_strm0_data_valid    ( std__pe56__lane22_strm0_data_valid ),      
               .std__pe56__lane22_strm0_data_mask     ( std__pe56__lane22_strm0_data_mask  ),      

               .pe56__std__lane22_strm1_ready         ( pe56__std__lane22_strm1_ready      ),      
               .std__pe56__lane22_strm1_cntl          ( std__pe56__lane22_strm1_cntl       ),      
               .std__pe56__lane22_strm1_data          ( std__pe56__lane22_strm1_data       ),      
               .std__pe56__lane22_strm1_data_valid    ( std__pe56__lane22_strm1_data_valid ),      
               .std__pe56__lane22_strm1_data_mask     ( std__pe56__lane22_strm1_data_mask  ),      

               // PE 56, Lane 23                 
               .pe56__std__lane23_strm0_ready         ( pe56__std__lane23_strm0_ready      ),      
               .std__pe56__lane23_strm0_cntl          ( std__pe56__lane23_strm0_cntl       ),      
               .std__pe56__lane23_strm0_data          ( std__pe56__lane23_strm0_data       ),      
               .std__pe56__lane23_strm0_data_valid    ( std__pe56__lane23_strm0_data_valid ),      
               .std__pe56__lane23_strm0_data_mask     ( std__pe56__lane23_strm0_data_mask  ),      

               .pe56__std__lane23_strm1_ready         ( pe56__std__lane23_strm1_ready      ),      
               .std__pe56__lane23_strm1_cntl          ( std__pe56__lane23_strm1_cntl       ),      
               .std__pe56__lane23_strm1_data          ( std__pe56__lane23_strm1_data       ),      
               .std__pe56__lane23_strm1_data_valid    ( std__pe56__lane23_strm1_data_valid ),      
               .std__pe56__lane23_strm1_data_mask     ( std__pe56__lane23_strm1_data_mask  ),      

               // PE 56, Lane 24                 
               .pe56__std__lane24_strm0_ready         ( pe56__std__lane24_strm0_ready      ),      
               .std__pe56__lane24_strm0_cntl          ( std__pe56__lane24_strm0_cntl       ),      
               .std__pe56__lane24_strm0_data          ( std__pe56__lane24_strm0_data       ),      
               .std__pe56__lane24_strm0_data_valid    ( std__pe56__lane24_strm0_data_valid ),      
               .std__pe56__lane24_strm0_data_mask     ( std__pe56__lane24_strm0_data_mask  ),      

               .pe56__std__lane24_strm1_ready         ( pe56__std__lane24_strm1_ready      ),      
               .std__pe56__lane24_strm1_cntl          ( std__pe56__lane24_strm1_cntl       ),      
               .std__pe56__lane24_strm1_data          ( std__pe56__lane24_strm1_data       ),      
               .std__pe56__lane24_strm1_data_valid    ( std__pe56__lane24_strm1_data_valid ),      
               .std__pe56__lane24_strm1_data_mask     ( std__pe56__lane24_strm1_data_mask  ),      

               // PE 56, Lane 25                 
               .pe56__std__lane25_strm0_ready         ( pe56__std__lane25_strm0_ready      ),      
               .std__pe56__lane25_strm0_cntl          ( std__pe56__lane25_strm0_cntl       ),      
               .std__pe56__lane25_strm0_data          ( std__pe56__lane25_strm0_data       ),      
               .std__pe56__lane25_strm0_data_valid    ( std__pe56__lane25_strm0_data_valid ),      
               .std__pe56__lane25_strm0_data_mask     ( std__pe56__lane25_strm0_data_mask  ),      

               .pe56__std__lane25_strm1_ready         ( pe56__std__lane25_strm1_ready      ),      
               .std__pe56__lane25_strm1_cntl          ( std__pe56__lane25_strm1_cntl       ),      
               .std__pe56__lane25_strm1_data          ( std__pe56__lane25_strm1_data       ),      
               .std__pe56__lane25_strm1_data_valid    ( std__pe56__lane25_strm1_data_valid ),      
               .std__pe56__lane25_strm1_data_mask     ( std__pe56__lane25_strm1_data_mask  ),      

               // PE 56, Lane 26                 
               .pe56__std__lane26_strm0_ready         ( pe56__std__lane26_strm0_ready      ),      
               .std__pe56__lane26_strm0_cntl          ( std__pe56__lane26_strm0_cntl       ),      
               .std__pe56__lane26_strm0_data          ( std__pe56__lane26_strm0_data       ),      
               .std__pe56__lane26_strm0_data_valid    ( std__pe56__lane26_strm0_data_valid ),      
               .std__pe56__lane26_strm0_data_mask     ( std__pe56__lane26_strm0_data_mask  ),      

               .pe56__std__lane26_strm1_ready         ( pe56__std__lane26_strm1_ready      ),      
               .std__pe56__lane26_strm1_cntl          ( std__pe56__lane26_strm1_cntl       ),      
               .std__pe56__lane26_strm1_data          ( std__pe56__lane26_strm1_data       ),      
               .std__pe56__lane26_strm1_data_valid    ( std__pe56__lane26_strm1_data_valid ),      
               .std__pe56__lane26_strm1_data_mask     ( std__pe56__lane26_strm1_data_mask  ),      

               // PE 56, Lane 27                 
               .pe56__std__lane27_strm0_ready         ( pe56__std__lane27_strm0_ready      ),      
               .std__pe56__lane27_strm0_cntl          ( std__pe56__lane27_strm0_cntl       ),      
               .std__pe56__lane27_strm0_data          ( std__pe56__lane27_strm0_data       ),      
               .std__pe56__lane27_strm0_data_valid    ( std__pe56__lane27_strm0_data_valid ),      
               .std__pe56__lane27_strm0_data_mask     ( std__pe56__lane27_strm0_data_mask  ),      

               .pe56__std__lane27_strm1_ready         ( pe56__std__lane27_strm1_ready      ),      
               .std__pe56__lane27_strm1_cntl          ( std__pe56__lane27_strm1_cntl       ),      
               .std__pe56__lane27_strm1_data          ( std__pe56__lane27_strm1_data       ),      
               .std__pe56__lane27_strm1_data_valid    ( std__pe56__lane27_strm1_data_valid ),      
               .std__pe56__lane27_strm1_data_mask     ( std__pe56__lane27_strm1_data_mask  ),      

               // PE 56, Lane 28                 
               .pe56__std__lane28_strm0_ready         ( pe56__std__lane28_strm0_ready      ),      
               .std__pe56__lane28_strm0_cntl          ( std__pe56__lane28_strm0_cntl       ),      
               .std__pe56__lane28_strm0_data          ( std__pe56__lane28_strm0_data       ),      
               .std__pe56__lane28_strm0_data_valid    ( std__pe56__lane28_strm0_data_valid ),      
               .std__pe56__lane28_strm0_data_mask     ( std__pe56__lane28_strm0_data_mask  ),      

               .pe56__std__lane28_strm1_ready         ( pe56__std__lane28_strm1_ready      ),      
               .std__pe56__lane28_strm1_cntl          ( std__pe56__lane28_strm1_cntl       ),      
               .std__pe56__lane28_strm1_data          ( std__pe56__lane28_strm1_data       ),      
               .std__pe56__lane28_strm1_data_valid    ( std__pe56__lane28_strm1_data_valid ),      
               .std__pe56__lane28_strm1_data_mask     ( std__pe56__lane28_strm1_data_mask  ),      

               // PE 56, Lane 29                 
               .pe56__std__lane29_strm0_ready         ( pe56__std__lane29_strm0_ready      ),      
               .std__pe56__lane29_strm0_cntl          ( std__pe56__lane29_strm0_cntl       ),      
               .std__pe56__lane29_strm0_data          ( std__pe56__lane29_strm0_data       ),      
               .std__pe56__lane29_strm0_data_valid    ( std__pe56__lane29_strm0_data_valid ),      
               .std__pe56__lane29_strm0_data_mask     ( std__pe56__lane29_strm0_data_mask  ),      

               .pe56__std__lane29_strm1_ready         ( pe56__std__lane29_strm1_ready      ),      
               .std__pe56__lane29_strm1_cntl          ( std__pe56__lane29_strm1_cntl       ),      
               .std__pe56__lane29_strm1_data          ( std__pe56__lane29_strm1_data       ),      
               .std__pe56__lane29_strm1_data_valid    ( std__pe56__lane29_strm1_data_valid ),      
               .std__pe56__lane29_strm1_data_mask     ( std__pe56__lane29_strm1_data_mask  ),      

               // PE 56, Lane 30                 
               .pe56__std__lane30_strm0_ready         ( pe56__std__lane30_strm0_ready      ),      
               .std__pe56__lane30_strm0_cntl          ( std__pe56__lane30_strm0_cntl       ),      
               .std__pe56__lane30_strm0_data          ( std__pe56__lane30_strm0_data       ),      
               .std__pe56__lane30_strm0_data_valid    ( std__pe56__lane30_strm0_data_valid ),      
               .std__pe56__lane30_strm0_data_mask     ( std__pe56__lane30_strm0_data_mask  ),      

               .pe56__std__lane30_strm1_ready         ( pe56__std__lane30_strm1_ready      ),      
               .std__pe56__lane30_strm1_cntl          ( std__pe56__lane30_strm1_cntl       ),      
               .std__pe56__lane30_strm1_data          ( std__pe56__lane30_strm1_data       ),      
               .std__pe56__lane30_strm1_data_valid    ( std__pe56__lane30_strm1_data_valid ),      
               .std__pe56__lane30_strm1_data_mask     ( std__pe56__lane30_strm1_data_mask  ),      

               // PE 56, Lane 31                 
               .pe56__std__lane31_strm0_ready         ( pe56__std__lane31_strm0_ready      ),      
               .std__pe56__lane31_strm0_cntl          ( std__pe56__lane31_strm0_cntl       ),      
               .std__pe56__lane31_strm0_data          ( std__pe56__lane31_strm0_data       ),      
               .std__pe56__lane31_strm0_data_valid    ( std__pe56__lane31_strm0_data_valid ),      
               .std__pe56__lane31_strm0_data_mask     ( std__pe56__lane31_strm0_data_mask  ),      

               .pe56__std__lane31_strm1_ready         ( pe56__std__lane31_strm1_ready      ),      
               .std__pe56__lane31_strm1_cntl          ( std__pe56__lane31_strm1_cntl       ),      
               .std__pe56__lane31_strm1_data          ( std__pe56__lane31_strm1_data       ),      
               .std__pe56__lane31_strm1_data_valid    ( std__pe56__lane31_strm1_data_valid ),      
               .std__pe56__lane31_strm1_data_mask     ( std__pe56__lane31_strm1_data_mask  ),      

               // PE 57, Lane 0                 
               .pe57__std__lane0_strm0_ready         ( pe57__std__lane0_strm0_ready      ),      
               .std__pe57__lane0_strm0_cntl          ( std__pe57__lane0_strm0_cntl       ),      
               .std__pe57__lane0_strm0_data          ( std__pe57__lane0_strm0_data       ),      
               .std__pe57__lane0_strm0_data_valid    ( std__pe57__lane0_strm0_data_valid ),      
               .std__pe57__lane0_strm0_data_mask     ( std__pe57__lane0_strm0_data_mask  ),      

               .pe57__std__lane0_strm1_ready         ( pe57__std__lane0_strm1_ready      ),      
               .std__pe57__lane0_strm1_cntl          ( std__pe57__lane0_strm1_cntl       ),      
               .std__pe57__lane0_strm1_data          ( std__pe57__lane0_strm1_data       ),      
               .std__pe57__lane0_strm1_data_valid    ( std__pe57__lane0_strm1_data_valid ),      
               .std__pe57__lane0_strm1_data_mask     ( std__pe57__lane0_strm1_data_mask  ),      

               // PE 57, Lane 1                 
               .pe57__std__lane1_strm0_ready         ( pe57__std__lane1_strm0_ready      ),      
               .std__pe57__lane1_strm0_cntl          ( std__pe57__lane1_strm0_cntl       ),      
               .std__pe57__lane1_strm0_data          ( std__pe57__lane1_strm0_data       ),      
               .std__pe57__lane1_strm0_data_valid    ( std__pe57__lane1_strm0_data_valid ),      
               .std__pe57__lane1_strm0_data_mask     ( std__pe57__lane1_strm0_data_mask  ),      

               .pe57__std__lane1_strm1_ready         ( pe57__std__lane1_strm1_ready      ),      
               .std__pe57__lane1_strm1_cntl          ( std__pe57__lane1_strm1_cntl       ),      
               .std__pe57__lane1_strm1_data          ( std__pe57__lane1_strm1_data       ),      
               .std__pe57__lane1_strm1_data_valid    ( std__pe57__lane1_strm1_data_valid ),      
               .std__pe57__lane1_strm1_data_mask     ( std__pe57__lane1_strm1_data_mask  ),      

               // PE 57, Lane 2                 
               .pe57__std__lane2_strm0_ready         ( pe57__std__lane2_strm0_ready      ),      
               .std__pe57__lane2_strm0_cntl          ( std__pe57__lane2_strm0_cntl       ),      
               .std__pe57__lane2_strm0_data          ( std__pe57__lane2_strm0_data       ),      
               .std__pe57__lane2_strm0_data_valid    ( std__pe57__lane2_strm0_data_valid ),      
               .std__pe57__lane2_strm0_data_mask     ( std__pe57__lane2_strm0_data_mask  ),      

               .pe57__std__lane2_strm1_ready         ( pe57__std__lane2_strm1_ready      ),      
               .std__pe57__lane2_strm1_cntl          ( std__pe57__lane2_strm1_cntl       ),      
               .std__pe57__lane2_strm1_data          ( std__pe57__lane2_strm1_data       ),      
               .std__pe57__lane2_strm1_data_valid    ( std__pe57__lane2_strm1_data_valid ),      
               .std__pe57__lane2_strm1_data_mask     ( std__pe57__lane2_strm1_data_mask  ),      

               // PE 57, Lane 3                 
               .pe57__std__lane3_strm0_ready         ( pe57__std__lane3_strm0_ready      ),      
               .std__pe57__lane3_strm0_cntl          ( std__pe57__lane3_strm0_cntl       ),      
               .std__pe57__lane3_strm0_data          ( std__pe57__lane3_strm0_data       ),      
               .std__pe57__lane3_strm0_data_valid    ( std__pe57__lane3_strm0_data_valid ),      
               .std__pe57__lane3_strm0_data_mask     ( std__pe57__lane3_strm0_data_mask  ),      

               .pe57__std__lane3_strm1_ready         ( pe57__std__lane3_strm1_ready      ),      
               .std__pe57__lane3_strm1_cntl          ( std__pe57__lane3_strm1_cntl       ),      
               .std__pe57__lane3_strm1_data          ( std__pe57__lane3_strm1_data       ),      
               .std__pe57__lane3_strm1_data_valid    ( std__pe57__lane3_strm1_data_valid ),      
               .std__pe57__lane3_strm1_data_mask     ( std__pe57__lane3_strm1_data_mask  ),      

               // PE 57, Lane 4                 
               .pe57__std__lane4_strm0_ready         ( pe57__std__lane4_strm0_ready      ),      
               .std__pe57__lane4_strm0_cntl          ( std__pe57__lane4_strm0_cntl       ),      
               .std__pe57__lane4_strm0_data          ( std__pe57__lane4_strm0_data       ),      
               .std__pe57__lane4_strm0_data_valid    ( std__pe57__lane4_strm0_data_valid ),      
               .std__pe57__lane4_strm0_data_mask     ( std__pe57__lane4_strm0_data_mask  ),      

               .pe57__std__lane4_strm1_ready         ( pe57__std__lane4_strm1_ready      ),      
               .std__pe57__lane4_strm1_cntl          ( std__pe57__lane4_strm1_cntl       ),      
               .std__pe57__lane4_strm1_data          ( std__pe57__lane4_strm1_data       ),      
               .std__pe57__lane4_strm1_data_valid    ( std__pe57__lane4_strm1_data_valid ),      
               .std__pe57__lane4_strm1_data_mask     ( std__pe57__lane4_strm1_data_mask  ),      

               // PE 57, Lane 5                 
               .pe57__std__lane5_strm0_ready         ( pe57__std__lane5_strm0_ready      ),      
               .std__pe57__lane5_strm0_cntl          ( std__pe57__lane5_strm0_cntl       ),      
               .std__pe57__lane5_strm0_data          ( std__pe57__lane5_strm0_data       ),      
               .std__pe57__lane5_strm0_data_valid    ( std__pe57__lane5_strm0_data_valid ),      
               .std__pe57__lane5_strm0_data_mask     ( std__pe57__lane5_strm0_data_mask  ),      

               .pe57__std__lane5_strm1_ready         ( pe57__std__lane5_strm1_ready      ),      
               .std__pe57__lane5_strm1_cntl          ( std__pe57__lane5_strm1_cntl       ),      
               .std__pe57__lane5_strm1_data          ( std__pe57__lane5_strm1_data       ),      
               .std__pe57__lane5_strm1_data_valid    ( std__pe57__lane5_strm1_data_valid ),      
               .std__pe57__lane5_strm1_data_mask     ( std__pe57__lane5_strm1_data_mask  ),      

               // PE 57, Lane 6                 
               .pe57__std__lane6_strm0_ready         ( pe57__std__lane6_strm0_ready      ),      
               .std__pe57__lane6_strm0_cntl          ( std__pe57__lane6_strm0_cntl       ),      
               .std__pe57__lane6_strm0_data          ( std__pe57__lane6_strm0_data       ),      
               .std__pe57__lane6_strm0_data_valid    ( std__pe57__lane6_strm0_data_valid ),      
               .std__pe57__lane6_strm0_data_mask     ( std__pe57__lane6_strm0_data_mask  ),      

               .pe57__std__lane6_strm1_ready         ( pe57__std__lane6_strm1_ready      ),      
               .std__pe57__lane6_strm1_cntl          ( std__pe57__lane6_strm1_cntl       ),      
               .std__pe57__lane6_strm1_data          ( std__pe57__lane6_strm1_data       ),      
               .std__pe57__lane6_strm1_data_valid    ( std__pe57__lane6_strm1_data_valid ),      
               .std__pe57__lane6_strm1_data_mask     ( std__pe57__lane6_strm1_data_mask  ),      

               // PE 57, Lane 7                 
               .pe57__std__lane7_strm0_ready         ( pe57__std__lane7_strm0_ready      ),      
               .std__pe57__lane7_strm0_cntl          ( std__pe57__lane7_strm0_cntl       ),      
               .std__pe57__lane7_strm0_data          ( std__pe57__lane7_strm0_data       ),      
               .std__pe57__lane7_strm0_data_valid    ( std__pe57__lane7_strm0_data_valid ),      
               .std__pe57__lane7_strm0_data_mask     ( std__pe57__lane7_strm0_data_mask  ),      

               .pe57__std__lane7_strm1_ready         ( pe57__std__lane7_strm1_ready      ),      
               .std__pe57__lane7_strm1_cntl          ( std__pe57__lane7_strm1_cntl       ),      
               .std__pe57__lane7_strm1_data          ( std__pe57__lane7_strm1_data       ),      
               .std__pe57__lane7_strm1_data_valid    ( std__pe57__lane7_strm1_data_valid ),      
               .std__pe57__lane7_strm1_data_mask     ( std__pe57__lane7_strm1_data_mask  ),      

               // PE 57, Lane 8                 
               .pe57__std__lane8_strm0_ready         ( pe57__std__lane8_strm0_ready      ),      
               .std__pe57__lane8_strm0_cntl          ( std__pe57__lane8_strm0_cntl       ),      
               .std__pe57__lane8_strm0_data          ( std__pe57__lane8_strm0_data       ),      
               .std__pe57__lane8_strm0_data_valid    ( std__pe57__lane8_strm0_data_valid ),      
               .std__pe57__lane8_strm0_data_mask     ( std__pe57__lane8_strm0_data_mask  ),      

               .pe57__std__lane8_strm1_ready         ( pe57__std__lane8_strm1_ready      ),      
               .std__pe57__lane8_strm1_cntl          ( std__pe57__lane8_strm1_cntl       ),      
               .std__pe57__lane8_strm1_data          ( std__pe57__lane8_strm1_data       ),      
               .std__pe57__lane8_strm1_data_valid    ( std__pe57__lane8_strm1_data_valid ),      
               .std__pe57__lane8_strm1_data_mask     ( std__pe57__lane8_strm1_data_mask  ),      

               // PE 57, Lane 9                 
               .pe57__std__lane9_strm0_ready         ( pe57__std__lane9_strm0_ready      ),      
               .std__pe57__lane9_strm0_cntl          ( std__pe57__lane9_strm0_cntl       ),      
               .std__pe57__lane9_strm0_data          ( std__pe57__lane9_strm0_data       ),      
               .std__pe57__lane9_strm0_data_valid    ( std__pe57__lane9_strm0_data_valid ),      
               .std__pe57__lane9_strm0_data_mask     ( std__pe57__lane9_strm0_data_mask  ),      

               .pe57__std__lane9_strm1_ready         ( pe57__std__lane9_strm1_ready      ),      
               .std__pe57__lane9_strm1_cntl          ( std__pe57__lane9_strm1_cntl       ),      
               .std__pe57__lane9_strm1_data          ( std__pe57__lane9_strm1_data       ),      
               .std__pe57__lane9_strm1_data_valid    ( std__pe57__lane9_strm1_data_valid ),      
               .std__pe57__lane9_strm1_data_mask     ( std__pe57__lane9_strm1_data_mask  ),      

               // PE 57, Lane 10                 
               .pe57__std__lane10_strm0_ready         ( pe57__std__lane10_strm0_ready      ),      
               .std__pe57__lane10_strm0_cntl          ( std__pe57__lane10_strm0_cntl       ),      
               .std__pe57__lane10_strm0_data          ( std__pe57__lane10_strm0_data       ),      
               .std__pe57__lane10_strm0_data_valid    ( std__pe57__lane10_strm0_data_valid ),      
               .std__pe57__lane10_strm0_data_mask     ( std__pe57__lane10_strm0_data_mask  ),      

               .pe57__std__lane10_strm1_ready         ( pe57__std__lane10_strm1_ready      ),      
               .std__pe57__lane10_strm1_cntl          ( std__pe57__lane10_strm1_cntl       ),      
               .std__pe57__lane10_strm1_data          ( std__pe57__lane10_strm1_data       ),      
               .std__pe57__lane10_strm1_data_valid    ( std__pe57__lane10_strm1_data_valid ),      
               .std__pe57__lane10_strm1_data_mask     ( std__pe57__lane10_strm1_data_mask  ),      

               // PE 57, Lane 11                 
               .pe57__std__lane11_strm0_ready         ( pe57__std__lane11_strm0_ready      ),      
               .std__pe57__lane11_strm0_cntl          ( std__pe57__lane11_strm0_cntl       ),      
               .std__pe57__lane11_strm0_data          ( std__pe57__lane11_strm0_data       ),      
               .std__pe57__lane11_strm0_data_valid    ( std__pe57__lane11_strm0_data_valid ),      
               .std__pe57__lane11_strm0_data_mask     ( std__pe57__lane11_strm0_data_mask  ),      

               .pe57__std__lane11_strm1_ready         ( pe57__std__lane11_strm1_ready      ),      
               .std__pe57__lane11_strm1_cntl          ( std__pe57__lane11_strm1_cntl       ),      
               .std__pe57__lane11_strm1_data          ( std__pe57__lane11_strm1_data       ),      
               .std__pe57__lane11_strm1_data_valid    ( std__pe57__lane11_strm1_data_valid ),      
               .std__pe57__lane11_strm1_data_mask     ( std__pe57__lane11_strm1_data_mask  ),      

               // PE 57, Lane 12                 
               .pe57__std__lane12_strm0_ready         ( pe57__std__lane12_strm0_ready      ),      
               .std__pe57__lane12_strm0_cntl          ( std__pe57__lane12_strm0_cntl       ),      
               .std__pe57__lane12_strm0_data          ( std__pe57__lane12_strm0_data       ),      
               .std__pe57__lane12_strm0_data_valid    ( std__pe57__lane12_strm0_data_valid ),      
               .std__pe57__lane12_strm0_data_mask     ( std__pe57__lane12_strm0_data_mask  ),      

               .pe57__std__lane12_strm1_ready         ( pe57__std__lane12_strm1_ready      ),      
               .std__pe57__lane12_strm1_cntl          ( std__pe57__lane12_strm1_cntl       ),      
               .std__pe57__lane12_strm1_data          ( std__pe57__lane12_strm1_data       ),      
               .std__pe57__lane12_strm1_data_valid    ( std__pe57__lane12_strm1_data_valid ),      
               .std__pe57__lane12_strm1_data_mask     ( std__pe57__lane12_strm1_data_mask  ),      

               // PE 57, Lane 13                 
               .pe57__std__lane13_strm0_ready         ( pe57__std__lane13_strm0_ready      ),      
               .std__pe57__lane13_strm0_cntl          ( std__pe57__lane13_strm0_cntl       ),      
               .std__pe57__lane13_strm0_data          ( std__pe57__lane13_strm0_data       ),      
               .std__pe57__lane13_strm0_data_valid    ( std__pe57__lane13_strm0_data_valid ),      
               .std__pe57__lane13_strm0_data_mask     ( std__pe57__lane13_strm0_data_mask  ),      

               .pe57__std__lane13_strm1_ready         ( pe57__std__lane13_strm1_ready      ),      
               .std__pe57__lane13_strm1_cntl          ( std__pe57__lane13_strm1_cntl       ),      
               .std__pe57__lane13_strm1_data          ( std__pe57__lane13_strm1_data       ),      
               .std__pe57__lane13_strm1_data_valid    ( std__pe57__lane13_strm1_data_valid ),      
               .std__pe57__lane13_strm1_data_mask     ( std__pe57__lane13_strm1_data_mask  ),      

               // PE 57, Lane 14                 
               .pe57__std__lane14_strm0_ready         ( pe57__std__lane14_strm0_ready      ),      
               .std__pe57__lane14_strm0_cntl          ( std__pe57__lane14_strm0_cntl       ),      
               .std__pe57__lane14_strm0_data          ( std__pe57__lane14_strm0_data       ),      
               .std__pe57__lane14_strm0_data_valid    ( std__pe57__lane14_strm0_data_valid ),      
               .std__pe57__lane14_strm0_data_mask     ( std__pe57__lane14_strm0_data_mask  ),      

               .pe57__std__lane14_strm1_ready         ( pe57__std__lane14_strm1_ready      ),      
               .std__pe57__lane14_strm1_cntl          ( std__pe57__lane14_strm1_cntl       ),      
               .std__pe57__lane14_strm1_data          ( std__pe57__lane14_strm1_data       ),      
               .std__pe57__lane14_strm1_data_valid    ( std__pe57__lane14_strm1_data_valid ),      
               .std__pe57__lane14_strm1_data_mask     ( std__pe57__lane14_strm1_data_mask  ),      

               // PE 57, Lane 15                 
               .pe57__std__lane15_strm0_ready         ( pe57__std__lane15_strm0_ready      ),      
               .std__pe57__lane15_strm0_cntl          ( std__pe57__lane15_strm0_cntl       ),      
               .std__pe57__lane15_strm0_data          ( std__pe57__lane15_strm0_data       ),      
               .std__pe57__lane15_strm0_data_valid    ( std__pe57__lane15_strm0_data_valid ),      
               .std__pe57__lane15_strm0_data_mask     ( std__pe57__lane15_strm0_data_mask  ),      

               .pe57__std__lane15_strm1_ready         ( pe57__std__lane15_strm1_ready      ),      
               .std__pe57__lane15_strm1_cntl          ( std__pe57__lane15_strm1_cntl       ),      
               .std__pe57__lane15_strm1_data          ( std__pe57__lane15_strm1_data       ),      
               .std__pe57__lane15_strm1_data_valid    ( std__pe57__lane15_strm1_data_valid ),      
               .std__pe57__lane15_strm1_data_mask     ( std__pe57__lane15_strm1_data_mask  ),      

               // PE 57, Lane 16                 
               .pe57__std__lane16_strm0_ready         ( pe57__std__lane16_strm0_ready      ),      
               .std__pe57__lane16_strm0_cntl          ( std__pe57__lane16_strm0_cntl       ),      
               .std__pe57__lane16_strm0_data          ( std__pe57__lane16_strm0_data       ),      
               .std__pe57__lane16_strm0_data_valid    ( std__pe57__lane16_strm0_data_valid ),      
               .std__pe57__lane16_strm0_data_mask     ( std__pe57__lane16_strm0_data_mask  ),      

               .pe57__std__lane16_strm1_ready         ( pe57__std__lane16_strm1_ready      ),      
               .std__pe57__lane16_strm1_cntl          ( std__pe57__lane16_strm1_cntl       ),      
               .std__pe57__lane16_strm1_data          ( std__pe57__lane16_strm1_data       ),      
               .std__pe57__lane16_strm1_data_valid    ( std__pe57__lane16_strm1_data_valid ),      
               .std__pe57__lane16_strm1_data_mask     ( std__pe57__lane16_strm1_data_mask  ),      

               // PE 57, Lane 17                 
               .pe57__std__lane17_strm0_ready         ( pe57__std__lane17_strm0_ready      ),      
               .std__pe57__lane17_strm0_cntl          ( std__pe57__lane17_strm0_cntl       ),      
               .std__pe57__lane17_strm0_data          ( std__pe57__lane17_strm0_data       ),      
               .std__pe57__lane17_strm0_data_valid    ( std__pe57__lane17_strm0_data_valid ),      
               .std__pe57__lane17_strm0_data_mask     ( std__pe57__lane17_strm0_data_mask  ),      

               .pe57__std__lane17_strm1_ready         ( pe57__std__lane17_strm1_ready      ),      
               .std__pe57__lane17_strm1_cntl          ( std__pe57__lane17_strm1_cntl       ),      
               .std__pe57__lane17_strm1_data          ( std__pe57__lane17_strm1_data       ),      
               .std__pe57__lane17_strm1_data_valid    ( std__pe57__lane17_strm1_data_valid ),      
               .std__pe57__lane17_strm1_data_mask     ( std__pe57__lane17_strm1_data_mask  ),      

               // PE 57, Lane 18                 
               .pe57__std__lane18_strm0_ready         ( pe57__std__lane18_strm0_ready      ),      
               .std__pe57__lane18_strm0_cntl          ( std__pe57__lane18_strm0_cntl       ),      
               .std__pe57__lane18_strm0_data          ( std__pe57__lane18_strm0_data       ),      
               .std__pe57__lane18_strm0_data_valid    ( std__pe57__lane18_strm0_data_valid ),      
               .std__pe57__lane18_strm0_data_mask     ( std__pe57__lane18_strm0_data_mask  ),      

               .pe57__std__lane18_strm1_ready         ( pe57__std__lane18_strm1_ready      ),      
               .std__pe57__lane18_strm1_cntl          ( std__pe57__lane18_strm1_cntl       ),      
               .std__pe57__lane18_strm1_data          ( std__pe57__lane18_strm1_data       ),      
               .std__pe57__lane18_strm1_data_valid    ( std__pe57__lane18_strm1_data_valid ),      
               .std__pe57__lane18_strm1_data_mask     ( std__pe57__lane18_strm1_data_mask  ),      

               // PE 57, Lane 19                 
               .pe57__std__lane19_strm0_ready         ( pe57__std__lane19_strm0_ready      ),      
               .std__pe57__lane19_strm0_cntl          ( std__pe57__lane19_strm0_cntl       ),      
               .std__pe57__lane19_strm0_data          ( std__pe57__lane19_strm0_data       ),      
               .std__pe57__lane19_strm0_data_valid    ( std__pe57__lane19_strm0_data_valid ),      
               .std__pe57__lane19_strm0_data_mask     ( std__pe57__lane19_strm0_data_mask  ),      

               .pe57__std__lane19_strm1_ready         ( pe57__std__lane19_strm1_ready      ),      
               .std__pe57__lane19_strm1_cntl          ( std__pe57__lane19_strm1_cntl       ),      
               .std__pe57__lane19_strm1_data          ( std__pe57__lane19_strm1_data       ),      
               .std__pe57__lane19_strm1_data_valid    ( std__pe57__lane19_strm1_data_valid ),      
               .std__pe57__lane19_strm1_data_mask     ( std__pe57__lane19_strm1_data_mask  ),      

               // PE 57, Lane 20                 
               .pe57__std__lane20_strm0_ready         ( pe57__std__lane20_strm0_ready      ),      
               .std__pe57__lane20_strm0_cntl          ( std__pe57__lane20_strm0_cntl       ),      
               .std__pe57__lane20_strm0_data          ( std__pe57__lane20_strm0_data       ),      
               .std__pe57__lane20_strm0_data_valid    ( std__pe57__lane20_strm0_data_valid ),      
               .std__pe57__lane20_strm0_data_mask     ( std__pe57__lane20_strm0_data_mask  ),      

               .pe57__std__lane20_strm1_ready         ( pe57__std__lane20_strm1_ready      ),      
               .std__pe57__lane20_strm1_cntl          ( std__pe57__lane20_strm1_cntl       ),      
               .std__pe57__lane20_strm1_data          ( std__pe57__lane20_strm1_data       ),      
               .std__pe57__lane20_strm1_data_valid    ( std__pe57__lane20_strm1_data_valid ),      
               .std__pe57__lane20_strm1_data_mask     ( std__pe57__lane20_strm1_data_mask  ),      

               // PE 57, Lane 21                 
               .pe57__std__lane21_strm0_ready         ( pe57__std__lane21_strm0_ready      ),      
               .std__pe57__lane21_strm0_cntl          ( std__pe57__lane21_strm0_cntl       ),      
               .std__pe57__lane21_strm0_data          ( std__pe57__lane21_strm0_data       ),      
               .std__pe57__lane21_strm0_data_valid    ( std__pe57__lane21_strm0_data_valid ),      
               .std__pe57__lane21_strm0_data_mask     ( std__pe57__lane21_strm0_data_mask  ),      

               .pe57__std__lane21_strm1_ready         ( pe57__std__lane21_strm1_ready      ),      
               .std__pe57__lane21_strm1_cntl          ( std__pe57__lane21_strm1_cntl       ),      
               .std__pe57__lane21_strm1_data          ( std__pe57__lane21_strm1_data       ),      
               .std__pe57__lane21_strm1_data_valid    ( std__pe57__lane21_strm1_data_valid ),      
               .std__pe57__lane21_strm1_data_mask     ( std__pe57__lane21_strm1_data_mask  ),      

               // PE 57, Lane 22                 
               .pe57__std__lane22_strm0_ready         ( pe57__std__lane22_strm0_ready      ),      
               .std__pe57__lane22_strm0_cntl          ( std__pe57__lane22_strm0_cntl       ),      
               .std__pe57__lane22_strm0_data          ( std__pe57__lane22_strm0_data       ),      
               .std__pe57__lane22_strm0_data_valid    ( std__pe57__lane22_strm0_data_valid ),      
               .std__pe57__lane22_strm0_data_mask     ( std__pe57__lane22_strm0_data_mask  ),      

               .pe57__std__lane22_strm1_ready         ( pe57__std__lane22_strm1_ready      ),      
               .std__pe57__lane22_strm1_cntl          ( std__pe57__lane22_strm1_cntl       ),      
               .std__pe57__lane22_strm1_data          ( std__pe57__lane22_strm1_data       ),      
               .std__pe57__lane22_strm1_data_valid    ( std__pe57__lane22_strm1_data_valid ),      
               .std__pe57__lane22_strm1_data_mask     ( std__pe57__lane22_strm1_data_mask  ),      

               // PE 57, Lane 23                 
               .pe57__std__lane23_strm0_ready         ( pe57__std__lane23_strm0_ready      ),      
               .std__pe57__lane23_strm0_cntl          ( std__pe57__lane23_strm0_cntl       ),      
               .std__pe57__lane23_strm0_data          ( std__pe57__lane23_strm0_data       ),      
               .std__pe57__lane23_strm0_data_valid    ( std__pe57__lane23_strm0_data_valid ),      
               .std__pe57__lane23_strm0_data_mask     ( std__pe57__lane23_strm0_data_mask  ),      

               .pe57__std__lane23_strm1_ready         ( pe57__std__lane23_strm1_ready      ),      
               .std__pe57__lane23_strm1_cntl          ( std__pe57__lane23_strm1_cntl       ),      
               .std__pe57__lane23_strm1_data          ( std__pe57__lane23_strm1_data       ),      
               .std__pe57__lane23_strm1_data_valid    ( std__pe57__lane23_strm1_data_valid ),      
               .std__pe57__lane23_strm1_data_mask     ( std__pe57__lane23_strm1_data_mask  ),      

               // PE 57, Lane 24                 
               .pe57__std__lane24_strm0_ready         ( pe57__std__lane24_strm0_ready      ),      
               .std__pe57__lane24_strm0_cntl          ( std__pe57__lane24_strm0_cntl       ),      
               .std__pe57__lane24_strm0_data          ( std__pe57__lane24_strm0_data       ),      
               .std__pe57__lane24_strm0_data_valid    ( std__pe57__lane24_strm0_data_valid ),      
               .std__pe57__lane24_strm0_data_mask     ( std__pe57__lane24_strm0_data_mask  ),      

               .pe57__std__lane24_strm1_ready         ( pe57__std__lane24_strm1_ready      ),      
               .std__pe57__lane24_strm1_cntl          ( std__pe57__lane24_strm1_cntl       ),      
               .std__pe57__lane24_strm1_data          ( std__pe57__lane24_strm1_data       ),      
               .std__pe57__lane24_strm1_data_valid    ( std__pe57__lane24_strm1_data_valid ),      
               .std__pe57__lane24_strm1_data_mask     ( std__pe57__lane24_strm1_data_mask  ),      

               // PE 57, Lane 25                 
               .pe57__std__lane25_strm0_ready         ( pe57__std__lane25_strm0_ready      ),      
               .std__pe57__lane25_strm0_cntl          ( std__pe57__lane25_strm0_cntl       ),      
               .std__pe57__lane25_strm0_data          ( std__pe57__lane25_strm0_data       ),      
               .std__pe57__lane25_strm0_data_valid    ( std__pe57__lane25_strm0_data_valid ),      
               .std__pe57__lane25_strm0_data_mask     ( std__pe57__lane25_strm0_data_mask  ),      

               .pe57__std__lane25_strm1_ready         ( pe57__std__lane25_strm1_ready      ),      
               .std__pe57__lane25_strm1_cntl          ( std__pe57__lane25_strm1_cntl       ),      
               .std__pe57__lane25_strm1_data          ( std__pe57__lane25_strm1_data       ),      
               .std__pe57__lane25_strm1_data_valid    ( std__pe57__lane25_strm1_data_valid ),      
               .std__pe57__lane25_strm1_data_mask     ( std__pe57__lane25_strm1_data_mask  ),      

               // PE 57, Lane 26                 
               .pe57__std__lane26_strm0_ready         ( pe57__std__lane26_strm0_ready      ),      
               .std__pe57__lane26_strm0_cntl          ( std__pe57__lane26_strm0_cntl       ),      
               .std__pe57__lane26_strm0_data          ( std__pe57__lane26_strm0_data       ),      
               .std__pe57__lane26_strm0_data_valid    ( std__pe57__lane26_strm0_data_valid ),      
               .std__pe57__lane26_strm0_data_mask     ( std__pe57__lane26_strm0_data_mask  ),      

               .pe57__std__lane26_strm1_ready         ( pe57__std__lane26_strm1_ready      ),      
               .std__pe57__lane26_strm1_cntl          ( std__pe57__lane26_strm1_cntl       ),      
               .std__pe57__lane26_strm1_data          ( std__pe57__lane26_strm1_data       ),      
               .std__pe57__lane26_strm1_data_valid    ( std__pe57__lane26_strm1_data_valid ),      
               .std__pe57__lane26_strm1_data_mask     ( std__pe57__lane26_strm1_data_mask  ),      

               // PE 57, Lane 27                 
               .pe57__std__lane27_strm0_ready         ( pe57__std__lane27_strm0_ready      ),      
               .std__pe57__lane27_strm0_cntl          ( std__pe57__lane27_strm0_cntl       ),      
               .std__pe57__lane27_strm0_data          ( std__pe57__lane27_strm0_data       ),      
               .std__pe57__lane27_strm0_data_valid    ( std__pe57__lane27_strm0_data_valid ),      
               .std__pe57__lane27_strm0_data_mask     ( std__pe57__lane27_strm0_data_mask  ),      

               .pe57__std__lane27_strm1_ready         ( pe57__std__lane27_strm1_ready      ),      
               .std__pe57__lane27_strm1_cntl          ( std__pe57__lane27_strm1_cntl       ),      
               .std__pe57__lane27_strm1_data          ( std__pe57__lane27_strm1_data       ),      
               .std__pe57__lane27_strm1_data_valid    ( std__pe57__lane27_strm1_data_valid ),      
               .std__pe57__lane27_strm1_data_mask     ( std__pe57__lane27_strm1_data_mask  ),      

               // PE 57, Lane 28                 
               .pe57__std__lane28_strm0_ready         ( pe57__std__lane28_strm0_ready      ),      
               .std__pe57__lane28_strm0_cntl          ( std__pe57__lane28_strm0_cntl       ),      
               .std__pe57__lane28_strm0_data          ( std__pe57__lane28_strm0_data       ),      
               .std__pe57__lane28_strm0_data_valid    ( std__pe57__lane28_strm0_data_valid ),      
               .std__pe57__lane28_strm0_data_mask     ( std__pe57__lane28_strm0_data_mask  ),      

               .pe57__std__lane28_strm1_ready         ( pe57__std__lane28_strm1_ready      ),      
               .std__pe57__lane28_strm1_cntl          ( std__pe57__lane28_strm1_cntl       ),      
               .std__pe57__lane28_strm1_data          ( std__pe57__lane28_strm1_data       ),      
               .std__pe57__lane28_strm1_data_valid    ( std__pe57__lane28_strm1_data_valid ),      
               .std__pe57__lane28_strm1_data_mask     ( std__pe57__lane28_strm1_data_mask  ),      

               // PE 57, Lane 29                 
               .pe57__std__lane29_strm0_ready         ( pe57__std__lane29_strm0_ready      ),      
               .std__pe57__lane29_strm0_cntl          ( std__pe57__lane29_strm0_cntl       ),      
               .std__pe57__lane29_strm0_data          ( std__pe57__lane29_strm0_data       ),      
               .std__pe57__lane29_strm0_data_valid    ( std__pe57__lane29_strm0_data_valid ),      
               .std__pe57__lane29_strm0_data_mask     ( std__pe57__lane29_strm0_data_mask  ),      

               .pe57__std__lane29_strm1_ready         ( pe57__std__lane29_strm1_ready      ),      
               .std__pe57__lane29_strm1_cntl          ( std__pe57__lane29_strm1_cntl       ),      
               .std__pe57__lane29_strm1_data          ( std__pe57__lane29_strm1_data       ),      
               .std__pe57__lane29_strm1_data_valid    ( std__pe57__lane29_strm1_data_valid ),      
               .std__pe57__lane29_strm1_data_mask     ( std__pe57__lane29_strm1_data_mask  ),      

               // PE 57, Lane 30                 
               .pe57__std__lane30_strm0_ready         ( pe57__std__lane30_strm0_ready      ),      
               .std__pe57__lane30_strm0_cntl          ( std__pe57__lane30_strm0_cntl       ),      
               .std__pe57__lane30_strm0_data          ( std__pe57__lane30_strm0_data       ),      
               .std__pe57__lane30_strm0_data_valid    ( std__pe57__lane30_strm0_data_valid ),      
               .std__pe57__lane30_strm0_data_mask     ( std__pe57__lane30_strm0_data_mask  ),      

               .pe57__std__lane30_strm1_ready         ( pe57__std__lane30_strm1_ready      ),      
               .std__pe57__lane30_strm1_cntl          ( std__pe57__lane30_strm1_cntl       ),      
               .std__pe57__lane30_strm1_data          ( std__pe57__lane30_strm1_data       ),      
               .std__pe57__lane30_strm1_data_valid    ( std__pe57__lane30_strm1_data_valid ),      
               .std__pe57__lane30_strm1_data_mask     ( std__pe57__lane30_strm1_data_mask  ),      

               // PE 57, Lane 31                 
               .pe57__std__lane31_strm0_ready         ( pe57__std__lane31_strm0_ready      ),      
               .std__pe57__lane31_strm0_cntl          ( std__pe57__lane31_strm0_cntl       ),      
               .std__pe57__lane31_strm0_data          ( std__pe57__lane31_strm0_data       ),      
               .std__pe57__lane31_strm0_data_valid    ( std__pe57__lane31_strm0_data_valid ),      
               .std__pe57__lane31_strm0_data_mask     ( std__pe57__lane31_strm0_data_mask  ),      

               .pe57__std__lane31_strm1_ready         ( pe57__std__lane31_strm1_ready      ),      
               .std__pe57__lane31_strm1_cntl          ( std__pe57__lane31_strm1_cntl       ),      
               .std__pe57__lane31_strm1_data          ( std__pe57__lane31_strm1_data       ),      
               .std__pe57__lane31_strm1_data_valid    ( std__pe57__lane31_strm1_data_valid ),      
               .std__pe57__lane31_strm1_data_mask     ( std__pe57__lane31_strm1_data_mask  ),      

               // PE 58, Lane 0                 
               .pe58__std__lane0_strm0_ready         ( pe58__std__lane0_strm0_ready      ),      
               .std__pe58__lane0_strm0_cntl          ( std__pe58__lane0_strm0_cntl       ),      
               .std__pe58__lane0_strm0_data          ( std__pe58__lane0_strm0_data       ),      
               .std__pe58__lane0_strm0_data_valid    ( std__pe58__lane0_strm0_data_valid ),      
               .std__pe58__lane0_strm0_data_mask     ( std__pe58__lane0_strm0_data_mask  ),      

               .pe58__std__lane0_strm1_ready         ( pe58__std__lane0_strm1_ready      ),      
               .std__pe58__lane0_strm1_cntl          ( std__pe58__lane0_strm1_cntl       ),      
               .std__pe58__lane0_strm1_data          ( std__pe58__lane0_strm1_data       ),      
               .std__pe58__lane0_strm1_data_valid    ( std__pe58__lane0_strm1_data_valid ),      
               .std__pe58__lane0_strm1_data_mask     ( std__pe58__lane0_strm1_data_mask  ),      

               // PE 58, Lane 1                 
               .pe58__std__lane1_strm0_ready         ( pe58__std__lane1_strm0_ready      ),      
               .std__pe58__lane1_strm0_cntl          ( std__pe58__lane1_strm0_cntl       ),      
               .std__pe58__lane1_strm0_data          ( std__pe58__lane1_strm0_data       ),      
               .std__pe58__lane1_strm0_data_valid    ( std__pe58__lane1_strm0_data_valid ),      
               .std__pe58__lane1_strm0_data_mask     ( std__pe58__lane1_strm0_data_mask  ),      

               .pe58__std__lane1_strm1_ready         ( pe58__std__lane1_strm1_ready      ),      
               .std__pe58__lane1_strm1_cntl          ( std__pe58__lane1_strm1_cntl       ),      
               .std__pe58__lane1_strm1_data          ( std__pe58__lane1_strm1_data       ),      
               .std__pe58__lane1_strm1_data_valid    ( std__pe58__lane1_strm1_data_valid ),      
               .std__pe58__lane1_strm1_data_mask     ( std__pe58__lane1_strm1_data_mask  ),      

               // PE 58, Lane 2                 
               .pe58__std__lane2_strm0_ready         ( pe58__std__lane2_strm0_ready      ),      
               .std__pe58__lane2_strm0_cntl          ( std__pe58__lane2_strm0_cntl       ),      
               .std__pe58__lane2_strm0_data          ( std__pe58__lane2_strm0_data       ),      
               .std__pe58__lane2_strm0_data_valid    ( std__pe58__lane2_strm0_data_valid ),      
               .std__pe58__lane2_strm0_data_mask     ( std__pe58__lane2_strm0_data_mask  ),      

               .pe58__std__lane2_strm1_ready         ( pe58__std__lane2_strm1_ready      ),      
               .std__pe58__lane2_strm1_cntl          ( std__pe58__lane2_strm1_cntl       ),      
               .std__pe58__lane2_strm1_data          ( std__pe58__lane2_strm1_data       ),      
               .std__pe58__lane2_strm1_data_valid    ( std__pe58__lane2_strm1_data_valid ),      
               .std__pe58__lane2_strm1_data_mask     ( std__pe58__lane2_strm1_data_mask  ),      

               // PE 58, Lane 3                 
               .pe58__std__lane3_strm0_ready         ( pe58__std__lane3_strm0_ready      ),      
               .std__pe58__lane3_strm0_cntl          ( std__pe58__lane3_strm0_cntl       ),      
               .std__pe58__lane3_strm0_data          ( std__pe58__lane3_strm0_data       ),      
               .std__pe58__lane3_strm0_data_valid    ( std__pe58__lane3_strm0_data_valid ),      
               .std__pe58__lane3_strm0_data_mask     ( std__pe58__lane3_strm0_data_mask  ),      

               .pe58__std__lane3_strm1_ready         ( pe58__std__lane3_strm1_ready      ),      
               .std__pe58__lane3_strm1_cntl          ( std__pe58__lane3_strm1_cntl       ),      
               .std__pe58__lane3_strm1_data          ( std__pe58__lane3_strm1_data       ),      
               .std__pe58__lane3_strm1_data_valid    ( std__pe58__lane3_strm1_data_valid ),      
               .std__pe58__lane3_strm1_data_mask     ( std__pe58__lane3_strm1_data_mask  ),      

               // PE 58, Lane 4                 
               .pe58__std__lane4_strm0_ready         ( pe58__std__lane4_strm0_ready      ),      
               .std__pe58__lane4_strm0_cntl          ( std__pe58__lane4_strm0_cntl       ),      
               .std__pe58__lane4_strm0_data          ( std__pe58__lane4_strm0_data       ),      
               .std__pe58__lane4_strm0_data_valid    ( std__pe58__lane4_strm0_data_valid ),      
               .std__pe58__lane4_strm0_data_mask     ( std__pe58__lane4_strm0_data_mask  ),      

               .pe58__std__lane4_strm1_ready         ( pe58__std__lane4_strm1_ready      ),      
               .std__pe58__lane4_strm1_cntl          ( std__pe58__lane4_strm1_cntl       ),      
               .std__pe58__lane4_strm1_data          ( std__pe58__lane4_strm1_data       ),      
               .std__pe58__lane4_strm1_data_valid    ( std__pe58__lane4_strm1_data_valid ),      
               .std__pe58__lane4_strm1_data_mask     ( std__pe58__lane4_strm1_data_mask  ),      

               // PE 58, Lane 5                 
               .pe58__std__lane5_strm0_ready         ( pe58__std__lane5_strm0_ready      ),      
               .std__pe58__lane5_strm0_cntl          ( std__pe58__lane5_strm0_cntl       ),      
               .std__pe58__lane5_strm0_data          ( std__pe58__lane5_strm0_data       ),      
               .std__pe58__lane5_strm0_data_valid    ( std__pe58__lane5_strm0_data_valid ),      
               .std__pe58__lane5_strm0_data_mask     ( std__pe58__lane5_strm0_data_mask  ),      

               .pe58__std__lane5_strm1_ready         ( pe58__std__lane5_strm1_ready      ),      
               .std__pe58__lane5_strm1_cntl          ( std__pe58__lane5_strm1_cntl       ),      
               .std__pe58__lane5_strm1_data          ( std__pe58__lane5_strm1_data       ),      
               .std__pe58__lane5_strm1_data_valid    ( std__pe58__lane5_strm1_data_valid ),      
               .std__pe58__lane5_strm1_data_mask     ( std__pe58__lane5_strm1_data_mask  ),      

               // PE 58, Lane 6                 
               .pe58__std__lane6_strm0_ready         ( pe58__std__lane6_strm0_ready      ),      
               .std__pe58__lane6_strm0_cntl          ( std__pe58__lane6_strm0_cntl       ),      
               .std__pe58__lane6_strm0_data          ( std__pe58__lane6_strm0_data       ),      
               .std__pe58__lane6_strm0_data_valid    ( std__pe58__lane6_strm0_data_valid ),      
               .std__pe58__lane6_strm0_data_mask     ( std__pe58__lane6_strm0_data_mask  ),      

               .pe58__std__lane6_strm1_ready         ( pe58__std__lane6_strm1_ready      ),      
               .std__pe58__lane6_strm1_cntl          ( std__pe58__lane6_strm1_cntl       ),      
               .std__pe58__lane6_strm1_data          ( std__pe58__lane6_strm1_data       ),      
               .std__pe58__lane6_strm1_data_valid    ( std__pe58__lane6_strm1_data_valid ),      
               .std__pe58__lane6_strm1_data_mask     ( std__pe58__lane6_strm1_data_mask  ),      

               // PE 58, Lane 7                 
               .pe58__std__lane7_strm0_ready         ( pe58__std__lane7_strm0_ready      ),      
               .std__pe58__lane7_strm0_cntl          ( std__pe58__lane7_strm0_cntl       ),      
               .std__pe58__lane7_strm0_data          ( std__pe58__lane7_strm0_data       ),      
               .std__pe58__lane7_strm0_data_valid    ( std__pe58__lane7_strm0_data_valid ),      
               .std__pe58__lane7_strm0_data_mask     ( std__pe58__lane7_strm0_data_mask  ),      

               .pe58__std__lane7_strm1_ready         ( pe58__std__lane7_strm1_ready      ),      
               .std__pe58__lane7_strm1_cntl          ( std__pe58__lane7_strm1_cntl       ),      
               .std__pe58__lane7_strm1_data          ( std__pe58__lane7_strm1_data       ),      
               .std__pe58__lane7_strm1_data_valid    ( std__pe58__lane7_strm1_data_valid ),      
               .std__pe58__lane7_strm1_data_mask     ( std__pe58__lane7_strm1_data_mask  ),      

               // PE 58, Lane 8                 
               .pe58__std__lane8_strm0_ready         ( pe58__std__lane8_strm0_ready      ),      
               .std__pe58__lane8_strm0_cntl          ( std__pe58__lane8_strm0_cntl       ),      
               .std__pe58__lane8_strm0_data          ( std__pe58__lane8_strm0_data       ),      
               .std__pe58__lane8_strm0_data_valid    ( std__pe58__lane8_strm0_data_valid ),      
               .std__pe58__lane8_strm0_data_mask     ( std__pe58__lane8_strm0_data_mask  ),      

               .pe58__std__lane8_strm1_ready         ( pe58__std__lane8_strm1_ready      ),      
               .std__pe58__lane8_strm1_cntl          ( std__pe58__lane8_strm1_cntl       ),      
               .std__pe58__lane8_strm1_data          ( std__pe58__lane8_strm1_data       ),      
               .std__pe58__lane8_strm1_data_valid    ( std__pe58__lane8_strm1_data_valid ),      
               .std__pe58__lane8_strm1_data_mask     ( std__pe58__lane8_strm1_data_mask  ),      

               // PE 58, Lane 9                 
               .pe58__std__lane9_strm0_ready         ( pe58__std__lane9_strm0_ready      ),      
               .std__pe58__lane9_strm0_cntl          ( std__pe58__lane9_strm0_cntl       ),      
               .std__pe58__lane9_strm0_data          ( std__pe58__lane9_strm0_data       ),      
               .std__pe58__lane9_strm0_data_valid    ( std__pe58__lane9_strm0_data_valid ),      
               .std__pe58__lane9_strm0_data_mask     ( std__pe58__lane9_strm0_data_mask  ),      

               .pe58__std__lane9_strm1_ready         ( pe58__std__lane9_strm1_ready      ),      
               .std__pe58__lane9_strm1_cntl          ( std__pe58__lane9_strm1_cntl       ),      
               .std__pe58__lane9_strm1_data          ( std__pe58__lane9_strm1_data       ),      
               .std__pe58__lane9_strm1_data_valid    ( std__pe58__lane9_strm1_data_valid ),      
               .std__pe58__lane9_strm1_data_mask     ( std__pe58__lane9_strm1_data_mask  ),      

               // PE 58, Lane 10                 
               .pe58__std__lane10_strm0_ready         ( pe58__std__lane10_strm0_ready      ),      
               .std__pe58__lane10_strm0_cntl          ( std__pe58__lane10_strm0_cntl       ),      
               .std__pe58__lane10_strm0_data          ( std__pe58__lane10_strm0_data       ),      
               .std__pe58__lane10_strm0_data_valid    ( std__pe58__lane10_strm0_data_valid ),      
               .std__pe58__lane10_strm0_data_mask     ( std__pe58__lane10_strm0_data_mask  ),      

               .pe58__std__lane10_strm1_ready         ( pe58__std__lane10_strm1_ready      ),      
               .std__pe58__lane10_strm1_cntl          ( std__pe58__lane10_strm1_cntl       ),      
               .std__pe58__lane10_strm1_data          ( std__pe58__lane10_strm1_data       ),      
               .std__pe58__lane10_strm1_data_valid    ( std__pe58__lane10_strm1_data_valid ),      
               .std__pe58__lane10_strm1_data_mask     ( std__pe58__lane10_strm1_data_mask  ),      

               // PE 58, Lane 11                 
               .pe58__std__lane11_strm0_ready         ( pe58__std__lane11_strm0_ready      ),      
               .std__pe58__lane11_strm0_cntl          ( std__pe58__lane11_strm0_cntl       ),      
               .std__pe58__lane11_strm0_data          ( std__pe58__lane11_strm0_data       ),      
               .std__pe58__lane11_strm0_data_valid    ( std__pe58__lane11_strm0_data_valid ),      
               .std__pe58__lane11_strm0_data_mask     ( std__pe58__lane11_strm0_data_mask  ),      

               .pe58__std__lane11_strm1_ready         ( pe58__std__lane11_strm1_ready      ),      
               .std__pe58__lane11_strm1_cntl          ( std__pe58__lane11_strm1_cntl       ),      
               .std__pe58__lane11_strm1_data          ( std__pe58__lane11_strm1_data       ),      
               .std__pe58__lane11_strm1_data_valid    ( std__pe58__lane11_strm1_data_valid ),      
               .std__pe58__lane11_strm1_data_mask     ( std__pe58__lane11_strm1_data_mask  ),      

               // PE 58, Lane 12                 
               .pe58__std__lane12_strm0_ready         ( pe58__std__lane12_strm0_ready      ),      
               .std__pe58__lane12_strm0_cntl          ( std__pe58__lane12_strm0_cntl       ),      
               .std__pe58__lane12_strm0_data          ( std__pe58__lane12_strm0_data       ),      
               .std__pe58__lane12_strm0_data_valid    ( std__pe58__lane12_strm0_data_valid ),      
               .std__pe58__lane12_strm0_data_mask     ( std__pe58__lane12_strm0_data_mask  ),      

               .pe58__std__lane12_strm1_ready         ( pe58__std__lane12_strm1_ready      ),      
               .std__pe58__lane12_strm1_cntl          ( std__pe58__lane12_strm1_cntl       ),      
               .std__pe58__lane12_strm1_data          ( std__pe58__lane12_strm1_data       ),      
               .std__pe58__lane12_strm1_data_valid    ( std__pe58__lane12_strm1_data_valid ),      
               .std__pe58__lane12_strm1_data_mask     ( std__pe58__lane12_strm1_data_mask  ),      

               // PE 58, Lane 13                 
               .pe58__std__lane13_strm0_ready         ( pe58__std__lane13_strm0_ready      ),      
               .std__pe58__lane13_strm0_cntl          ( std__pe58__lane13_strm0_cntl       ),      
               .std__pe58__lane13_strm0_data          ( std__pe58__lane13_strm0_data       ),      
               .std__pe58__lane13_strm0_data_valid    ( std__pe58__lane13_strm0_data_valid ),      
               .std__pe58__lane13_strm0_data_mask     ( std__pe58__lane13_strm0_data_mask  ),      

               .pe58__std__lane13_strm1_ready         ( pe58__std__lane13_strm1_ready      ),      
               .std__pe58__lane13_strm1_cntl          ( std__pe58__lane13_strm1_cntl       ),      
               .std__pe58__lane13_strm1_data          ( std__pe58__lane13_strm1_data       ),      
               .std__pe58__lane13_strm1_data_valid    ( std__pe58__lane13_strm1_data_valid ),      
               .std__pe58__lane13_strm1_data_mask     ( std__pe58__lane13_strm1_data_mask  ),      

               // PE 58, Lane 14                 
               .pe58__std__lane14_strm0_ready         ( pe58__std__lane14_strm0_ready      ),      
               .std__pe58__lane14_strm0_cntl          ( std__pe58__lane14_strm0_cntl       ),      
               .std__pe58__lane14_strm0_data          ( std__pe58__lane14_strm0_data       ),      
               .std__pe58__lane14_strm0_data_valid    ( std__pe58__lane14_strm0_data_valid ),      
               .std__pe58__lane14_strm0_data_mask     ( std__pe58__lane14_strm0_data_mask  ),      

               .pe58__std__lane14_strm1_ready         ( pe58__std__lane14_strm1_ready      ),      
               .std__pe58__lane14_strm1_cntl          ( std__pe58__lane14_strm1_cntl       ),      
               .std__pe58__lane14_strm1_data          ( std__pe58__lane14_strm1_data       ),      
               .std__pe58__lane14_strm1_data_valid    ( std__pe58__lane14_strm1_data_valid ),      
               .std__pe58__lane14_strm1_data_mask     ( std__pe58__lane14_strm1_data_mask  ),      

               // PE 58, Lane 15                 
               .pe58__std__lane15_strm0_ready         ( pe58__std__lane15_strm0_ready      ),      
               .std__pe58__lane15_strm0_cntl          ( std__pe58__lane15_strm0_cntl       ),      
               .std__pe58__lane15_strm0_data          ( std__pe58__lane15_strm0_data       ),      
               .std__pe58__lane15_strm0_data_valid    ( std__pe58__lane15_strm0_data_valid ),      
               .std__pe58__lane15_strm0_data_mask     ( std__pe58__lane15_strm0_data_mask  ),      

               .pe58__std__lane15_strm1_ready         ( pe58__std__lane15_strm1_ready      ),      
               .std__pe58__lane15_strm1_cntl          ( std__pe58__lane15_strm1_cntl       ),      
               .std__pe58__lane15_strm1_data          ( std__pe58__lane15_strm1_data       ),      
               .std__pe58__lane15_strm1_data_valid    ( std__pe58__lane15_strm1_data_valid ),      
               .std__pe58__lane15_strm1_data_mask     ( std__pe58__lane15_strm1_data_mask  ),      

               // PE 58, Lane 16                 
               .pe58__std__lane16_strm0_ready         ( pe58__std__lane16_strm0_ready      ),      
               .std__pe58__lane16_strm0_cntl          ( std__pe58__lane16_strm0_cntl       ),      
               .std__pe58__lane16_strm0_data          ( std__pe58__lane16_strm0_data       ),      
               .std__pe58__lane16_strm0_data_valid    ( std__pe58__lane16_strm0_data_valid ),      
               .std__pe58__lane16_strm0_data_mask     ( std__pe58__lane16_strm0_data_mask  ),      

               .pe58__std__lane16_strm1_ready         ( pe58__std__lane16_strm1_ready      ),      
               .std__pe58__lane16_strm1_cntl          ( std__pe58__lane16_strm1_cntl       ),      
               .std__pe58__lane16_strm1_data          ( std__pe58__lane16_strm1_data       ),      
               .std__pe58__lane16_strm1_data_valid    ( std__pe58__lane16_strm1_data_valid ),      
               .std__pe58__lane16_strm1_data_mask     ( std__pe58__lane16_strm1_data_mask  ),      

               // PE 58, Lane 17                 
               .pe58__std__lane17_strm0_ready         ( pe58__std__lane17_strm0_ready      ),      
               .std__pe58__lane17_strm0_cntl          ( std__pe58__lane17_strm0_cntl       ),      
               .std__pe58__lane17_strm0_data          ( std__pe58__lane17_strm0_data       ),      
               .std__pe58__lane17_strm0_data_valid    ( std__pe58__lane17_strm0_data_valid ),      
               .std__pe58__lane17_strm0_data_mask     ( std__pe58__lane17_strm0_data_mask  ),      

               .pe58__std__lane17_strm1_ready         ( pe58__std__lane17_strm1_ready      ),      
               .std__pe58__lane17_strm1_cntl          ( std__pe58__lane17_strm1_cntl       ),      
               .std__pe58__lane17_strm1_data          ( std__pe58__lane17_strm1_data       ),      
               .std__pe58__lane17_strm1_data_valid    ( std__pe58__lane17_strm1_data_valid ),      
               .std__pe58__lane17_strm1_data_mask     ( std__pe58__lane17_strm1_data_mask  ),      

               // PE 58, Lane 18                 
               .pe58__std__lane18_strm0_ready         ( pe58__std__lane18_strm0_ready      ),      
               .std__pe58__lane18_strm0_cntl          ( std__pe58__lane18_strm0_cntl       ),      
               .std__pe58__lane18_strm0_data          ( std__pe58__lane18_strm0_data       ),      
               .std__pe58__lane18_strm0_data_valid    ( std__pe58__lane18_strm0_data_valid ),      
               .std__pe58__lane18_strm0_data_mask     ( std__pe58__lane18_strm0_data_mask  ),      

               .pe58__std__lane18_strm1_ready         ( pe58__std__lane18_strm1_ready      ),      
               .std__pe58__lane18_strm1_cntl          ( std__pe58__lane18_strm1_cntl       ),      
               .std__pe58__lane18_strm1_data          ( std__pe58__lane18_strm1_data       ),      
               .std__pe58__lane18_strm1_data_valid    ( std__pe58__lane18_strm1_data_valid ),      
               .std__pe58__lane18_strm1_data_mask     ( std__pe58__lane18_strm1_data_mask  ),      

               // PE 58, Lane 19                 
               .pe58__std__lane19_strm0_ready         ( pe58__std__lane19_strm0_ready      ),      
               .std__pe58__lane19_strm0_cntl          ( std__pe58__lane19_strm0_cntl       ),      
               .std__pe58__lane19_strm0_data          ( std__pe58__lane19_strm0_data       ),      
               .std__pe58__lane19_strm0_data_valid    ( std__pe58__lane19_strm0_data_valid ),      
               .std__pe58__lane19_strm0_data_mask     ( std__pe58__lane19_strm0_data_mask  ),      

               .pe58__std__lane19_strm1_ready         ( pe58__std__lane19_strm1_ready      ),      
               .std__pe58__lane19_strm1_cntl          ( std__pe58__lane19_strm1_cntl       ),      
               .std__pe58__lane19_strm1_data          ( std__pe58__lane19_strm1_data       ),      
               .std__pe58__lane19_strm1_data_valid    ( std__pe58__lane19_strm1_data_valid ),      
               .std__pe58__lane19_strm1_data_mask     ( std__pe58__lane19_strm1_data_mask  ),      

               // PE 58, Lane 20                 
               .pe58__std__lane20_strm0_ready         ( pe58__std__lane20_strm0_ready      ),      
               .std__pe58__lane20_strm0_cntl          ( std__pe58__lane20_strm0_cntl       ),      
               .std__pe58__lane20_strm0_data          ( std__pe58__lane20_strm0_data       ),      
               .std__pe58__lane20_strm0_data_valid    ( std__pe58__lane20_strm0_data_valid ),      
               .std__pe58__lane20_strm0_data_mask     ( std__pe58__lane20_strm0_data_mask  ),      

               .pe58__std__lane20_strm1_ready         ( pe58__std__lane20_strm1_ready      ),      
               .std__pe58__lane20_strm1_cntl          ( std__pe58__lane20_strm1_cntl       ),      
               .std__pe58__lane20_strm1_data          ( std__pe58__lane20_strm1_data       ),      
               .std__pe58__lane20_strm1_data_valid    ( std__pe58__lane20_strm1_data_valid ),      
               .std__pe58__lane20_strm1_data_mask     ( std__pe58__lane20_strm1_data_mask  ),      

               // PE 58, Lane 21                 
               .pe58__std__lane21_strm0_ready         ( pe58__std__lane21_strm0_ready      ),      
               .std__pe58__lane21_strm0_cntl          ( std__pe58__lane21_strm0_cntl       ),      
               .std__pe58__lane21_strm0_data          ( std__pe58__lane21_strm0_data       ),      
               .std__pe58__lane21_strm0_data_valid    ( std__pe58__lane21_strm0_data_valid ),      
               .std__pe58__lane21_strm0_data_mask     ( std__pe58__lane21_strm0_data_mask  ),      

               .pe58__std__lane21_strm1_ready         ( pe58__std__lane21_strm1_ready      ),      
               .std__pe58__lane21_strm1_cntl          ( std__pe58__lane21_strm1_cntl       ),      
               .std__pe58__lane21_strm1_data          ( std__pe58__lane21_strm1_data       ),      
               .std__pe58__lane21_strm1_data_valid    ( std__pe58__lane21_strm1_data_valid ),      
               .std__pe58__lane21_strm1_data_mask     ( std__pe58__lane21_strm1_data_mask  ),      

               // PE 58, Lane 22                 
               .pe58__std__lane22_strm0_ready         ( pe58__std__lane22_strm0_ready      ),      
               .std__pe58__lane22_strm0_cntl          ( std__pe58__lane22_strm0_cntl       ),      
               .std__pe58__lane22_strm0_data          ( std__pe58__lane22_strm0_data       ),      
               .std__pe58__lane22_strm0_data_valid    ( std__pe58__lane22_strm0_data_valid ),      
               .std__pe58__lane22_strm0_data_mask     ( std__pe58__lane22_strm0_data_mask  ),      

               .pe58__std__lane22_strm1_ready         ( pe58__std__lane22_strm1_ready      ),      
               .std__pe58__lane22_strm1_cntl          ( std__pe58__lane22_strm1_cntl       ),      
               .std__pe58__lane22_strm1_data          ( std__pe58__lane22_strm1_data       ),      
               .std__pe58__lane22_strm1_data_valid    ( std__pe58__lane22_strm1_data_valid ),      
               .std__pe58__lane22_strm1_data_mask     ( std__pe58__lane22_strm1_data_mask  ),      

               // PE 58, Lane 23                 
               .pe58__std__lane23_strm0_ready         ( pe58__std__lane23_strm0_ready      ),      
               .std__pe58__lane23_strm0_cntl          ( std__pe58__lane23_strm0_cntl       ),      
               .std__pe58__lane23_strm0_data          ( std__pe58__lane23_strm0_data       ),      
               .std__pe58__lane23_strm0_data_valid    ( std__pe58__lane23_strm0_data_valid ),      
               .std__pe58__lane23_strm0_data_mask     ( std__pe58__lane23_strm0_data_mask  ),      

               .pe58__std__lane23_strm1_ready         ( pe58__std__lane23_strm1_ready      ),      
               .std__pe58__lane23_strm1_cntl          ( std__pe58__lane23_strm1_cntl       ),      
               .std__pe58__lane23_strm1_data          ( std__pe58__lane23_strm1_data       ),      
               .std__pe58__lane23_strm1_data_valid    ( std__pe58__lane23_strm1_data_valid ),      
               .std__pe58__lane23_strm1_data_mask     ( std__pe58__lane23_strm1_data_mask  ),      

               // PE 58, Lane 24                 
               .pe58__std__lane24_strm0_ready         ( pe58__std__lane24_strm0_ready      ),      
               .std__pe58__lane24_strm0_cntl          ( std__pe58__lane24_strm0_cntl       ),      
               .std__pe58__lane24_strm0_data          ( std__pe58__lane24_strm0_data       ),      
               .std__pe58__lane24_strm0_data_valid    ( std__pe58__lane24_strm0_data_valid ),      
               .std__pe58__lane24_strm0_data_mask     ( std__pe58__lane24_strm0_data_mask  ),      

               .pe58__std__lane24_strm1_ready         ( pe58__std__lane24_strm1_ready      ),      
               .std__pe58__lane24_strm1_cntl          ( std__pe58__lane24_strm1_cntl       ),      
               .std__pe58__lane24_strm1_data          ( std__pe58__lane24_strm1_data       ),      
               .std__pe58__lane24_strm1_data_valid    ( std__pe58__lane24_strm1_data_valid ),      
               .std__pe58__lane24_strm1_data_mask     ( std__pe58__lane24_strm1_data_mask  ),      

               // PE 58, Lane 25                 
               .pe58__std__lane25_strm0_ready         ( pe58__std__lane25_strm0_ready      ),      
               .std__pe58__lane25_strm0_cntl          ( std__pe58__lane25_strm0_cntl       ),      
               .std__pe58__lane25_strm0_data          ( std__pe58__lane25_strm0_data       ),      
               .std__pe58__lane25_strm0_data_valid    ( std__pe58__lane25_strm0_data_valid ),      
               .std__pe58__lane25_strm0_data_mask     ( std__pe58__lane25_strm0_data_mask  ),      

               .pe58__std__lane25_strm1_ready         ( pe58__std__lane25_strm1_ready      ),      
               .std__pe58__lane25_strm1_cntl          ( std__pe58__lane25_strm1_cntl       ),      
               .std__pe58__lane25_strm1_data          ( std__pe58__lane25_strm1_data       ),      
               .std__pe58__lane25_strm1_data_valid    ( std__pe58__lane25_strm1_data_valid ),      
               .std__pe58__lane25_strm1_data_mask     ( std__pe58__lane25_strm1_data_mask  ),      

               // PE 58, Lane 26                 
               .pe58__std__lane26_strm0_ready         ( pe58__std__lane26_strm0_ready      ),      
               .std__pe58__lane26_strm0_cntl          ( std__pe58__lane26_strm0_cntl       ),      
               .std__pe58__lane26_strm0_data          ( std__pe58__lane26_strm0_data       ),      
               .std__pe58__lane26_strm0_data_valid    ( std__pe58__lane26_strm0_data_valid ),      
               .std__pe58__lane26_strm0_data_mask     ( std__pe58__lane26_strm0_data_mask  ),      

               .pe58__std__lane26_strm1_ready         ( pe58__std__lane26_strm1_ready      ),      
               .std__pe58__lane26_strm1_cntl          ( std__pe58__lane26_strm1_cntl       ),      
               .std__pe58__lane26_strm1_data          ( std__pe58__lane26_strm1_data       ),      
               .std__pe58__lane26_strm1_data_valid    ( std__pe58__lane26_strm1_data_valid ),      
               .std__pe58__lane26_strm1_data_mask     ( std__pe58__lane26_strm1_data_mask  ),      

               // PE 58, Lane 27                 
               .pe58__std__lane27_strm0_ready         ( pe58__std__lane27_strm0_ready      ),      
               .std__pe58__lane27_strm0_cntl          ( std__pe58__lane27_strm0_cntl       ),      
               .std__pe58__lane27_strm0_data          ( std__pe58__lane27_strm0_data       ),      
               .std__pe58__lane27_strm0_data_valid    ( std__pe58__lane27_strm0_data_valid ),      
               .std__pe58__lane27_strm0_data_mask     ( std__pe58__lane27_strm0_data_mask  ),      

               .pe58__std__lane27_strm1_ready         ( pe58__std__lane27_strm1_ready      ),      
               .std__pe58__lane27_strm1_cntl          ( std__pe58__lane27_strm1_cntl       ),      
               .std__pe58__lane27_strm1_data          ( std__pe58__lane27_strm1_data       ),      
               .std__pe58__lane27_strm1_data_valid    ( std__pe58__lane27_strm1_data_valid ),      
               .std__pe58__lane27_strm1_data_mask     ( std__pe58__lane27_strm1_data_mask  ),      

               // PE 58, Lane 28                 
               .pe58__std__lane28_strm0_ready         ( pe58__std__lane28_strm0_ready      ),      
               .std__pe58__lane28_strm0_cntl          ( std__pe58__lane28_strm0_cntl       ),      
               .std__pe58__lane28_strm0_data          ( std__pe58__lane28_strm0_data       ),      
               .std__pe58__lane28_strm0_data_valid    ( std__pe58__lane28_strm0_data_valid ),      
               .std__pe58__lane28_strm0_data_mask     ( std__pe58__lane28_strm0_data_mask  ),      

               .pe58__std__lane28_strm1_ready         ( pe58__std__lane28_strm1_ready      ),      
               .std__pe58__lane28_strm1_cntl          ( std__pe58__lane28_strm1_cntl       ),      
               .std__pe58__lane28_strm1_data          ( std__pe58__lane28_strm1_data       ),      
               .std__pe58__lane28_strm1_data_valid    ( std__pe58__lane28_strm1_data_valid ),      
               .std__pe58__lane28_strm1_data_mask     ( std__pe58__lane28_strm1_data_mask  ),      

               // PE 58, Lane 29                 
               .pe58__std__lane29_strm0_ready         ( pe58__std__lane29_strm0_ready      ),      
               .std__pe58__lane29_strm0_cntl          ( std__pe58__lane29_strm0_cntl       ),      
               .std__pe58__lane29_strm0_data          ( std__pe58__lane29_strm0_data       ),      
               .std__pe58__lane29_strm0_data_valid    ( std__pe58__lane29_strm0_data_valid ),      
               .std__pe58__lane29_strm0_data_mask     ( std__pe58__lane29_strm0_data_mask  ),      

               .pe58__std__lane29_strm1_ready         ( pe58__std__lane29_strm1_ready      ),      
               .std__pe58__lane29_strm1_cntl          ( std__pe58__lane29_strm1_cntl       ),      
               .std__pe58__lane29_strm1_data          ( std__pe58__lane29_strm1_data       ),      
               .std__pe58__lane29_strm1_data_valid    ( std__pe58__lane29_strm1_data_valid ),      
               .std__pe58__lane29_strm1_data_mask     ( std__pe58__lane29_strm1_data_mask  ),      

               // PE 58, Lane 30                 
               .pe58__std__lane30_strm0_ready         ( pe58__std__lane30_strm0_ready      ),      
               .std__pe58__lane30_strm0_cntl          ( std__pe58__lane30_strm0_cntl       ),      
               .std__pe58__lane30_strm0_data          ( std__pe58__lane30_strm0_data       ),      
               .std__pe58__lane30_strm0_data_valid    ( std__pe58__lane30_strm0_data_valid ),      
               .std__pe58__lane30_strm0_data_mask     ( std__pe58__lane30_strm0_data_mask  ),      

               .pe58__std__lane30_strm1_ready         ( pe58__std__lane30_strm1_ready      ),      
               .std__pe58__lane30_strm1_cntl          ( std__pe58__lane30_strm1_cntl       ),      
               .std__pe58__lane30_strm1_data          ( std__pe58__lane30_strm1_data       ),      
               .std__pe58__lane30_strm1_data_valid    ( std__pe58__lane30_strm1_data_valid ),      
               .std__pe58__lane30_strm1_data_mask     ( std__pe58__lane30_strm1_data_mask  ),      

               // PE 58, Lane 31                 
               .pe58__std__lane31_strm0_ready         ( pe58__std__lane31_strm0_ready      ),      
               .std__pe58__lane31_strm0_cntl          ( std__pe58__lane31_strm0_cntl       ),      
               .std__pe58__lane31_strm0_data          ( std__pe58__lane31_strm0_data       ),      
               .std__pe58__lane31_strm0_data_valid    ( std__pe58__lane31_strm0_data_valid ),      
               .std__pe58__lane31_strm0_data_mask     ( std__pe58__lane31_strm0_data_mask  ),      

               .pe58__std__lane31_strm1_ready         ( pe58__std__lane31_strm1_ready      ),      
               .std__pe58__lane31_strm1_cntl          ( std__pe58__lane31_strm1_cntl       ),      
               .std__pe58__lane31_strm1_data          ( std__pe58__lane31_strm1_data       ),      
               .std__pe58__lane31_strm1_data_valid    ( std__pe58__lane31_strm1_data_valid ),      
               .std__pe58__lane31_strm1_data_mask     ( std__pe58__lane31_strm1_data_mask  ),      

               // PE 59, Lane 0                 
               .pe59__std__lane0_strm0_ready         ( pe59__std__lane0_strm0_ready      ),      
               .std__pe59__lane0_strm0_cntl          ( std__pe59__lane0_strm0_cntl       ),      
               .std__pe59__lane0_strm0_data          ( std__pe59__lane0_strm0_data       ),      
               .std__pe59__lane0_strm0_data_valid    ( std__pe59__lane0_strm0_data_valid ),      
               .std__pe59__lane0_strm0_data_mask     ( std__pe59__lane0_strm0_data_mask  ),      

               .pe59__std__lane0_strm1_ready         ( pe59__std__lane0_strm1_ready      ),      
               .std__pe59__lane0_strm1_cntl          ( std__pe59__lane0_strm1_cntl       ),      
               .std__pe59__lane0_strm1_data          ( std__pe59__lane0_strm1_data       ),      
               .std__pe59__lane0_strm1_data_valid    ( std__pe59__lane0_strm1_data_valid ),      
               .std__pe59__lane0_strm1_data_mask     ( std__pe59__lane0_strm1_data_mask  ),      

               // PE 59, Lane 1                 
               .pe59__std__lane1_strm0_ready         ( pe59__std__lane1_strm0_ready      ),      
               .std__pe59__lane1_strm0_cntl          ( std__pe59__lane1_strm0_cntl       ),      
               .std__pe59__lane1_strm0_data          ( std__pe59__lane1_strm0_data       ),      
               .std__pe59__lane1_strm0_data_valid    ( std__pe59__lane1_strm0_data_valid ),      
               .std__pe59__lane1_strm0_data_mask     ( std__pe59__lane1_strm0_data_mask  ),      

               .pe59__std__lane1_strm1_ready         ( pe59__std__lane1_strm1_ready      ),      
               .std__pe59__lane1_strm1_cntl          ( std__pe59__lane1_strm1_cntl       ),      
               .std__pe59__lane1_strm1_data          ( std__pe59__lane1_strm1_data       ),      
               .std__pe59__lane1_strm1_data_valid    ( std__pe59__lane1_strm1_data_valid ),      
               .std__pe59__lane1_strm1_data_mask     ( std__pe59__lane1_strm1_data_mask  ),      

               // PE 59, Lane 2                 
               .pe59__std__lane2_strm0_ready         ( pe59__std__lane2_strm0_ready      ),      
               .std__pe59__lane2_strm0_cntl          ( std__pe59__lane2_strm0_cntl       ),      
               .std__pe59__lane2_strm0_data          ( std__pe59__lane2_strm0_data       ),      
               .std__pe59__lane2_strm0_data_valid    ( std__pe59__lane2_strm0_data_valid ),      
               .std__pe59__lane2_strm0_data_mask     ( std__pe59__lane2_strm0_data_mask  ),      

               .pe59__std__lane2_strm1_ready         ( pe59__std__lane2_strm1_ready      ),      
               .std__pe59__lane2_strm1_cntl          ( std__pe59__lane2_strm1_cntl       ),      
               .std__pe59__lane2_strm1_data          ( std__pe59__lane2_strm1_data       ),      
               .std__pe59__lane2_strm1_data_valid    ( std__pe59__lane2_strm1_data_valid ),      
               .std__pe59__lane2_strm1_data_mask     ( std__pe59__lane2_strm1_data_mask  ),      

               // PE 59, Lane 3                 
               .pe59__std__lane3_strm0_ready         ( pe59__std__lane3_strm0_ready      ),      
               .std__pe59__lane3_strm0_cntl          ( std__pe59__lane3_strm0_cntl       ),      
               .std__pe59__lane3_strm0_data          ( std__pe59__lane3_strm0_data       ),      
               .std__pe59__lane3_strm0_data_valid    ( std__pe59__lane3_strm0_data_valid ),      
               .std__pe59__lane3_strm0_data_mask     ( std__pe59__lane3_strm0_data_mask  ),      

               .pe59__std__lane3_strm1_ready         ( pe59__std__lane3_strm1_ready      ),      
               .std__pe59__lane3_strm1_cntl          ( std__pe59__lane3_strm1_cntl       ),      
               .std__pe59__lane3_strm1_data          ( std__pe59__lane3_strm1_data       ),      
               .std__pe59__lane3_strm1_data_valid    ( std__pe59__lane3_strm1_data_valid ),      
               .std__pe59__lane3_strm1_data_mask     ( std__pe59__lane3_strm1_data_mask  ),      

               // PE 59, Lane 4                 
               .pe59__std__lane4_strm0_ready         ( pe59__std__lane4_strm0_ready      ),      
               .std__pe59__lane4_strm0_cntl          ( std__pe59__lane4_strm0_cntl       ),      
               .std__pe59__lane4_strm0_data          ( std__pe59__lane4_strm0_data       ),      
               .std__pe59__lane4_strm0_data_valid    ( std__pe59__lane4_strm0_data_valid ),      
               .std__pe59__lane4_strm0_data_mask     ( std__pe59__lane4_strm0_data_mask  ),      

               .pe59__std__lane4_strm1_ready         ( pe59__std__lane4_strm1_ready      ),      
               .std__pe59__lane4_strm1_cntl          ( std__pe59__lane4_strm1_cntl       ),      
               .std__pe59__lane4_strm1_data          ( std__pe59__lane4_strm1_data       ),      
               .std__pe59__lane4_strm1_data_valid    ( std__pe59__lane4_strm1_data_valid ),      
               .std__pe59__lane4_strm1_data_mask     ( std__pe59__lane4_strm1_data_mask  ),      

               // PE 59, Lane 5                 
               .pe59__std__lane5_strm0_ready         ( pe59__std__lane5_strm0_ready      ),      
               .std__pe59__lane5_strm0_cntl          ( std__pe59__lane5_strm0_cntl       ),      
               .std__pe59__lane5_strm0_data          ( std__pe59__lane5_strm0_data       ),      
               .std__pe59__lane5_strm0_data_valid    ( std__pe59__lane5_strm0_data_valid ),      
               .std__pe59__lane5_strm0_data_mask     ( std__pe59__lane5_strm0_data_mask  ),      

               .pe59__std__lane5_strm1_ready         ( pe59__std__lane5_strm1_ready      ),      
               .std__pe59__lane5_strm1_cntl          ( std__pe59__lane5_strm1_cntl       ),      
               .std__pe59__lane5_strm1_data          ( std__pe59__lane5_strm1_data       ),      
               .std__pe59__lane5_strm1_data_valid    ( std__pe59__lane5_strm1_data_valid ),      
               .std__pe59__lane5_strm1_data_mask     ( std__pe59__lane5_strm1_data_mask  ),      

               // PE 59, Lane 6                 
               .pe59__std__lane6_strm0_ready         ( pe59__std__lane6_strm0_ready      ),      
               .std__pe59__lane6_strm0_cntl          ( std__pe59__lane6_strm0_cntl       ),      
               .std__pe59__lane6_strm0_data          ( std__pe59__lane6_strm0_data       ),      
               .std__pe59__lane6_strm0_data_valid    ( std__pe59__lane6_strm0_data_valid ),      
               .std__pe59__lane6_strm0_data_mask     ( std__pe59__lane6_strm0_data_mask  ),      

               .pe59__std__lane6_strm1_ready         ( pe59__std__lane6_strm1_ready      ),      
               .std__pe59__lane6_strm1_cntl          ( std__pe59__lane6_strm1_cntl       ),      
               .std__pe59__lane6_strm1_data          ( std__pe59__lane6_strm1_data       ),      
               .std__pe59__lane6_strm1_data_valid    ( std__pe59__lane6_strm1_data_valid ),      
               .std__pe59__lane6_strm1_data_mask     ( std__pe59__lane6_strm1_data_mask  ),      

               // PE 59, Lane 7                 
               .pe59__std__lane7_strm0_ready         ( pe59__std__lane7_strm0_ready      ),      
               .std__pe59__lane7_strm0_cntl          ( std__pe59__lane7_strm0_cntl       ),      
               .std__pe59__lane7_strm0_data          ( std__pe59__lane7_strm0_data       ),      
               .std__pe59__lane7_strm0_data_valid    ( std__pe59__lane7_strm0_data_valid ),      
               .std__pe59__lane7_strm0_data_mask     ( std__pe59__lane7_strm0_data_mask  ),      

               .pe59__std__lane7_strm1_ready         ( pe59__std__lane7_strm1_ready      ),      
               .std__pe59__lane7_strm1_cntl          ( std__pe59__lane7_strm1_cntl       ),      
               .std__pe59__lane7_strm1_data          ( std__pe59__lane7_strm1_data       ),      
               .std__pe59__lane7_strm1_data_valid    ( std__pe59__lane7_strm1_data_valid ),      
               .std__pe59__lane7_strm1_data_mask     ( std__pe59__lane7_strm1_data_mask  ),      

               // PE 59, Lane 8                 
               .pe59__std__lane8_strm0_ready         ( pe59__std__lane8_strm0_ready      ),      
               .std__pe59__lane8_strm0_cntl          ( std__pe59__lane8_strm0_cntl       ),      
               .std__pe59__lane8_strm0_data          ( std__pe59__lane8_strm0_data       ),      
               .std__pe59__lane8_strm0_data_valid    ( std__pe59__lane8_strm0_data_valid ),      
               .std__pe59__lane8_strm0_data_mask     ( std__pe59__lane8_strm0_data_mask  ),      

               .pe59__std__lane8_strm1_ready         ( pe59__std__lane8_strm1_ready      ),      
               .std__pe59__lane8_strm1_cntl          ( std__pe59__lane8_strm1_cntl       ),      
               .std__pe59__lane8_strm1_data          ( std__pe59__lane8_strm1_data       ),      
               .std__pe59__lane8_strm1_data_valid    ( std__pe59__lane8_strm1_data_valid ),      
               .std__pe59__lane8_strm1_data_mask     ( std__pe59__lane8_strm1_data_mask  ),      

               // PE 59, Lane 9                 
               .pe59__std__lane9_strm0_ready         ( pe59__std__lane9_strm0_ready      ),      
               .std__pe59__lane9_strm0_cntl          ( std__pe59__lane9_strm0_cntl       ),      
               .std__pe59__lane9_strm0_data          ( std__pe59__lane9_strm0_data       ),      
               .std__pe59__lane9_strm0_data_valid    ( std__pe59__lane9_strm0_data_valid ),      
               .std__pe59__lane9_strm0_data_mask     ( std__pe59__lane9_strm0_data_mask  ),      

               .pe59__std__lane9_strm1_ready         ( pe59__std__lane9_strm1_ready      ),      
               .std__pe59__lane9_strm1_cntl          ( std__pe59__lane9_strm1_cntl       ),      
               .std__pe59__lane9_strm1_data          ( std__pe59__lane9_strm1_data       ),      
               .std__pe59__lane9_strm1_data_valid    ( std__pe59__lane9_strm1_data_valid ),      
               .std__pe59__lane9_strm1_data_mask     ( std__pe59__lane9_strm1_data_mask  ),      

               // PE 59, Lane 10                 
               .pe59__std__lane10_strm0_ready         ( pe59__std__lane10_strm0_ready      ),      
               .std__pe59__lane10_strm0_cntl          ( std__pe59__lane10_strm0_cntl       ),      
               .std__pe59__lane10_strm0_data          ( std__pe59__lane10_strm0_data       ),      
               .std__pe59__lane10_strm0_data_valid    ( std__pe59__lane10_strm0_data_valid ),      
               .std__pe59__lane10_strm0_data_mask     ( std__pe59__lane10_strm0_data_mask  ),      

               .pe59__std__lane10_strm1_ready         ( pe59__std__lane10_strm1_ready      ),      
               .std__pe59__lane10_strm1_cntl          ( std__pe59__lane10_strm1_cntl       ),      
               .std__pe59__lane10_strm1_data          ( std__pe59__lane10_strm1_data       ),      
               .std__pe59__lane10_strm1_data_valid    ( std__pe59__lane10_strm1_data_valid ),      
               .std__pe59__lane10_strm1_data_mask     ( std__pe59__lane10_strm1_data_mask  ),      

               // PE 59, Lane 11                 
               .pe59__std__lane11_strm0_ready         ( pe59__std__lane11_strm0_ready      ),      
               .std__pe59__lane11_strm0_cntl          ( std__pe59__lane11_strm0_cntl       ),      
               .std__pe59__lane11_strm0_data          ( std__pe59__lane11_strm0_data       ),      
               .std__pe59__lane11_strm0_data_valid    ( std__pe59__lane11_strm0_data_valid ),      
               .std__pe59__lane11_strm0_data_mask     ( std__pe59__lane11_strm0_data_mask  ),      

               .pe59__std__lane11_strm1_ready         ( pe59__std__lane11_strm1_ready      ),      
               .std__pe59__lane11_strm1_cntl          ( std__pe59__lane11_strm1_cntl       ),      
               .std__pe59__lane11_strm1_data          ( std__pe59__lane11_strm1_data       ),      
               .std__pe59__lane11_strm1_data_valid    ( std__pe59__lane11_strm1_data_valid ),      
               .std__pe59__lane11_strm1_data_mask     ( std__pe59__lane11_strm1_data_mask  ),      

               // PE 59, Lane 12                 
               .pe59__std__lane12_strm0_ready         ( pe59__std__lane12_strm0_ready      ),      
               .std__pe59__lane12_strm0_cntl          ( std__pe59__lane12_strm0_cntl       ),      
               .std__pe59__lane12_strm0_data          ( std__pe59__lane12_strm0_data       ),      
               .std__pe59__lane12_strm0_data_valid    ( std__pe59__lane12_strm0_data_valid ),      
               .std__pe59__lane12_strm0_data_mask     ( std__pe59__lane12_strm0_data_mask  ),      

               .pe59__std__lane12_strm1_ready         ( pe59__std__lane12_strm1_ready      ),      
               .std__pe59__lane12_strm1_cntl          ( std__pe59__lane12_strm1_cntl       ),      
               .std__pe59__lane12_strm1_data          ( std__pe59__lane12_strm1_data       ),      
               .std__pe59__lane12_strm1_data_valid    ( std__pe59__lane12_strm1_data_valid ),      
               .std__pe59__lane12_strm1_data_mask     ( std__pe59__lane12_strm1_data_mask  ),      

               // PE 59, Lane 13                 
               .pe59__std__lane13_strm0_ready         ( pe59__std__lane13_strm0_ready      ),      
               .std__pe59__lane13_strm0_cntl          ( std__pe59__lane13_strm0_cntl       ),      
               .std__pe59__lane13_strm0_data          ( std__pe59__lane13_strm0_data       ),      
               .std__pe59__lane13_strm0_data_valid    ( std__pe59__lane13_strm0_data_valid ),      
               .std__pe59__lane13_strm0_data_mask     ( std__pe59__lane13_strm0_data_mask  ),      

               .pe59__std__lane13_strm1_ready         ( pe59__std__lane13_strm1_ready      ),      
               .std__pe59__lane13_strm1_cntl          ( std__pe59__lane13_strm1_cntl       ),      
               .std__pe59__lane13_strm1_data          ( std__pe59__lane13_strm1_data       ),      
               .std__pe59__lane13_strm1_data_valid    ( std__pe59__lane13_strm1_data_valid ),      
               .std__pe59__lane13_strm1_data_mask     ( std__pe59__lane13_strm1_data_mask  ),      

               // PE 59, Lane 14                 
               .pe59__std__lane14_strm0_ready         ( pe59__std__lane14_strm0_ready      ),      
               .std__pe59__lane14_strm0_cntl          ( std__pe59__lane14_strm0_cntl       ),      
               .std__pe59__lane14_strm0_data          ( std__pe59__lane14_strm0_data       ),      
               .std__pe59__lane14_strm0_data_valid    ( std__pe59__lane14_strm0_data_valid ),      
               .std__pe59__lane14_strm0_data_mask     ( std__pe59__lane14_strm0_data_mask  ),      

               .pe59__std__lane14_strm1_ready         ( pe59__std__lane14_strm1_ready      ),      
               .std__pe59__lane14_strm1_cntl          ( std__pe59__lane14_strm1_cntl       ),      
               .std__pe59__lane14_strm1_data          ( std__pe59__lane14_strm1_data       ),      
               .std__pe59__lane14_strm1_data_valid    ( std__pe59__lane14_strm1_data_valid ),      
               .std__pe59__lane14_strm1_data_mask     ( std__pe59__lane14_strm1_data_mask  ),      

               // PE 59, Lane 15                 
               .pe59__std__lane15_strm0_ready         ( pe59__std__lane15_strm0_ready      ),      
               .std__pe59__lane15_strm0_cntl          ( std__pe59__lane15_strm0_cntl       ),      
               .std__pe59__lane15_strm0_data          ( std__pe59__lane15_strm0_data       ),      
               .std__pe59__lane15_strm0_data_valid    ( std__pe59__lane15_strm0_data_valid ),      
               .std__pe59__lane15_strm0_data_mask     ( std__pe59__lane15_strm0_data_mask  ),      

               .pe59__std__lane15_strm1_ready         ( pe59__std__lane15_strm1_ready      ),      
               .std__pe59__lane15_strm1_cntl          ( std__pe59__lane15_strm1_cntl       ),      
               .std__pe59__lane15_strm1_data          ( std__pe59__lane15_strm1_data       ),      
               .std__pe59__lane15_strm1_data_valid    ( std__pe59__lane15_strm1_data_valid ),      
               .std__pe59__lane15_strm1_data_mask     ( std__pe59__lane15_strm1_data_mask  ),      

               // PE 59, Lane 16                 
               .pe59__std__lane16_strm0_ready         ( pe59__std__lane16_strm0_ready      ),      
               .std__pe59__lane16_strm0_cntl          ( std__pe59__lane16_strm0_cntl       ),      
               .std__pe59__lane16_strm0_data          ( std__pe59__lane16_strm0_data       ),      
               .std__pe59__lane16_strm0_data_valid    ( std__pe59__lane16_strm0_data_valid ),      
               .std__pe59__lane16_strm0_data_mask     ( std__pe59__lane16_strm0_data_mask  ),      

               .pe59__std__lane16_strm1_ready         ( pe59__std__lane16_strm1_ready      ),      
               .std__pe59__lane16_strm1_cntl          ( std__pe59__lane16_strm1_cntl       ),      
               .std__pe59__lane16_strm1_data          ( std__pe59__lane16_strm1_data       ),      
               .std__pe59__lane16_strm1_data_valid    ( std__pe59__lane16_strm1_data_valid ),      
               .std__pe59__lane16_strm1_data_mask     ( std__pe59__lane16_strm1_data_mask  ),      

               // PE 59, Lane 17                 
               .pe59__std__lane17_strm0_ready         ( pe59__std__lane17_strm0_ready      ),      
               .std__pe59__lane17_strm0_cntl          ( std__pe59__lane17_strm0_cntl       ),      
               .std__pe59__lane17_strm0_data          ( std__pe59__lane17_strm0_data       ),      
               .std__pe59__lane17_strm0_data_valid    ( std__pe59__lane17_strm0_data_valid ),      
               .std__pe59__lane17_strm0_data_mask     ( std__pe59__lane17_strm0_data_mask  ),      

               .pe59__std__lane17_strm1_ready         ( pe59__std__lane17_strm1_ready      ),      
               .std__pe59__lane17_strm1_cntl          ( std__pe59__lane17_strm1_cntl       ),      
               .std__pe59__lane17_strm1_data          ( std__pe59__lane17_strm1_data       ),      
               .std__pe59__lane17_strm1_data_valid    ( std__pe59__lane17_strm1_data_valid ),      
               .std__pe59__lane17_strm1_data_mask     ( std__pe59__lane17_strm1_data_mask  ),      

               // PE 59, Lane 18                 
               .pe59__std__lane18_strm0_ready         ( pe59__std__lane18_strm0_ready      ),      
               .std__pe59__lane18_strm0_cntl          ( std__pe59__lane18_strm0_cntl       ),      
               .std__pe59__lane18_strm0_data          ( std__pe59__lane18_strm0_data       ),      
               .std__pe59__lane18_strm0_data_valid    ( std__pe59__lane18_strm0_data_valid ),      
               .std__pe59__lane18_strm0_data_mask     ( std__pe59__lane18_strm0_data_mask  ),      

               .pe59__std__lane18_strm1_ready         ( pe59__std__lane18_strm1_ready      ),      
               .std__pe59__lane18_strm1_cntl          ( std__pe59__lane18_strm1_cntl       ),      
               .std__pe59__lane18_strm1_data          ( std__pe59__lane18_strm1_data       ),      
               .std__pe59__lane18_strm1_data_valid    ( std__pe59__lane18_strm1_data_valid ),      
               .std__pe59__lane18_strm1_data_mask     ( std__pe59__lane18_strm1_data_mask  ),      

               // PE 59, Lane 19                 
               .pe59__std__lane19_strm0_ready         ( pe59__std__lane19_strm0_ready      ),      
               .std__pe59__lane19_strm0_cntl          ( std__pe59__lane19_strm0_cntl       ),      
               .std__pe59__lane19_strm0_data          ( std__pe59__lane19_strm0_data       ),      
               .std__pe59__lane19_strm0_data_valid    ( std__pe59__lane19_strm0_data_valid ),      
               .std__pe59__lane19_strm0_data_mask     ( std__pe59__lane19_strm0_data_mask  ),      

               .pe59__std__lane19_strm1_ready         ( pe59__std__lane19_strm1_ready      ),      
               .std__pe59__lane19_strm1_cntl          ( std__pe59__lane19_strm1_cntl       ),      
               .std__pe59__lane19_strm1_data          ( std__pe59__lane19_strm1_data       ),      
               .std__pe59__lane19_strm1_data_valid    ( std__pe59__lane19_strm1_data_valid ),      
               .std__pe59__lane19_strm1_data_mask     ( std__pe59__lane19_strm1_data_mask  ),      

               // PE 59, Lane 20                 
               .pe59__std__lane20_strm0_ready         ( pe59__std__lane20_strm0_ready      ),      
               .std__pe59__lane20_strm0_cntl          ( std__pe59__lane20_strm0_cntl       ),      
               .std__pe59__lane20_strm0_data          ( std__pe59__lane20_strm0_data       ),      
               .std__pe59__lane20_strm0_data_valid    ( std__pe59__lane20_strm0_data_valid ),      
               .std__pe59__lane20_strm0_data_mask     ( std__pe59__lane20_strm0_data_mask  ),      

               .pe59__std__lane20_strm1_ready         ( pe59__std__lane20_strm1_ready      ),      
               .std__pe59__lane20_strm1_cntl          ( std__pe59__lane20_strm1_cntl       ),      
               .std__pe59__lane20_strm1_data          ( std__pe59__lane20_strm1_data       ),      
               .std__pe59__lane20_strm1_data_valid    ( std__pe59__lane20_strm1_data_valid ),      
               .std__pe59__lane20_strm1_data_mask     ( std__pe59__lane20_strm1_data_mask  ),      

               // PE 59, Lane 21                 
               .pe59__std__lane21_strm0_ready         ( pe59__std__lane21_strm0_ready      ),      
               .std__pe59__lane21_strm0_cntl          ( std__pe59__lane21_strm0_cntl       ),      
               .std__pe59__lane21_strm0_data          ( std__pe59__lane21_strm0_data       ),      
               .std__pe59__lane21_strm0_data_valid    ( std__pe59__lane21_strm0_data_valid ),      
               .std__pe59__lane21_strm0_data_mask     ( std__pe59__lane21_strm0_data_mask  ),      

               .pe59__std__lane21_strm1_ready         ( pe59__std__lane21_strm1_ready      ),      
               .std__pe59__lane21_strm1_cntl          ( std__pe59__lane21_strm1_cntl       ),      
               .std__pe59__lane21_strm1_data          ( std__pe59__lane21_strm1_data       ),      
               .std__pe59__lane21_strm1_data_valid    ( std__pe59__lane21_strm1_data_valid ),      
               .std__pe59__lane21_strm1_data_mask     ( std__pe59__lane21_strm1_data_mask  ),      

               // PE 59, Lane 22                 
               .pe59__std__lane22_strm0_ready         ( pe59__std__lane22_strm0_ready      ),      
               .std__pe59__lane22_strm0_cntl          ( std__pe59__lane22_strm0_cntl       ),      
               .std__pe59__lane22_strm0_data          ( std__pe59__lane22_strm0_data       ),      
               .std__pe59__lane22_strm0_data_valid    ( std__pe59__lane22_strm0_data_valid ),      
               .std__pe59__lane22_strm0_data_mask     ( std__pe59__lane22_strm0_data_mask  ),      

               .pe59__std__lane22_strm1_ready         ( pe59__std__lane22_strm1_ready      ),      
               .std__pe59__lane22_strm1_cntl          ( std__pe59__lane22_strm1_cntl       ),      
               .std__pe59__lane22_strm1_data          ( std__pe59__lane22_strm1_data       ),      
               .std__pe59__lane22_strm1_data_valid    ( std__pe59__lane22_strm1_data_valid ),      
               .std__pe59__lane22_strm1_data_mask     ( std__pe59__lane22_strm1_data_mask  ),      

               // PE 59, Lane 23                 
               .pe59__std__lane23_strm0_ready         ( pe59__std__lane23_strm0_ready      ),      
               .std__pe59__lane23_strm0_cntl          ( std__pe59__lane23_strm0_cntl       ),      
               .std__pe59__lane23_strm0_data          ( std__pe59__lane23_strm0_data       ),      
               .std__pe59__lane23_strm0_data_valid    ( std__pe59__lane23_strm0_data_valid ),      
               .std__pe59__lane23_strm0_data_mask     ( std__pe59__lane23_strm0_data_mask  ),      

               .pe59__std__lane23_strm1_ready         ( pe59__std__lane23_strm1_ready      ),      
               .std__pe59__lane23_strm1_cntl          ( std__pe59__lane23_strm1_cntl       ),      
               .std__pe59__lane23_strm1_data          ( std__pe59__lane23_strm1_data       ),      
               .std__pe59__lane23_strm1_data_valid    ( std__pe59__lane23_strm1_data_valid ),      
               .std__pe59__lane23_strm1_data_mask     ( std__pe59__lane23_strm1_data_mask  ),      

               // PE 59, Lane 24                 
               .pe59__std__lane24_strm0_ready         ( pe59__std__lane24_strm0_ready      ),      
               .std__pe59__lane24_strm0_cntl          ( std__pe59__lane24_strm0_cntl       ),      
               .std__pe59__lane24_strm0_data          ( std__pe59__lane24_strm0_data       ),      
               .std__pe59__lane24_strm0_data_valid    ( std__pe59__lane24_strm0_data_valid ),      
               .std__pe59__lane24_strm0_data_mask     ( std__pe59__lane24_strm0_data_mask  ),      

               .pe59__std__lane24_strm1_ready         ( pe59__std__lane24_strm1_ready      ),      
               .std__pe59__lane24_strm1_cntl          ( std__pe59__lane24_strm1_cntl       ),      
               .std__pe59__lane24_strm1_data          ( std__pe59__lane24_strm1_data       ),      
               .std__pe59__lane24_strm1_data_valid    ( std__pe59__lane24_strm1_data_valid ),      
               .std__pe59__lane24_strm1_data_mask     ( std__pe59__lane24_strm1_data_mask  ),      

               // PE 59, Lane 25                 
               .pe59__std__lane25_strm0_ready         ( pe59__std__lane25_strm0_ready      ),      
               .std__pe59__lane25_strm0_cntl          ( std__pe59__lane25_strm0_cntl       ),      
               .std__pe59__lane25_strm0_data          ( std__pe59__lane25_strm0_data       ),      
               .std__pe59__lane25_strm0_data_valid    ( std__pe59__lane25_strm0_data_valid ),      
               .std__pe59__lane25_strm0_data_mask     ( std__pe59__lane25_strm0_data_mask  ),      

               .pe59__std__lane25_strm1_ready         ( pe59__std__lane25_strm1_ready      ),      
               .std__pe59__lane25_strm1_cntl          ( std__pe59__lane25_strm1_cntl       ),      
               .std__pe59__lane25_strm1_data          ( std__pe59__lane25_strm1_data       ),      
               .std__pe59__lane25_strm1_data_valid    ( std__pe59__lane25_strm1_data_valid ),      
               .std__pe59__lane25_strm1_data_mask     ( std__pe59__lane25_strm1_data_mask  ),      

               // PE 59, Lane 26                 
               .pe59__std__lane26_strm0_ready         ( pe59__std__lane26_strm0_ready      ),      
               .std__pe59__lane26_strm0_cntl          ( std__pe59__lane26_strm0_cntl       ),      
               .std__pe59__lane26_strm0_data          ( std__pe59__lane26_strm0_data       ),      
               .std__pe59__lane26_strm0_data_valid    ( std__pe59__lane26_strm0_data_valid ),      
               .std__pe59__lane26_strm0_data_mask     ( std__pe59__lane26_strm0_data_mask  ),      

               .pe59__std__lane26_strm1_ready         ( pe59__std__lane26_strm1_ready      ),      
               .std__pe59__lane26_strm1_cntl          ( std__pe59__lane26_strm1_cntl       ),      
               .std__pe59__lane26_strm1_data          ( std__pe59__lane26_strm1_data       ),      
               .std__pe59__lane26_strm1_data_valid    ( std__pe59__lane26_strm1_data_valid ),      
               .std__pe59__lane26_strm1_data_mask     ( std__pe59__lane26_strm1_data_mask  ),      

               // PE 59, Lane 27                 
               .pe59__std__lane27_strm0_ready         ( pe59__std__lane27_strm0_ready      ),      
               .std__pe59__lane27_strm0_cntl          ( std__pe59__lane27_strm0_cntl       ),      
               .std__pe59__lane27_strm0_data          ( std__pe59__lane27_strm0_data       ),      
               .std__pe59__lane27_strm0_data_valid    ( std__pe59__lane27_strm0_data_valid ),      
               .std__pe59__lane27_strm0_data_mask     ( std__pe59__lane27_strm0_data_mask  ),      

               .pe59__std__lane27_strm1_ready         ( pe59__std__lane27_strm1_ready      ),      
               .std__pe59__lane27_strm1_cntl          ( std__pe59__lane27_strm1_cntl       ),      
               .std__pe59__lane27_strm1_data          ( std__pe59__lane27_strm1_data       ),      
               .std__pe59__lane27_strm1_data_valid    ( std__pe59__lane27_strm1_data_valid ),      
               .std__pe59__lane27_strm1_data_mask     ( std__pe59__lane27_strm1_data_mask  ),      

               // PE 59, Lane 28                 
               .pe59__std__lane28_strm0_ready         ( pe59__std__lane28_strm0_ready      ),      
               .std__pe59__lane28_strm0_cntl          ( std__pe59__lane28_strm0_cntl       ),      
               .std__pe59__lane28_strm0_data          ( std__pe59__lane28_strm0_data       ),      
               .std__pe59__lane28_strm0_data_valid    ( std__pe59__lane28_strm0_data_valid ),      
               .std__pe59__lane28_strm0_data_mask     ( std__pe59__lane28_strm0_data_mask  ),      

               .pe59__std__lane28_strm1_ready         ( pe59__std__lane28_strm1_ready      ),      
               .std__pe59__lane28_strm1_cntl          ( std__pe59__lane28_strm1_cntl       ),      
               .std__pe59__lane28_strm1_data          ( std__pe59__lane28_strm1_data       ),      
               .std__pe59__lane28_strm1_data_valid    ( std__pe59__lane28_strm1_data_valid ),      
               .std__pe59__lane28_strm1_data_mask     ( std__pe59__lane28_strm1_data_mask  ),      

               // PE 59, Lane 29                 
               .pe59__std__lane29_strm0_ready         ( pe59__std__lane29_strm0_ready      ),      
               .std__pe59__lane29_strm0_cntl          ( std__pe59__lane29_strm0_cntl       ),      
               .std__pe59__lane29_strm0_data          ( std__pe59__lane29_strm0_data       ),      
               .std__pe59__lane29_strm0_data_valid    ( std__pe59__lane29_strm0_data_valid ),      
               .std__pe59__lane29_strm0_data_mask     ( std__pe59__lane29_strm0_data_mask  ),      

               .pe59__std__lane29_strm1_ready         ( pe59__std__lane29_strm1_ready      ),      
               .std__pe59__lane29_strm1_cntl          ( std__pe59__lane29_strm1_cntl       ),      
               .std__pe59__lane29_strm1_data          ( std__pe59__lane29_strm1_data       ),      
               .std__pe59__lane29_strm1_data_valid    ( std__pe59__lane29_strm1_data_valid ),      
               .std__pe59__lane29_strm1_data_mask     ( std__pe59__lane29_strm1_data_mask  ),      

               // PE 59, Lane 30                 
               .pe59__std__lane30_strm0_ready         ( pe59__std__lane30_strm0_ready      ),      
               .std__pe59__lane30_strm0_cntl          ( std__pe59__lane30_strm0_cntl       ),      
               .std__pe59__lane30_strm0_data          ( std__pe59__lane30_strm0_data       ),      
               .std__pe59__lane30_strm0_data_valid    ( std__pe59__lane30_strm0_data_valid ),      
               .std__pe59__lane30_strm0_data_mask     ( std__pe59__lane30_strm0_data_mask  ),      

               .pe59__std__lane30_strm1_ready         ( pe59__std__lane30_strm1_ready      ),      
               .std__pe59__lane30_strm1_cntl          ( std__pe59__lane30_strm1_cntl       ),      
               .std__pe59__lane30_strm1_data          ( std__pe59__lane30_strm1_data       ),      
               .std__pe59__lane30_strm1_data_valid    ( std__pe59__lane30_strm1_data_valid ),      
               .std__pe59__lane30_strm1_data_mask     ( std__pe59__lane30_strm1_data_mask  ),      

               // PE 59, Lane 31                 
               .pe59__std__lane31_strm0_ready         ( pe59__std__lane31_strm0_ready      ),      
               .std__pe59__lane31_strm0_cntl          ( std__pe59__lane31_strm0_cntl       ),      
               .std__pe59__lane31_strm0_data          ( std__pe59__lane31_strm0_data       ),      
               .std__pe59__lane31_strm0_data_valid    ( std__pe59__lane31_strm0_data_valid ),      
               .std__pe59__lane31_strm0_data_mask     ( std__pe59__lane31_strm0_data_mask  ),      

               .pe59__std__lane31_strm1_ready         ( pe59__std__lane31_strm1_ready      ),      
               .std__pe59__lane31_strm1_cntl          ( std__pe59__lane31_strm1_cntl       ),      
               .std__pe59__lane31_strm1_data          ( std__pe59__lane31_strm1_data       ),      
               .std__pe59__lane31_strm1_data_valid    ( std__pe59__lane31_strm1_data_valid ),      
               .std__pe59__lane31_strm1_data_mask     ( std__pe59__lane31_strm1_data_mask  ),      

               // PE 60, Lane 0                 
               .pe60__std__lane0_strm0_ready         ( pe60__std__lane0_strm0_ready      ),      
               .std__pe60__lane0_strm0_cntl          ( std__pe60__lane0_strm0_cntl       ),      
               .std__pe60__lane0_strm0_data          ( std__pe60__lane0_strm0_data       ),      
               .std__pe60__lane0_strm0_data_valid    ( std__pe60__lane0_strm0_data_valid ),      
               .std__pe60__lane0_strm0_data_mask     ( std__pe60__lane0_strm0_data_mask  ),      

               .pe60__std__lane0_strm1_ready         ( pe60__std__lane0_strm1_ready      ),      
               .std__pe60__lane0_strm1_cntl          ( std__pe60__lane0_strm1_cntl       ),      
               .std__pe60__lane0_strm1_data          ( std__pe60__lane0_strm1_data       ),      
               .std__pe60__lane0_strm1_data_valid    ( std__pe60__lane0_strm1_data_valid ),      
               .std__pe60__lane0_strm1_data_mask     ( std__pe60__lane0_strm1_data_mask  ),      

               // PE 60, Lane 1                 
               .pe60__std__lane1_strm0_ready         ( pe60__std__lane1_strm0_ready      ),      
               .std__pe60__lane1_strm0_cntl          ( std__pe60__lane1_strm0_cntl       ),      
               .std__pe60__lane1_strm0_data          ( std__pe60__lane1_strm0_data       ),      
               .std__pe60__lane1_strm0_data_valid    ( std__pe60__lane1_strm0_data_valid ),      
               .std__pe60__lane1_strm0_data_mask     ( std__pe60__lane1_strm0_data_mask  ),      

               .pe60__std__lane1_strm1_ready         ( pe60__std__lane1_strm1_ready      ),      
               .std__pe60__lane1_strm1_cntl          ( std__pe60__lane1_strm1_cntl       ),      
               .std__pe60__lane1_strm1_data          ( std__pe60__lane1_strm1_data       ),      
               .std__pe60__lane1_strm1_data_valid    ( std__pe60__lane1_strm1_data_valid ),      
               .std__pe60__lane1_strm1_data_mask     ( std__pe60__lane1_strm1_data_mask  ),      

               // PE 60, Lane 2                 
               .pe60__std__lane2_strm0_ready         ( pe60__std__lane2_strm0_ready      ),      
               .std__pe60__lane2_strm0_cntl          ( std__pe60__lane2_strm0_cntl       ),      
               .std__pe60__lane2_strm0_data          ( std__pe60__lane2_strm0_data       ),      
               .std__pe60__lane2_strm0_data_valid    ( std__pe60__lane2_strm0_data_valid ),      
               .std__pe60__lane2_strm0_data_mask     ( std__pe60__lane2_strm0_data_mask  ),      

               .pe60__std__lane2_strm1_ready         ( pe60__std__lane2_strm1_ready      ),      
               .std__pe60__lane2_strm1_cntl          ( std__pe60__lane2_strm1_cntl       ),      
               .std__pe60__lane2_strm1_data          ( std__pe60__lane2_strm1_data       ),      
               .std__pe60__lane2_strm1_data_valid    ( std__pe60__lane2_strm1_data_valid ),      
               .std__pe60__lane2_strm1_data_mask     ( std__pe60__lane2_strm1_data_mask  ),      

               // PE 60, Lane 3                 
               .pe60__std__lane3_strm0_ready         ( pe60__std__lane3_strm0_ready      ),      
               .std__pe60__lane3_strm0_cntl          ( std__pe60__lane3_strm0_cntl       ),      
               .std__pe60__lane3_strm0_data          ( std__pe60__lane3_strm0_data       ),      
               .std__pe60__lane3_strm0_data_valid    ( std__pe60__lane3_strm0_data_valid ),      
               .std__pe60__lane3_strm0_data_mask     ( std__pe60__lane3_strm0_data_mask  ),      

               .pe60__std__lane3_strm1_ready         ( pe60__std__lane3_strm1_ready      ),      
               .std__pe60__lane3_strm1_cntl          ( std__pe60__lane3_strm1_cntl       ),      
               .std__pe60__lane3_strm1_data          ( std__pe60__lane3_strm1_data       ),      
               .std__pe60__lane3_strm1_data_valid    ( std__pe60__lane3_strm1_data_valid ),      
               .std__pe60__lane3_strm1_data_mask     ( std__pe60__lane3_strm1_data_mask  ),      

               // PE 60, Lane 4                 
               .pe60__std__lane4_strm0_ready         ( pe60__std__lane4_strm0_ready      ),      
               .std__pe60__lane4_strm0_cntl          ( std__pe60__lane4_strm0_cntl       ),      
               .std__pe60__lane4_strm0_data          ( std__pe60__lane4_strm0_data       ),      
               .std__pe60__lane4_strm0_data_valid    ( std__pe60__lane4_strm0_data_valid ),      
               .std__pe60__lane4_strm0_data_mask     ( std__pe60__lane4_strm0_data_mask  ),      

               .pe60__std__lane4_strm1_ready         ( pe60__std__lane4_strm1_ready      ),      
               .std__pe60__lane4_strm1_cntl          ( std__pe60__lane4_strm1_cntl       ),      
               .std__pe60__lane4_strm1_data          ( std__pe60__lane4_strm1_data       ),      
               .std__pe60__lane4_strm1_data_valid    ( std__pe60__lane4_strm1_data_valid ),      
               .std__pe60__lane4_strm1_data_mask     ( std__pe60__lane4_strm1_data_mask  ),      

               // PE 60, Lane 5                 
               .pe60__std__lane5_strm0_ready         ( pe60__std__lane5_strm0_ready      ),      
               .std__pe60__lane5_strm0_cntl          ( std__pe60__lane5_strm0_cntl       ),      
               .std__pe60__lane5_strm0_data          ( std__pe60__lane5_strm0_data       ),      
               .std__pe60__lane5_strm0_data_valid    ( std__pe60__lane5_strm0_data_valid ),      
               .std__pe60__lane5_strm0_data_mask     ( std__pe60__lane5_strm0_data_mask  ),      

               .pe60__std__lane5_strm1_ready         ( pe60__std__lane5_strm1_ready      ),      
               .std__pe60__lane5_strm1_cntl          ( std__pe60__lane5_strm1_cntl       ),      
               .std__pe60__lane5_strm1_data          ( std__pe60__lane5_strm1_data       ),      
               .std__pe60__lane5_strm1_data_valid    ( std__pe60__lane5_strm1_data_valid ),      
               .std__pe60__lane5_strm1_data_mask     ( std__pe60__lane5_strm1_data_mask  ),      

               // PE 60, Lane 6                 
               .pe60__std__lane6_strm0_ready         ( pe60__std__lane6_strm0_ready      ),      
               .std__pe60__lane6_strm0_cntl          ( std__pe60__lane6_strm0_cntl       ),      
               .std__pe60__lane6_strm0_data          ( std__pe60__lane6_strm0_data       ),      
               .std__pe60__lane6_strm0_data_valid    ( std__pe60__lane6_strm0_data_valid ),      
               .std__pe60__lane6_strm0_data_mask     ( std__pe60__lane6_strm0_data_mask  ),      

               .pe60__std__lane6_strm1_ready         ( pe60__std__lane6_strm1_ready      ),      
               .std__pe60__lane6_strm1_cntl          ( std__pe60__lane6_strm1_cntl       ),      
               .std__pe60__lane6_strm1_data          ( std__pe60__lane6_strm1_data       ),      
               .std__pe60__lane6_strm1_data_valid    ( std__pe60__lane6_strm1_data_valid ),      
               .std__pe60__lane6_strm1_data_mask     ( std__pe60__lane6_strm1_data_mask  ),      

               // PE 60, Lane 7                 
               .pe60__std__lane7_strm0_ready         ( pe60__std__lane7_strm0_ready      ),      
               .std__pe60__lane7_strm0_cntl          ( std__pe60__lane7_strm0_cntl       ),      
               .std__pe60__lane7_strm0_data          ( std__pe60__lane7_strm0_data       ),      
               .std__pe60__lane7_strm0_data_valid    ( std__pe60__lane7_strm0_data_valid ),      
               .std__pe60__lane7_strm0_data_mask     ( std__pe60__lane7_strm0_data_mask  ),      

               .pe60__std__lane7_strm1_ready         ( pe60__std__lane7_strm1_ready      ),      
               .std__pe60__lane7_strm1_cntl          ( std__pe60__lane7_strm1_cntl       ),      
               .std__pe60__lane7_strm1_data          ( std__pe60__lane7_strm1_data       ),      
               .std__pe60__lane7_strm1_data_valid    ( std__pe60__lane7_strm1_data_valid ),      
               .std__pe60__lane7_strm1_data_mask     ( std__pe60__lane7_strm1_data_mask  ),      

               // PE 60, Lane 8                 
               .pe60__std__lane8_strm0_ready         ( pe60__std__lane8_strm0_ready      ),      
               .std__pe60__lane8_strm0_cntl          ( std__pe60__lane8_strm0_cntl       ),      
               .std__pe60__lane8_strm0_data          ( std__pe60__lane8_strm0_data       ),      
               .std__pe60__lane8_strm0_data_valid    ( std__pe60__lane8_strm0_data_valid ),      
               .std__pe60__lane8_strm0_data_mask     ( std__pe60__lane8_strm0_data_mask  ),      

               .pe60__std__lane8_strm1_ready         ( pe60__std__lane8_strm1_ready      ),      
               .std__pe60__lane8_strm1_cntl          ( std__pe60__lane8_strm1_cntl       ),      
               .std__pe60__lane8_strm1_data          ( std__pe60__lane8_strm1_data       ),      
               .std__pe60__lane8_strm1_data_valid    ( std__pe60__lane8_strm1_data_valid ),      
               .std__pe60__lane8_strm1_data_mask     ( std__pe60__lane8_strm1_data_mask  ),      

               // PE 60, Lane 9                 
               .pe60__std__lane9_strm0_ready         ( pe60__std__lane9_strm0_ready      ),      
               .std__pe60__lane9_strm0_cntl          ( std__pe60__lane9_strm0_cntl       ),      
               .std__pe60__lane9_strm0_data          ( std__pe60__lane9_strm0_data       ),      
               .std__pe60__lane9_strm0_data_valid    ( std__pe60__lane9_strm0_data_valid ),      
               .std__pe60__lane9_strm0_data_mask     ( std__pe60__lane9_strm0_data_mask  ),      

               .pe60__std__lane9_strm1_ready         ( pe60__std__lane9_strm1_ready      ),      
               .std__pe60__lane9_strm1_cntl          ( std__pe60__lane9_strm1_cntl       ),      
               .std__pe60__lane9_strm1_data          ( std__pe60__lane9_strm1_data       ),      
               .std__pe60__lane9_strm1_data_valid    ( std__pe60__lane9_strm1_data_valid ),      
               .std__pe60__lane9_strm1_data_mask     ( std__pe60__lane9_strm1_data_mask  ),      

               // PE 60, Lane 10                 
               .pe60__std__lane10_strm0_ready         ( pe60__std__lane10_strm0_ready      ),      
               .std__pe60__lane10_strm0_cntl          ( std__pe60__lane10_strm0_cntl       ),      
               .std__pe60__lane10_strm0_data          ( std__pe60__lane10_strm0_data       ),      
               .std__pe60__lane10_strm0_data_valid    ( std__pe60__lane10_strm0_data_valid ),      
               .std__pe60__lane10_strm0_data_mask     ( std__pe60__lane10_strm0_data_mask  ),      

               .pe60__std__lane10_strm1_ready         ( pe60__std__lane10_strm1_ready      ),      
               .std__pe60__lane10_strm1_cntl          ( std__pe60__lane10_strm1_cntl       ),      
               .std__pe60__lane10_strm1_data          ( std__pe60__lane10_strm1_data       ),      
               .std__pe60__lane10_strm1_data_valid    ( std__pe60__lane10_strm1_data_valid ),      
               .std__pe60__lane10_strm1_data_mask     ( std__pe60__lane10_strm1_data_mask  ),      

               // PE 60, Lane 11                 
               .pe60__std__lane11_strm0_ready         ( pe60__std__lane11_strm0_ready      ),      
               .std__pe60__lane11_strm0_cntl          ( std__pe60__lane11_strm0_cntl       ),      
               .std__pe60__lane11_strm0_data          ( std__pe60__lane11_strm0_data       ),      
               .std__pe60__lane11_strm0_data_valid    ( std__pe60__lane11_strm0_data_valid ),      
               .std__pe60__lane11_strm0_data_mask     ( std__pe60__lane11_strm0_data_mask  ),      

               .pe60__std__lane11_strm1_ready         ( pe60__std__lane11_strm1_ready      ),      
               .std__pe60__lane11_strm1_cntl          ( std__pe60__lane11_strm1_cntl       ),      
               .std__pe60__lane11_strm1_data          ( std__pe60__lane11_strm1_data       ),      
               .std__pe60__lane11_strm1_data_valid    ( std__pe60__lane11_strm1_data_valid ),      
               .std__pe60__lane11_strm1_data_mask     ( std__pe60__lane11_strm1_data_mask  ),      

               // PE 60, Lane 12                 
               .pe60__std__lane12_strm0_ready         ( pe60__std__lane12_strm0_ready      ),      
               .std__pe60__lane12_strm0_cntl          ( std__pe60__lane12_strm0_cntl       ),      
               .std__pe60__lane12_strm0_data          ( std__pe60__lane12_strm0_data       ),      
               .std__pe60__lane12_strm0_data_valid    ( std__pe60__lane12_strm0_data_valid ),      
               .std__pe60__lane12_strm0_data_mask     ( std__pe60__lane12_strm0_data_mask  ),      

               .pe60__std__lane12_strm1_ready         ( pe60__std__lane12_strm1_ready      ),      
               .std__pe60__lane12_strm1_cntl          ( std__pe60__lane12_strm1_cntl       ),      
               .std__pe60__lane12_strm1_data          ( std__pe60__lane12_strm1_data       ),      
               .std__pe60__lane12_strm1_data_valid    ( std__pe60__lane12_strm1_data_valid ),      
               .std__pe60__lane12_strm1_data_mask     ( std__pe60__lane12_strm1_data_mask  ),      

               // PE 60, Lane 13                 
               .pe60__std__lane13_strm0_ready         ( pe60__std__lane13_strm0_ready      ),      
               .std__pe60__lane13_strm0_cntl          ( std__pe60__lane13_strm0_cntl       ),      
               .std__pe60__lane13_strm0_data          ( std__pe60__lane13_strm0_data       ),      
               .std__pe60__lane13_strm0_data_valid    ( std__pe60__lane13_strm0_data_valid ),      
               .std__pe60__lane13_strm0_data_mask     ( std__pe60__lane13_strm0_data_mask  ),      

               .pe60__std__lane13_strm1_ready         ( pe60__std__lane13_strm1_ready      ),      
               .std__pe60__lane13_strm1_cntl          ( std__pe60__lane13_strm1_cntl       ),      
               .std__pe60__lane13_strm1_data          ( std__pe60__lane13_strm1_data       ),      
               .std__pe60__lane13_strm1_data_valid    ( std__pe60__lane13_strm1_data_valid ),      
               .std__pe60__lane13_strm1_data_mask     ( std__pe60__lane13_strm1_data_mask  ),      

               // PE 60, Lane 14                 
               .pe60__std__lane14_strm0_ready         ( pe60__std__lane14_strm0_ready      ),      
               .std__pe60__lane14_strm0_cntl          ( std__pe60__lane14_strm0_cntl       ),      
               .std__pe60__lane14_strm0_data          ( std__pe60__lane14_strm0_data       ),      
               .std__pe60__lane14_strm0_data_valid    ( std__pe60__lane14_strm0_data_valid ),      
               .std__pe60__lane14_strm0_data_mask     ( std__pe60__lane14_strm0_data_mask  ),      

               .pe60__std__lane14_strm1_ready         ( pe60__std__lane14_strm1_ready      ),      
               .std__pe60__lane14_strm1_cntl          ( std__pe60__lane14_strm1_cntl       ),      
               .std__pe60__lane14_strm1_data          ( std__pe60__lane14_strm1_data       ),      
               .std__pe60__lane14_strm1_data_valid    ( std__pe60__lane14_strm1_data_valid ),      
               .std__pe60__lane14_strm1_data_mask     ( std__pe60__lane14_strm1_data_mask  ),      

               // PE 60, Lane 15                 
               .pe60__std__lane15_strm0_ready         ( pe60__std__lane15_strm0_ready      ),      
               .std__pe60__lane15_strm0_cntl          ( std__pe60__lane15_strm0_cntl       ),      
               .std__pe60__lane15_strm0_data          ( std__pe60__lane15_strm0_data       ),      
               .std__pe60__lane15_strm0_data_valid    ( std__pe60__lane15_strm0_data_valid ),      
               .std__pe60__lane15_strm0_data_mask     ( std__pe60__lane15_strm0_data_mask  ),      

               .pe60__std__lane15_strm1_ready         ( pe60__std__lane15_strm1_ready      ),      
               .std__pe60__lane15_strm1_cntl          ( std__pe60__lane15_strm1_cntl       ),      
               .std__pe60__lane15_strm1_data          ( std__pe60__lane15_strm1_data       ),      
               .std__pe60__lane15_strm1_data_valid    ( std__pe60__lane15_strm1_data_valid ),      
               .std__pe60__lane15_strm1_data_mask     ( std__pe60__lane15_strm1_data_mask  ),      

               // PE 60, Lane 16                 
               .pe60__std__lane16_strm0_ready         ( pe60__std__lane16_strm0_ready      ),      
               .std__pe60__lane16_strm0_cntl          ( std__pe60__lane16_strm0_cntl       ),      
               .std__pe60__lane16_strm0_data          ( std__pe60__lane16_strm0_data       ),      
               .std__pe60__lane16_strm0_data_valid    ( std__pe60__lane16_strm0_data_valid ),      
               .std__pe60__lane16_strm0_data_mask     ( std__pe60__lane16_strm0_data_mask  ),      

               .pe60__std__lane16_strm1_ready         ( pe60__std__lane16_strm1_ready      ),      
               .std__pe60__lane16_strm1_cntl          ( std__pe60__lane16_strm1_cntl       ),      
               .std__pe60__lane16_strm1_data          ( std__pe60__lane16_strm1_data       ),      
               .std__pe60__lane16_strm1_data_valid    ( std__pe60__lane16_strm1_data_valid ),      
               .std__pe60__lane16_strm1_data_mask     ( std__pe60__lane16_strm1_data_mask  ),      

               // PE 60, Lane 17                 
               .pe60__std__lane17_strm0_ready         ( pe60__std__lane17_strm0_ready      ),      
               .std__pe60__lane17_strm0_cntl          ( std__pe60__lane17_strm0_cntl       ),      
               .std__pe60__lane17_strm0_data          ( std__pe60__lane17_strm0_data       ),      
               .std__pe60__lane17_strm0_data_valid    ( std__pe60__lane17_strm0_data_valid ),      
               .std__pe60__lane17_strm0_data_mask     ( std__pe60__lane17_strm0_data_mask  ),      

               .pe60__std__lane17_strm1_ready         ( pe60__std__lane17_strm1_ready      ),      
               .std__pe60__lane17_strm1_cntl          ( std__pe60__lane17_strm1_cntl       ),      
               .std__pe60__lane17_strm1_data          ( std__pe60__lane17_strm1_data       ),      
               .std__pe60__lane17_strm1_data_valid    ( std__pe60__lane17_strm1_data_valid ),      
               .std__pe60__lane17_strm1_data_mask     ( std__pe60__lane17_strm1_data_mask  ),      

               // PE 60, Lane 18                 
               .pe60__std__lane18_strm0_ready         ( pe60__std__lane18_strm0_ready      ),      
               .std__pe60__lane18_strm0_cntl          ( std__pe60__lane18_strm0_cntl       ),      
               .std__pe60__lane18_strm0_data          ( std__pe60__lane18_strm0_data       ),      
               .std__pe60__lane18_strm0_data_valid    ( std__pe60__lane18_strm0_data_valid ),      
               .std__pe60__lane18_strm0_data_mask     ( std__pe60__lane18_strm0_data_mask  ),      

               .pe60__std__lane18_strm1_ready         ( pe60__std__lane18_strm1_ready      ),      
               .std__pe60__lane18_strm1_cntl          ( std__pe60__lane18_strm1_cntl       ),      
               .std__pe60__lane18_strm1_data          ( std__pe60__lane18_strm1_data       ),      
               .std__pe60__lane18_strm1_data_valid    ( std__pe60__lane18_strm1_data_valid ),      
               .std__pe60__lane18_strm1_data_mask     ( std__pe60__lane18_strm1_data_mask  ),      

               // PE 60, Lane 19                 
               .pe60__std__lane19_strm0_ready         ( pe60__std__lane19_strm0_ready      ),      
               .std__pe60__lane19_strm0_cntl          ( std__pe60__lane19_strm0_cntl       ),      
               .std__pe60__lane19_strm0_data          ( std__pe60__lane19_strm0_data       ),      
               .std__pe60__lane19_strm0_data_valid    ( std__pe60__lane19_strm0_data_valid ),      
               .std__pe60__lane19_strm0_data_mask     ( std__pe60__lane19_strm0_data_mask  ),      

               .pe60__std__lane19_strm1_ready         ( pe60__std__lane19_strm1_ready      ),      
               .std__pe60__lane19_strm1_cntl          ( std__pe60__lane19_strm1_cntl       ),      
               .std__pe60__lane19_strm1_data          ( std__pe60__lane19_strm1_data       ),      
               .std__pe60__lane19_strm1_data_valid    ( std__pe60__lane19_strm1_data_valid ),      
               .std__pe60__lane19_strm1_data_mask     ( std__pe60__lane19_strm1_data_mask  ),      

               // PE 60, Lane 20                 
               .pe60__std__lane20_strm0_ready         ( pe60__std__lane20_strm0_ready      ),      
               .std__pe60__lane20_strm0_cntl          ( std__pe60__lane20_strm0_cntl       ),      
               .std__pe60__lane20_strm0_data          ( std__pe60__lane20_strm0_data       ),      
               .std__pe60__lane20_strm0_data_valid    ( std__pe60__lane20_strm0_data_valid ),      
               .std__pe60__lane20_strm0_data_mask     ( std__pe60__lane20_strm0_data_mask  ),      

               .pe60__std__lane20_strm1_ready         ( pe60__std__lane20_strm1_ready      ),      
               .std__pe60__lane20_strm1_cntl          ( std__pe60__lane20_strm1_cntl       ),      
               .std__pe60__lane20_strm1_data          ( std__pe60__lane20_strm1_data       ),      
               .std__pe60__lane20_strm1_data_valid    ( std__pe60__lane20_strm1_data_valid ),      
               .std__pe60__lane20_strm1_data_mask     ( std__pe60__lane20_strm1_data_mask  ),      

               // PE 60, Lane 21                 
               .pe60__std__lane21_strm0_ready         ( pe60__std__lane21_strm0_ready      ),      
               .std__pe60__lane21_strm0_cntl          ( std__pe60__lane21_strm0_cntl       ),      
               .std__pe60__lane21_strm0_data          ( std__pe60__lane21_strm0_data       ),      
               .std__pe60__lane21_strm0_data_valid    ( std__pe60__lane21_strm0_data_valid ),      
               .std__pe60__lane21_strm0_data_mask     ( std__pe60__lane21_strm0_data_mask  ),      

               .pe60__std__lane21_strm1_ready         ( pe60__std__lane21_strm1_ready      ),      
               .std__pe60__lane21_strm1_cntl          ( std__pe60__lane21_strm1_cntl       ),      
               .std__pe60__lane21_strm1_data          ( std__pe60__lane21_strm1_data       ),      
               .std__pe60__lane21_strm1_data_valid    ( std__pe60__lane21_strm1_data_valid ),      
               .std__pe60__lane21_strm1_data_mask     ( std__pe60__lane21_strm1_data_mask  ),      

               // PE 60, Lane 22                 
               .pe60__std__lane22_strm0_ready         ( pe60__std__lane22_strm0_ready      ),      
               .std__pe60__lane22_strm0_cntl          ( std__pe60__lane22_strm0_cntl       ),      
               .std__pe60__lane22_strm0_data          ( std__pe60__lane22_strm0_data       ),      
               .std__pe60__lane22_strm0_data_valid    ( std__pe60__lane22_strm0_data_valid ),      
               .std__pe60__lane22_strm0_data_mask     ( std__pe60__lane22_strm0_data_mask  ),      

               .pe60__std__lane22_strm1_ready         ( pe60__std__lane22_strm1_ready      ),      
               .std__pe60__lane22_strm1_cntl          ( std__pe60__lane22_strm1_cntl       ),      
               .std__pe60__lane22_strm1_data          ( std__pe60__lane22_strm1_data       ),      
               .std__pe60__lane22_strm1_data_valid    ( std__pe60__lane22_strm1_data_valid ),      
               .std__pe60__lane22_strm1_data_mask     ( std__pe60__lane22_strm1_data_mask  ),      

               // PE 60, Lane 23                 
               .pe60__std__lane23_strm0_ready         ( pe60__std__lane23_strm0_ready      ),      
               .std__pe60__lane23_strm0_cntl          ( std__pe60__lane23_strm0_cntl       ),      
               .std__pe60__lane23_strm0_data          ( std__pe60__lane23_strm0_data       ),      
               .std__pe60__lane23_strm0_data_valid    ( std__pe60__lane23_strm0_data_valid ),      
               .std__pe60__lane23_strm0_data_mask     ( std__pe60__lane23_strm0_data_mask  ),      

               .pe60__std__lane23_strm1_ready         ( pe60__std__lane23_strm1_ready      ),      
               .std__pe60__lane23_strm1_cntl          ( std__pe60__lane23_strm1_cntl       ),      
               .std__pe60__lane23_strm1_data          ( std__pe60__lane23_strm1_data       ),      
               .std__pe60__lane23_strm1_data_valid    ( std__pe60__lane23_strm1_data_valid ),      
               .std__pe60__lane23_strm1_data_mask     ( std__pe60__lane23_strm1_data_mask  ),      

               // PE 60, Lane 24                 
               .pe60__std__lane24_strm0_ready         ( pe60__std__lane24_strm0_ready      ),      
               .std__pe60__lane24_strm0_cntl          ( std__pe60__lane24_strm0_cntl       ),      
               .std__pe60__lane24_strm0_data          ( std__pe60__lane24_strm0_data       ),      
               .std__pe60__lane24_strm0_data_valid    ( std__pe60__lane24_strm0_data_valid ),      
               .std__pe60__lane24_strm0_data_mask     ( std__pe60__lane24_strm0_data_mask  ),      

               .pe60__std__lane24_strm1_ready         ( pe60__std__lane24_strm1_ready      ),      
               .std__pe60__lane24_strm1_cntl          ( std__pe60__lane24_strm1_cntl       ),      
               .std__pe60__lane24_strm1_data          ( std__pe60__lane24_strm1_data       ),      
               .std__pe60__lane24_strm1_data_valid    ( std__pe60__lane24_strm1_data_valid ),      
               .std__pe60__lane24_strm1_data_mask     ( std__pe60__lane24_strm1_data_mask  ),      

               // PE 60, Lane 25                 
               .pe60__std__lane25_strm0_ready         ( pe60__std__lane25_strm0_ready      ),      
               .std__pe60__lane25_strm0_cntl          ( std__pe60__lane25_strm0_cntl       ),      
               .std__pe60__lane25_strm0_data          ( std__pe60__lane25_strm0_data       ),      
               .std__pe60__lane25_strm0_data_valid    ( std__pe60__lane25_strm0_data_valid ),      
               .std__pe60__lane25_strm0_data_mask     ( std__pe60__lane25_strm0_data_mask  ),      

               .pe60__std__lane25_strm1_ready         ( pe60__std__lane25_strm1_ready      ),      
               .std__pe60__lane25_strm1_cntl          ( std__pe60__lane25_strm1_cntl       ),      
               .std__pe60__lane25_strm1_data          ( std__pe60__lane25_strm1_data       ),      
               .std__pe60__lane25_strm1_data_valid    ( std__pe60__lane25_strm1_data_valid ),      
               .std__pe60__lane25_strm1_data_mask     ( std__pe60__lane25_strm1_data_mask  ),      

               // PE 60, Lane 26                 
               .pe60__std__lane26_strm0_ready         ( pe60__std__lane26_strm0_ready      ),      
               .std__pe60__lane26_strm0_cntl          ( std__pe60__lane26_strm0_cntl       ),      
               .std__pe60__lane26_strm0_data          ( std__pe60__lane26_strm0_data       ),      
               .std__pe60__lane26_strm0_data_valid    ( std__pe60__lane26_strm0_data_valid ),      
               .std__pe60__lane26_strm0_data_mask     ( std__pe60__lane26_strm0_data_mask  ),      

               .pe60__std__lane26_strm1_ready         ( pe60__std__lane26_strm1_ready      ),      
               .std__pe60__lane26_strm1_cntl          ( std__pe60__lane26_strm1_cntl       ),      
               .std__pe60__lane26_strm1_data          ( std__pe60__lane26_strm1_data       ),      
               .std__pe60__lane26_strm1_data_valid    ( std__pe60__lane26_strm1_data_valid ),      
               .std__pe60__lane26_strm1_data_mask     ( std__pe60__lane26_strm1_data_mask  ),      

               // PE 60, Lane 27                 
               .pe60__std__lane27_strm0_ready         ( pe60__std__lane27_strm0_ready      ),      
               .std__pe60__lane27_strm0_cntl          ( std__pe60__lane27_strm0_cntl       ),      
               .std__pe60__lane27_strm0_data          ( std__pe60__lane27_strm0_data       ),      
               .std__pe60__lane27_strm0_data_valid    ( std__pe60__lane27_strm0_data_valid ),      
               .std__pe60__lane27_strm0_data_mask     ( std__pe60__lane27_strm0_data_mask  ),      

               .pe60__std__lane27_strm1_ready         ( pe60__std__lane27_strm1_ready      ),      
               .std__pe60__lane27_strm1_cntl          ( std__pe60__lane27_strm1_cntl       ),      
               .std__pe60__lane27_strm1_data          ( std__pe60__lane27_strm1_data       ),      
               .std__pe60__lane27_strm1_data_valid    ( std__pe60__lane27_strm1_data_valid ),      
               .std__pe60__lane27_strm1_data_mask     ( std__pe60__lane27_strm1_data_mask  ),      

               // PE 60, Lane 28                 
               .pe60__std__lane28_strm0_ready         ( pe60__std__lane28_strm0_ready      ),      
               .std__pe60__lane28_strm0_cntl          ( std__pe60__lane28_strm0_cntl       ),      
               .std__pe60__lane28_strm0_data          ( std__pe60__lane28_strm0_data       ),      
               .std__pe60__lane28_strm0_data_valid    ( std__pe60__lane28_strm0_data_valid ),      
               .std__pe60__lane28_strm0_data_mask     ( std__pe60__lane28_strm0_data_mask  ),      

               .pe60__std__lane28_strm1_ready         ( pe60__std__lane28_strm1_ready      ),      
               .std__pe60__lane28_strm1_cntl          ( std__pe60__lane28_strm1_cntl       ),      
               .std__pe60__lane28_strm1_data          ( std__pe60__lane28_strm1_data       ),      
               .std__pe60__lane28_strm1_data_valid    ( std__pe60__lane28_strm1_data_valid ),      
               .std__pe60__lane28_strm1_data_mask     ( std__pe60__lane28_strm1_data_mask  ),      

               // PE 60, Lane 29                 
               .pe60__std__lane29_strm0_ready         ( pe60__std__lane29_strm0_ready      ),      
               .std__pe60__lane29_strm0_cntl          ( std__pe60__lane29_strm0_cntl       ),      
               .std__pe60__lane29_strm0_data          ( std__pe60__lane29_strm0_data       ),      
               .std__pe60__lane29_strm0_data_valid    ( std__pe60__lane29_strm0_data_valid ),      
               .std__pe60__lane29_strm0_data_mask     ( std__pe60__lane29_strm0_data_mask  ),      

               .pe60__std__lane29_strm1_ready         ( pe60__std__lane29_strm1_ready      ),      
               .std__pe60__lane29_strm1_cntl          ( std__pe60__lane29_strm1_cntl       ),      
               .std__pe60__lane29_strm1_data          ( std__pe60__lane29_strm1_data       ),      
               .std__pe60__lane29_strm1_data_valid    ( std__pe60__lane29_strm1_data_valid ),      
               .std__pe60__lane29_strm1_data_mask     ( std__pe60__lane29_strm1_data_mask  ),      

               // PE 60, Lane 30                 
               .pe60__std__lane30_strm0_ready         ( pe60__std__lane30_strm0_ready      ),      
               .std__pe60__lane30_strm0_cntl          ( std__pe60__lane30_strm0_cntl       ),      
               .std__pe60__lane30_strm0_data          ( std__pe60__lane30_strm0_data       ),      
               .std__pe60__lane30_strm0_data_valid    ( std__pe60__lane30_strm0_data_valid ),      
               .std__pe60__lane30_strm0_data_mask     ( std__pe60__lane30_strm0_data_mask  ),      

               .pe60__std__lane30_strm1_ready         ( pe60__std__lane30_strm1_ready      ),      
               .std__pe60__lane30_strm1_cntl          ( std__pe60__lane30_strm1_cntl       ),      
               .std__pe60__lane30_strm1_data          ( std__pe60__lane30_strm1_data       ),      
               .std__pe60__lane30_strm1_data_valid    ( std__pe60__lane30_strm1_data_valid ),      
               .std__pe60__lane30_strm1_data_mask     ( std__pe60__lane30_strm1_data_mask  ),      

               // PE 60, Lane 31                 
               .pe60__std__lane31_strm0_ready         ( pe60__std__lane31_strm0_ready      ),      
               .std__pe60__lane31_strm0_cntl          ( std__pe60__lane31_strm0_cntl       ),      
               .std__pe60__lane31_strm0_data          ( std__pe60__lane31_strm0_data       ),      
               .std__pe60__lane31_strm0_data_valid    ( std__pe60__lane31_strm0_data_valid ),      
               .std__pe60__lane31_strm0_data_mask     ( std__pe60__lane31_strm0_data_mask  ),      

               .pe60__std__lane31_strm1_ready         ( pe60__std__lane31_strm1_ready      ),      
               .std__pe60__lane31_strm1_cntl          ( std__pe60__lane31_strm1_cntl       ),      
               .std__pe60__lane31_strm1_data          ( std__pe60__lane31_strm1_data       ),      
               .std__pe60__lane31_strm1_data_valid    ( std__pe60__lane31_strm1_data_valid ),      
               .std__pe60__lane31_strm1_data_mask     ( std__pe60__lane31_strm1_data_mask  ),      

               // PE 61, Lane 0                 
               .pe61__std__lane0_strm0_ready         ( pe61__std__lane0_strm0_ready      ),      
               .std__pe61__lane0_strm0_cntl          ( std__pe61__lane0_strm0_cntl       ),      
               .std__pe61__lane0_strm0_data          ( std__pe61__lane0_strm0_data       ),      
               .std__pe61__lane0_strm0_data_valid    ( std__pe61__lane0_strm0_data_valid ),      
               .std__pe61__lane0_strm0_data_mask     ( std__pe61__lane0_strm0_data_mask  ),      

               .pe61__std__lane0_strm1_ready         ( pe61__std__lane0_strm1_ready      ),      
               .std__pe61__lane0_strm1_cntl          ( std__pe61__lane0_strm1_cntl       ),      
               .std__pe61__lane0_strm1_data          ( std__pe61__lane0_strm1_data       ),      
               .std__pe61__lane0_strm1_data_valid    ( std__pe61__lane0_strm1_data_valid ),      
               .std__pe61__lane0_strm1_data_mask     ( std__pe61__lane0_strm1_data_mask  ),      

               // PE 61, Lane 1                 
               .pe61__std__lane1_strm0_ready         ( pe61__std__lane1_strm0_ready      ),      
               .std__pe61__lane1_strm0_cntl          ( std__pe61__lane1_strm0_cntl       ),      
               .std__pe61__lane1_strm0_data          ( std__pe61__lane1_strm0_data       ),      
               .std__pe61__lane1_strm0_data_valid    ( std__pe61__lane1_strm0_data_valid ),      
               .std__pe61__lane1_strm0_data_mask     ( std__pe61__lane1_strm0_data_mask  ),      

               .pe61__std__lane1_strm1_ready         ( pe61__std__lane1_strm1_ready      ),      
               .std__pe61__lane1_strm1_cntl          ( std__pe61__lane1_strm1_cntl       ),      
               .std__pe61__lane1_strm1_data          ( std__pe61__lane1_strm1_data       ),      
               .std__pe61__lane1_strm1_data_valid    ( std__pe61__lane1_strm1_data_valid ),      
               .std__pe61__lane1_strm1_data_mask     ( std__pe61__lane1_strm1_data_mask  ),      

               // PE 61, Lane 2                 
               .pe61__std__lane2_strm0_ready         ( pe61__std__lane2_strm0_ready      ),      
               .std__pe61__lane2_strm0_cntl          ( std__pe61__lane2_strm0_cntl       ),      
               .std__pe61__lane2_strm0_data          ( std__pe61__lane2_strm0_data       ),      
               .std__pe61__lane2_strm0_data_valid    ( std__pe61__lane2_strm0_data_valid ),      
               .std__pe61__lane2_strm0_data_mask     ( std__pe61__lane2_strm0_data_mask  ),      

               .pe61__std__lane2_strm1_ready         ( pe61__std__lane2_strm1_ready      ),      
               .std__pe61__lane2_strm1_cntl          ( std__pe61__lane2_strm1_cntl       ),      
               .std__pe61__lane2_strm1_data          ( std__pe61__lane2_strm1_data       ),      
               .std__pe61__lane2_strm1_data_valid    ( std__pe61__lane2_strm1_data_valid ),      
               .std__pe61__lane2_strm1_data_mask     ( std__pe61__lane2_strm1_data_mask  ),      

               // PE 61, Lane 3                 
               .pe61__std__lane3_strm0_ready         ( pe61__std__lane3_strm0_ready      ),      
               .std__pe61__lane3_strm0_cntl          ( std__pe61__lane3_strm0_cntl       ),      
               .std__pe61__lane3_strm0_data          ( std__pe61__lane3_strm0_data       ),      
               .std__pe61__lane3_strm0_data_valid    ( std__pe61__lane3_strm0_data_valid ),      
               .std__pe61__lane3_strm0_data_mask     ( std__pe61__lane3_strm0_data_mask  ),      

               .pe61__std__lane3_strm1_ready         ( pe61__std__lane3_strm1_ready      ),      
               .std__pe61__lane3_strm1_cntl          ( std__pe61__lane3_strm1_cntl       ),      
               .std__pe61__lane3_strm1_data          ( std__pe61__lane3_strm1_data       ),      
               .std__pe61__lane3_strm1_data_valid    ( std__pe61__lane3_strm1_data_valid ),      
               .std__pe61__lane3_strm1_data_mask     ( std__pe61__lane3_strm1_data_mask  ),      

               // PE 61, Lane 4                 
               .pe61__std__lane4_strm0_ready         ( pe61__std__lane4_strm0_ready      ),      
               .std__pe61__lane4_strm0_cntl          ( std__pe61__lane4_strm0_cntl       ),      
               .std__pe61__lane4_strm0_data          ( std__pe61__lane4_strm0_data       ),      
               .std__pe61__lane4_strm0_data_valid    ( std__pe61__lane4_strm0_data_valid ),      
               .std__pe61__lane4_strm0_data_mask     ( std__pe61__lane4_strm0_data_mask  ),      

               .pe61__std__lane4_strm1_ready         ( pe61__std__lane4_strm1_ready      ),      
               .std__pe61__lane4_strm1_cntl          ( std__pe61__lane4_strm1_cntl       ),      
               .std__pe61__lane4_strm1_data          ( std__pe61__lane4_strm1_data       ),      
               .std__pe61__lane4_strm1_data_valid    ( std__pe61__lane4_strm1_data_valid ),      
               .std__pe61__lane4_strm1_data_mask     ( std__pe61__lane4_strm1_data_mask  ),      

               // PE 61, Lane 5                 
               .pe61__std__lane5_strm0_ready         ( pe61__std__lane5_strm0_ready      ),      
               .std__pe61__lane5_strm0_cntl          ( std__pe61__lane5_strm0_cntl       ),      
               .std__pe61__lane5_strm0_data          ( std__pe61__lane5_strm0_data       ),      
               .std__pe61__lane5_strm0_data_valid    ( std__pe61__lane5_strm0_data_valid ),      
               .std__pe61__lane5_strm0_data_mask     ( std__pe61__lane5_strm0_data_mask  ),      

               .pe61__std__lane5_strm1_ready         ( pe61__std__lane5_strm1_ready      ),      
               .std__pe61__lane5_strm1_cntl          ( std__pe61__lane5_strm1_cntl       ),      
               .std__pe61__lane5_strm1_data          ( std__pe61__lane5_strm1_data       ),      
               .std__pe61__lane5_strm1_data_valid    ( std__pe61__lane5_strm1_data_valid ),      
               .std__pe61__lane5_strm1_data_mask     ( std__pe61__lane5_strm1_data_mask  ),      

               // PE 61, Lane 6                 
               .pe61__std__lane6_strm0_ready         ( pe61__std__lane6_strm0_ready      ),      
               .std__pe61__lane6_strm0_cntl          ( std__pe61__lane6_strm0_cntl       ),      
               .std__pe61__lane6_strm0_data          ( std__pe61__lane6_strm0_data       ),      
               .std__pe61__lane6_strm0_data_valid    ( std__pe61__lane6_strm0_data_valid ),      
               .std__pe61__lane6_strm0_data_mask     ( std__pe61__lane6_strm0_data_mask  ),      

               .pe61__std__lane6_strm1_ready         ( pe61__std__lane6_strm1_ready      ),      
               .std__pe61__lane6_strm1_cntl          ( std__pe61__lane6_strm1_cntl       ),      
               .std__pe61__lane6_strm1_data          ( std__pe61__lane6_strm1_data       ),      
               .std__pe61__lane6_strm1_data_valid    ( std__pe61__lane6_strm1_data_valid ),      
               .std__pe61__lane6_strm1_data_mask     ( std__pe61__lane6_strm1_data_mask  ),      

               // PE 61, Lane 7                 
               .pe61__std__lane7_strm0_ready         ( pe61__std__lane7_strm0_ready      ),      
               .std__pe61__lane7_strm0_cntl          ( std__pe61__lane7_strm0_cntl       ),      
               .std__pe61__lane7_strm0_data          ( std__pe61__lane7_strm0_data       ),      
               .std__pe61__lane7_strm0_data_valid    ( std__pe61__lane7_strm0_data_valid ),      
               .std__pe61__lane7_strm0_data_mask     ( std__pe61__lane7_strm0_data_mask  ),      

               .pe61__std__lane7_strm1_ready         ( pe61__std__lane7_strm1_ready      ),      
               .std__pe61__lane7_strm1_cntl          ( std__pe61__lane7_strm1_cntl       ),      
               .std__pe61__lane7_strm1_data          ( std__pe61__lane7_strm1_data       ),      
               .std__pe61__lane7_strm1_data_valid    ( std__pe61__lane7_strm1_data_valid ),      
               .std__pe61__lane7_strm1_data_mask     ( std__pe61__lane7_strm1_data_mask  ),      

               // PE 61, Lane 8                 
               .pe61__std__lane8_strm0_ready         ( pe61__std__lane8_strm0_ready      ),      
               .std__pe61__lane8_strm0_cntl          ( std__pe61__lane8_strm0_cntl       ),      
               .std__pe61__lane8_strm0_data          ( std__pe61__lane8_strm0_data       ),      
               .std__pe61__lane8_strm0_data_valid    ( std__pe61__lane8_strm0_data_valid ),      
               .std__pe61__lane8_strm0_data_mask     ( std__pe61__lane8_strm0_data_mask  ),      

               .pe61__std__lane8_strm1_ready         ( pe61__std__lane8_strm1_ready      ),      
               .std__pe61__lane8_strm1_cntl          ( std__pe61__lane8_strm1_cntl       ),      
               .std__pe61__lane8_strm1_data          ( std__pe61__lane8_strm1_data       ),      
               .std__pe61__lane8_strm1_data_valid    ( std__pe61__lane8_strm1_data_valid ),      
               .std__pe61__lane8_strm1_data_mask     ( std__pe61__lane8_strm1_data_mask  ),      

               // PE 61, Lane 9                 
               .pe61__std__lane9_strm0_ready         ( pe61__std__lane9_strm0_ready      ),      
               .std__pe61__lane9_strm0_cntl          ( std__pe61__lane9_strm0_cntl       ),      
               .std__pe61__lane9_strm0_data          ( std__pe61__lane9_strm0_data       ),      
               .std__pe61__lane9_strm0_data_valid    ( std__pe61__lane9_strm0_data_valid ),      
               .std__pe61__lane9_strm0_data_mask     ( std__pe61__lane9_strm0_data_mask  ),      

               .pe61__std__lane9_strm1_ready         ( pe61__std__lane9_strm1_ready      ),      
               .std__pe61__lane9_strm1_cntl          ( std__pe61__lane9_strm1_cntl       ),      
               .std__pe61__lane9_strm1_data          ( std__pe61__lane9_strm1_data       ),      
               .std__pe61__lane9_strm1_data_valid    ( std__pe61__lane9_strm1_data_valid ),      
               .std__pe61__lane9_strm1_data_mask     ( std__pe61__lane9_strm1_data_mask  ),      

               // PE 61, Lane 10                 
               .pe61__std__lane10_strm0_ready         ( pe61__std__lane10_strm0_ready      ),      
               .std__pe61__lane10_strm0_cntl          ( std__pe61__lane10_strm0_cntl       ),      
               .std__pe61__lane10_strm0_data          ( std__pe61__lane10_strm0_data       ),      
               .std__pe61__lane10_strm0_data_valid    ( std__pe61__lane10_strm0_data_valid ),      
               .std__pe61__lane10_strm0_data_mask     ( std__pe61__lane10_strm0_data_mask  ),      

               .pe61__std__lane10_strm1_ready         ( pe61__std__lane10_strm1_ready      ),      
               .std__pe61__lane10_strm1_cntl          ( std__pe61__lane10_strm1_cntl       ),      
               .std__pe61__lane10_strm1_data          ( std__pe61__lane10_strm1_data       ),      
               .std__pe61__lane10_strm1_data_valid    ( std__pe61__lane10_strm1_data_valid ),      
               .std__pe61__lane10_strm1_data_mask     ( std__pe61__lane10_strm1_data_mask  ),      

               // PE 61, Lane 11                 
               .pe61__std__lane11_strm0_ready         ( pe61__std__lane11_strm0_ready      ),      
               .std__pe61__lane11_strm0_cntl          ( std__pe61__lane11_strm0_cntl       ),      
               .std__pe61__lane11_strm0_data          ( std__pe61__lane11_strm0_data       ),      
               .std__pe61__lane11_strm0_data_valid    ( std__pe61__lane11_strm0_data_valid ),      
               .std__pe61__lane11_strm0_data_mask     ( std__pe61__lane11_strm0_data_mask  ),      

               .pe61__std__lane11_strm1_ready         ( pe61__std__lane11_strm1_ready      ),      
               .std__pe61__lane11_strm1_cntl          ( std__pe61__lane11_strm1_cntl       ),      
               .std__pe61__lane11_strm1_data          ( std__pe61__lane11_strm1_data       ),      
               .std__pe61__lane11_strm1_data_valid    ( std__pe61__lane11_strm1_data_valid ),      
               .std__pe61__lane11_strm1_data_mask     ( std__pe61__lane11_strm1_data_mask  ),      

               // PE 61, Lane 12                 
               .pe61__std__lane12_strm0_ready         ( pe61__std__lane12_strm0_ready      ),      
               .std__pe61__lane12_strm0_cntl          ( std__pe61__lane12_strm0_cntl       ),      
               .std__pe61__lane12_strm0_data          ( std__pe61__lane12_strm0_data       ),      
               .std__pe61__lane12_strm0_data_valid    ( std__pe61__lane12_strm0_data_valid ),      
               .std__pe61__lane12_strm0_data_mask     ( std__pe61__lane12_strm0_data_mask  ),      

               .pe61__std__lane12_strm1_ready         ( pe61__std__lane12_strm1_ready      ),      
               .std__pe61__lane12_strm1_cntl          ( std__pe61__lane12_strm1_cntl       ),      
               .std__pe61__lane12_strm1_data          ( std__pe61__lane12_strm1_data       ),      
               .std__pe61__lane12_strm1_data_valid    ( std__pe61__lane12_strm1_data_valid ),      
               .std__pe61__lane12_strm1_data_mask     ( std__pe61__lane12_strm1_data_mask  ),      

               // PE 61, Lane 13                 
               .pe61__std__lane13_strm0_ready         ( pe61__std__lane13_strm0_ready      ),      
               .std__pe61__lane13_strm0_cntl          ( std__pe61__lane13_strm0_cntl       ),      
               .std__pe61__lane13_strm0_data          ( std__pe61__lane13_strm0_data       ),      
               .std__pe61__lane13_strm0_data_valid    ( std__pe61__lane13_strm0_data_valid ),      
               .std__pe61__lane13_strm0_data_mask     ( std__pe61__lane13_strm0_data_mask  ),      

               .pe61__std__lane13_strm1_ready         ( pe61__std__lane13_strm1_ready      ),      
               .std__pe61__lane13_strm1_cntl          ( std__pe61__lane13_strm1_cntl       ),      
               .std__pe61__lane13_strm1_data          ( std__pe61__lane13_strm1_data       ),      
               .std__pe61__lane13_strm1_data_valid    ( std__pe61__lane13_strm1_data_valid ),      
               .std__pe61__lane13_strm1_data_mask     ( std__pe61__lane13_strm1_data_mask  ),      

               // PE 61, Lane 14                 
               .pe61__std__lane14_strm0_ready         ( pe61__std__lane14_strm0_ready      ),      
               .std__pe61__lane14_strm0_cntl          ( std__pe61__lane14_strm0_cntl       ),      
               .std__pe61__lane14_strm0_data          ( std__pe61__lane14_strm0_data       ),      
               .std__pe61__lane14_strm0_data_valid    ( std__pe61__lane14_strm0_data_valid ),      
               .std__pe61__lane14_strm0_data_mask     ( std__pe61__lane14_strm0_data_mask  ),      

               .pe61__std__lane14_strm1_ready         ( pe61__std__lane14_strm1_ready      ),      
               .std__pe61__lane14_strm1_cntl          ( std__pe61__lane14_strm1_cntl       ),      
               .std__pe61__lane14_strm1_data          ( std__pe61__lane14_strm1_data       ),      
               .std__pe61__lane14_strm1_data_valid    ( std__pe61__lane14_strm1_data_valid ),      
               .std__pe61__lane14_strm1_data_mask     ( std__pe61__lane14_strm1_data_mask  ),      

               // PE 61, Lane 15                 
               .pe61__std__lane15_strm0_ready         ( pe61__std__lane15_strm0_ready      ),      
               .std__pe61__lane15_strm0_cntl          ( std__pe61__lane15_strm0_cntl       ),      
               .std__pe61__lane15_strm0_data          ( std__pe61__lane15_strm0_data       ),      
               .std__pe61__lane15_strm0_data_valid    ( std__pe61__lane15_strm0_data_valid ),      
               .std__pe61__lane15_strm0_data_mask     ( std__pe61__lane15_strm0_data_mask  ),      

               .pe61__std__lane15_strm1_ready         ( pe61__std__lane15_strm1_ready      ),      
               .std__pe61__lane15_strm1_cntl          ( std__pe61__lane15_strm1_cntl       ),      
               .std__pe61__lane15_strm1_data          ( std__pe61__lane15_strm1_data       ),      
               .std__pe61__lane15_strm1_data_valid    ( std__pe61__lane15_strm1_data_valid ),      
               .std__pe61__lane15_strm1_data_mask     ( std__pe61__lane15_strm1_data_mask  ),      

               // PE 61, Lane 16                 
               .pe61__std__lane16_strm0_ready         ( pe61__std__lane16_strm0_ready      ),      
               .std__pe61__lane16_strm0_cntl          ( std__pe61__lane16_strm0_cntl       ),      
               .std__pe61__lane16_strm0_data          ( std__pe61__lane16_strm0_data       ),      
               .std__pe61__lane16_strm0_data_valid    ( std__pe61__lane16_strm0_data_valid ),      
               .std__pe61__lane16_strm0_data_mask     ( std__pe61__lane16_strm0_data_mask  ),      

               .pe61__std__lane16_strm1_ready         ( pe61__std__lane16_strm1_ready      ),      
               .std__pe61__lane16_strm1_cntl          ( std__pe61__lane16_strm1_cntl       ),      
               .std__pe61__lane16_strm1_data          ( std__pe61__lane16_strm1_data       ),      
               .std__pe61__lane16_strm1_data_valid    ( std__pe61__lane16_strm1_data_valid ),      
               .std__pe61__lane16_strm1_data_mask     ( std__pe61__lane16_strm1_data_mask  ),      

               // PE 61, Lane 17                 
               .pe61__std__lane17_strm0_ready         ( pe61__std__lane17_strm0_ready      ),      
               .std__pe61__lane17_strm0_cntl          ( std__pe61__lane17_strm0_cntl       ),      
               .std__pe61__lane17_strm0_data          ( std__pe61__lane17_strm0_data       ),      
               .std__pe61__lane17_strm0_data_valid    ( std__pe61__lane17_strm0_data_valid ),      
               .std__pe61__lane17_strm0_data_mask     ( std__pe61__lane17_strm0_data_mask  ),      

               .pe61__std__lane17_strm1_ready         ( pe61__std__lane17_strm1_ready      ),      
               .std__pe61__lane17_strm1_cntl          ( std__pe61__lane17_strm1_cntl       ),      
               .std__pe61__lane17_strm1_data          ( std__pe61__lane17_strm1_data       ),      
               .std__pe61__lane17_strm1_data_valid    ( std__pe61__lane17_strm1_data_valid ),      
               .std__pe61__lane17_strm1_data_mask     ( std__pe61__lane17_strm1_data_mask  ),      

               // PE 61, Lane 18                 
               .pe61__std__lane18_strm0_ready         ( pe61__std__lane18_strm0_ready      ),      
               .std__pe61__lane18_strm0_cntl          ( std__pe61__lane18_strm0_cntl       ),      
               .std__pe61__lane18_strm0_data          ( std__pe61__lane18_strm0_data       ),      
               .std__pe61__lane18_strm0_data_valid    ( std__pe61__lane18_strm0_data_valid ),      
               .std__pe61__lane18_strm0_data_mask     ( std__pe61__lane18_strm0_data_mask  ),      

               .pe61__std__lane18_strm1_ready         ( pe61__std__lane18_strm1_ready      ),      
               .std__pe61__lane18_strm1_cntl          ( std__pe61__lane18_strm1_cntl       ),      
               .std__pe61__lane18_strm1_data          ( std__pe61__lane18_strm1_data       ),      
               .std__pe61__lane18_strm1_data_valid    ( std__pe61__lane18_strm1_data_valid ),      
               .std__pe61__lane18_strm1_data_mask     ( std__pe61__lane18_strm1_data_mask  ),      

               // PE 61, Lane 19                 
               .pe61__std__lane19_strm0_ready         ( pe61__std__lane19_strm0_ready      ),      
               .std__pe61__lane19_strm0_cntl          ( std__pe61__lane19_strm0_cntl       ),      
               .std__pe61__lane19_strm0_data          ( std__pe61__lane19_strm0_data       ),      
               .std__pe61__lane19_strm0_data_valid    ( std__pe61__lane19_strm0_data_valid ),      
               .std__pe61__lane19_strm0_data_mask     ( std__pe61__lane19_strm0_data_mask  ),      

               .pe61__std__lane19_strm1_ready         ( pe61__std__lane19_strm1_ready      ),      
               .std__pe61__lane19_strm1_cntl          ( std__pe61__lane19_strm1_cntl       ),      
               .std__pe61__lane19_strm1_data          ( std__pe61__lane19_strm1_data       ),      
               .std__pe61__lane19_strm1_data_valid    ( std__pe61__lane19_strm1_data_valid ),      
               .std__pe61__lane19_strm1_data_mask     ( std__pe61__lane19_strm1_data_mask  ),      

               // PE 61, Lane 20                 
               .pe61__std__lane20_strm0_ready         ( pe61__std__lane20_strm0_ready      ),      
               .std__pe61__lane20_strm0_cntl          ( std__pe61__lane20_strm0_cntl       ),      
               .std__pe61__lane20_strm0_data          ( std__pe61__lane20_strm0_data       ),      
               .std__pe61__lane20_strm0_data_valid    ( std__pe61__lane20_strm0_data_valid ),      
               .std__pe61__lane20_strm0_data_mask     ( std__pe61__lane20_strm0_data_mask  ),      

               .pe61__std__lane20_strm1_ready         ( pe61__std__lane20_strm1_ready      ),      
               .std__pe61__lane20_strm1_cntl          ( std__pe61__lane20_strm1_cntl       ),      
               .std__pe61__lane20_strm1_data          ( std__pe61__lane20_strm1_data       ),      
               .std__pe61__lane20_strm1_data_valid    ( std__pe61__lane20_strm1_data_valid ),      
               .std__pe61__lane20_strm1_data_mask     ( std__pe61__lane20_strm1_data_mask  ),      

               // PE 61, Lane 21                 
               .pe61__std__lane21_strm0_ready         ( pe61__std__lane21_strm0_ready      ),      
               .std__pe61__lane21_strm0_cntl          ( std__pe61__lane21_strm0_cntl       ),      
               .std__pe61__lane21_strm0_data          ( std__pe61__lane21_strm0_data       ),      
               .std__pe61__lane21_strm0_data_valid    ( std__pe61__lane21_strm0_data_valid ),      
               .std__pe61__lane21_strm0_data_mask     ( std__pe61__lane21_strm0_data_mask  ),      

               .pe61__std__lane21_strm1_ready         ( pe61__std__lane21_strm1_ready      ),      
               .std__pe61__lane21_strm1_cntl          ( std__pe61__lane21_strm1_cntl       ),      
               .std__pe61__lane21_strm1_data          ( std__pe61__lane21_strm1_data       ),      
               .std__pe61__lane21_strm1_data_valid    ( std__pe61__lane21_strm1_data_valid ),      
               .std__pe61__lane21_strm1_data_mask     ( std__pe61__lane21_strm1_data_mask  ),      

               // PE 61, Lane 22                 
               .pe61__std__lane22_strm0_ready         ( pe61__std__lane22_strm0_ready      ),      
               .std__pe61__lane22_strm0_cntl          ( std__pe61__lane22_strm0_cntl       ),      
               .std__pe61__lane22_strm0_data          ( std__pe61__lane22_strm0_data       ),      
               .std__pe61__lane22_strm0_data_valid    ( std__pe61__lane22_strm0_data_valid ),      
               .std__pe61__lane22_strm0_data_mask     ( std__pe61__lane22_strm0_data_mask  ),      

               .pe61__std__lane22_strm1_ready         ( pe61__std__lane22_strm1_ready      ),      
               .std__pe61__lane22_strm1_cntl          ( std__pe61__lane22_strm1_cntl       ),      
               .std__pe61__lane22_strm1_data          ( std__pe61__lane22_strm1_data       ),      
               .std__pe61__lane22_strm1_data_valid    ( std__pe61__lane22_strm1_data_valid ),      
               .std__pe61__lane22_strm1_data_mask     ( std__pe61__lane22_strm1_data_mask  ),      

               // PE 61, Lane 23                 
               .pe61__std__lane23_strm0_ready         ( pe61__std__lane23_strm0_ready      ),      
               .std__pe61__lane23_strm0_cntl          ( std__pe61__lane23_strm0_cntl       ),      
               .std__pe61__lane23_strm0_data          ( std__pe61__lane23_strm0_data       ),      
               .std__pe61__lane23_strm0_data_valid    ( std__pe61__lane23_strm0_data_valid ),      
               .std__pe61__lane23_strm0_data_mask     ( std__pe61__lane23_strm0_data_mask  ),      

               .pe61__std__lane23_strm1_ready         ( pe61__std__lane23_strm1_ready      ),      
               .std__pe61__lane23_strm1_cntl          ( std__pe61__lane23_strm1_cntl       ),      
               .std__pe61__lane23_strm1_data          ( std__pe61__lane23_strm1_data       ),      
               .std__pe61__lane23_strm1_data_valid    ( std__pe61__lane23_strm1_data_valid ),      
               .std__pe61__lane23_strm1_data_mask     ( std__pe61__lane23_strm1_data_mask  ),      

               // PE 61, Lane 24                 
               .pe61__std__lane24_strm0_ready         ( pe61__std__lane24_strm0_ready      ),      
               .std__pe61__lane24_strm0_cntl          ( std__pe61__lane24_strm0_cntl       ),      
               .std__pe61__lane24_strm0_data          ( std__pe61__lane24_strm0_data       ),      
               .std__pe61__lane24_strm0_data_valid    ( std__pe61__lane24_strm0_data_valid ),      
               .std__pe61__lane24_strm0_data_mask     ( std__pe61__lane24_strm0_data_mask  ),      

               .pe61__std__lane24_strm1_ready         ( pe61__std__lane24_strm1_ready      ),      
               .std__pe61__lane24_strm1_cntl          ( std__pe61__lane24_strm1_cntl       ),      
               .std__pe61__lane24_strm1_data          ( std__pe61__lane24_strm1_data       ),      
               .std__pe61__lane24_strm1_data_valid    ( std__pe61__lane24_strm1_data_valid ),      
               .std__pe61__lane24_strm1_data_mask     ( std__pe61__lane24_strm1_data_mask  ),      

               // PE 61, Lane 25                 
               .pe61__std__lane25_strm0_ready         ( pe61__std__lane25_strm0_ready      ),      
               .std__pe61__lane25_strm0_cntl          ( std__pe61__lane25_strm0_cntl       ),      
               .std__pe61__lane25_strm0_data          ( std__pe61__lane25_strm0_data       ),      
               .std__pe61__lane25_strm0_data_valid    ( std__pe61__lane25_strm0_data_valid ),      
               .std__pe61__lane25_strm0_data_mask     ( std__pe61__lane25_strm0_data_mask  ),      

               .pe61__std__lane25_strm1_ready         ( pe61__std__lane25_strm1_ready      ),      
               .std__pe61__lane25_strm1_cntl          ( std__pe61__lane25_strm1_cntl       ),      
               .std__pe61__lane25_strm1_data          ( std__pe61__lane25_strm1_data       ),      
               .std__pe61__lane25_strm1_data_valid    ( std__pe61__lane25_strm1_data_valid ),      
               .std__pe61__lane25_strm1_data_mask     ( std__pe61__lane25_strm1_data_mask  ),      

               // PE 61, Lane 26                 
               .pe61__std__lane26_strm0_ready         ( pe61__std__lane26_strm0_ready      ),      
               .std__pe61__lane26_strm0_cntl          ( std__pe61__lane26_strm0_cntl       ),      
               .std__pe61__lane26_strm0_data          ( std__pe61__lane26_strm0_data       ),      
               .std__pe61__lane26_strm0_data_valid    ( std__pe61__lane26_strm0_data_valid ),      
               .std__pe61__lane26_strm0_data_mask     ( std__pe61__lane26_strm0_data_mask  ),      

               .pe61__std__lane26_strm1_ready         ( pe61__std__lane26_strm1_ready      ),      
               .std__pe61__lane26_strm1_cntl          ( std__pe61__lane26_strm1_cntl       ),      
               .std__pe61__lane26_strm1_data          ( std__pe61__lane26_strm1_data       ),      
               .std__pe61__lane26_strm1_data_valid    ( std__pe61__lane26_strm1_data_valid ),      
               .std__pe61__lane26_strm1_data_mask     ( std__pe61__lane26_strm1_data_mask  ),      

               // PE 61, Lane 27                 
               .pe61__std__lane27_strm0_ready         ( pe61__std__lane27_strm0_ready      ),      
               .std__pe61__lane27_strm0_cntl          ( std__pe61__lane27_strm0_cntl       ),      
               .std__pe61__lane27_strm0_data          ( std__pe61__lane27_strm0_data       ),      
               .std__pe61__lane27_strm0_data_valid    ( std__pe61__lane27_strm0_data_valid ),      
               .std__pe61__lane27_strm0_data_mask     ( std__pe61__lane27_strm0_data_mask  ),      

               .pe61__std__lane27_strm1_ready         ( pe61__std__lane27_strm1_ready      ),      
               .std__pe61__lane27_strm1_cntl          ( std__pe61__lane27_strm1_cntl       ),      
               .std__pe61__lane27_strm1_data          ( std__pe61__lane27_strm1_data       ),      
               .std__pe61__lane27_strm1_data_valid    ( std__pe61__lane27_strm1_data_valid ),      
               .std__pe61__lane27_strm1_data_mask     ( std__pe61__lane27_strm1_data_mask  ),      

               // PE 61, Lane 28                 
               .pe61__std__lane28_strm0_ready         ( pe61__std__lane28_strm0_ready      ),      
               .std__pe61__lane28_strm0_cntl          ( std__pe61__lane28_strm0_cntl       ),      
               .std__pe61__lane28_strm0_data          ( std__pe61__lane28_strm0_data       ),      
               .std__pe61__lane28_strm0_data_valid    ( std__pe61__lane28_strm0_data_valid ),      
               .std__pe61__lane28_strm0_data_mask     ( std__pe61__lane28_strm0_data_mask  ),      

               .pe61__std__lane28_strm1_ready         ( pe61__std__lane28_strm1_ready      ),      
               .std__pe61__lane28_strm1_cntl          ( std__pe61__lane28_strm1_cntl       ),      
               .std__pe61__lane28_strm1_data          ( std__pe61__lane28_strm1_data       ),      
               .std__pe61__lane28_strm1_data_valid    ( std__pe61__lane28_strm1_data_valid ),      
               .std__pe61__lane28_strm1_data_mask     ( std__pe61__lane28_strm1_data_mask  ),      

               // PE 61, Lane 29                 
               .pe61__std__lane29_strm0_ready         ( pe61__std__lane29_strm0_ready      ),      
               .std__pe61__lane29_strm0_cntl          ( std__pe61__lane29_strm0_cntl       ),      
               .std__pe61__lane29_strm0_data          ( std__pe61__lane29_strm0_data       ),      
               .std__pe61__lane29_strm0_data_valid    ( std__pe61__lane29_strm0_data_valid ),      
               .std__pe61__lane29_strm0_data_mask     ( std__pe61__lane29_strm0_data_mask  ),      

               .pe61__std__lane29_strm1_ready         ( pe61__std__lane29_strm1_ready      ),      
               .std__pe61__lane29_strm1_cntl          ( std__pe61__lane29_strm1_cntl       ),      
               .std__pe61__lane29_strm1_data          ( std__pe61__lane29_strm1_data       ),      
               .std__pe61__lane29_strm1_data_valid    ( std__pe61__lane29_strm1_data_valid ),      
               .std__pe61__lane29_strm1_data_mask     ( std__pe61__lane29_strm1_data_mask  ),      

               // PE 61, Lane 30                 
               .pe61__std__lane30_strm0_ready         ( pe61__std__lane30_strm0_ready      ),      
               .std__pe61__lane30_strm0_cntl          ( std__pe61__lane30_strm0_cntl       ),      
               .std__pe61__lane30_strm0_data          ( std__pe61__lane30_strm0_data       ),      
               .std__pe61__lane30_strm0_data_valid    ( std__pe61__lane30_strm0_data_valid ),      
               .std__pe61__lane30_strm0_data_mask     ( std__pe61__lane30_strm0_data_mask  ),      

               .pe61__std__lane30_strm1_ready         ( pe61__std__lane30_strm1_ready      ),      
               .std__pe61__lane30_strm1_cntl          ( std__pe61__lane30_strm1_cntl       ),      
               .std__pe61__lane30_strm1_data          ( std__pe61__lane30_strm1_data       ),      
               .std__pe61__lane30_strm1_data_valid    ( std__pe61__lane30_strm1_data_valid ),      
               .std__pe61__lane30_strm1_data_mask     ( std__pe61__lane30_strm1_data_mask  ),      

               // PE 61, Lane 31                 
               .pe61__std__lane31_strm0_ready         ( pe61__std__lane31_strm0_ready      ),      
               .std__pe61__lane31_strm0_cntl          ( std__pe61__lane31_strm0_cntl       ),      
               .std__pe61__lane31_strm0_data          ( std__pe61__lane31_strm0_data       ),      
               .std__pe61__lane31_strm0_data_valid    ( std__pe61__lane31_strm0_data_valid ),      
               .std__pe61__lane31_strm0_data_mask     ( std__pe61__lane31_strm0_data_mask  ),      

               .pe61__std__lane31_strm1_ready         ( pe61__std__lane31_strm1_ready      ),      
               .std__pe61__lane31_strm1_cntl          ( std__pe61__lane31_strm1_cntl       ),      
               .std__pe61__lane31_strm1_data          ( std__pe61__lane31_strm1_data       ),      
               .std__pe61__lane31_strm1_data_valid    ( std__pe61__lane31_strm1_data_valid ),      
               .std__pe61__lane31_strm1_data_mask     ( std__pe61__lane31_strm1_data_mask  ),      

               // PE 62, Lane 0                 
               .pe62__std__lane0_strm0_ready         ( pe62__std__lane0_strm0_ready      ),      
               .std__pe62__lane0_strm0_cntl          ( std__pe62__lane0_strm0_cntl       ),      
               .std__pe62__lane0_strm0_data          ( std__pe62__lane0_strm0_data       ),      
               .std__pe62__lane0_strm0_data_valid    ( std__pe62__lane0_strm0_data_valid ),      
               .std__pe62__lane0_strm0_data_mask     ( std__pe62__lane0_strm0_data_mask  ),      

               .pe62__std__lane0_strm1_ready         ( pe62__std__lane0_strm1_ready      ),      
               .std__pe62__lane0_strm1_cntl          ( std__pe62__lane0_strm1_cntl       ),      
               .std__pe62__lane0_strm1_data          ( std__pe62__lane0_strm1_data       ),      
               .std__pe62__lane0_strm1_data_valid    ( std__pe62__lane0_strm1_data_valid ),      
               .std__pe62__lane0_strm1_data_mask     ( std__pe62__lane0_strm1_data_mask  ),      

               // PE 62, Lane 1                 
               .pe62__std__lane1_strm0_ready         ( pe62__std__lane1_strm0_ready      ),      
               .std__pe62__lane1_strm0_cntl          ( std__pe62__lane1_strm0_cntl       ),      
               .std__pe62__lane1_strm0_data          ( std__pe62__lane1_strm0_data       ),      
               .std__pe62__lane1_strm0_data_valid    ( std__pe62__lane1_strm0_data_valid ),      
               .std__pe62__lane1_strm0_data_mask     ( std__pe62__lane1_strm0_data_mask  ),      

               .pe62__std__lane1_strm1_ready         ( pe62__std__lane1_strm1_ready      ),      
               .std__pe62__lane1_strm1_cntl          ( std__pe62__lane1_strm1_cntl       ),      
               .std__pe62__lane1_strm1_data          ( std__pe62__lane1_strm1_data       ),      
               .std__pe62__lane1_strm1_data_valid    ( std__pe62__lane1_strm1_data_valid ),      
               .std__pe62__lane1_strm1_data_mask     ( std__pe62__lane1_strm1_data_mask  ),      

               // PE 62, Lane 2                 
               .pe62__std__lane2_strm0_ready         ( pe62__std__lane2_strm0_ready      ),      
               .std__pe62__lane2_strm0_cntl          ( std__pe62__lane2_strm0_cntl       ),      
               .std__pe62__lane2_strm0_data          ( std__pe62__lane2_strm0_data       ),      
               .std__pe62__lane2_strm0_data_valid    ( std__pe62__lane2_strm0_data_valid ),      
               .std__pe62__lane2_strm0_data_mask     ( std__pe62__lane2_strm0_data_mask  ),      

               .pe62__std__lane2_strm1_ready         ( pe62__std__lane2_strm1_ready      ),      
               .std__pe62__lane2_strm1_cntl          ( std__pe62__lane2_strm1_cntl       ),      
               .std__pe62__lane2_strm1_data          ( std__pe62__lane2_strm1_data       ),      
               .std__pe62__lane2_strm1_data_valid    ( std__pe62__lane2_strm1_data_valid ),      
               .std__pe62__lane2_strm1_data_mask     ( std__pe62__lane2_strm1_data_mask  ),      

               // PE 62, Lane 3                 
               .pe62__std__lane3_strm0_ready         ( pe62__std__lane3_strm0_ready      ),      
               .std__pe62__lane3_strm0_cntl          ( std__pe62__lane3_strm0_cntl       ),      
               .std__pe62__lane3_strm0_data          ( std__pe62__lane3_strm0_data       ),      
               .std__pe62__lane3_strm0_data_valid    ( std__pe62__lane3_strm0_data_valid ),      
               .std__pe62__lane3_strm0_data_mask     ( std__pe62__lane3_strm0_data_mask  ),      

               .pe62__std__lane3_strm1_ready         ( pe62__std__lane3_strm1_ready      ),      
               .std__pe62__lane3_strm1_cntl          ( std__pe62__lane3_strm1_cntl       ),      
               .std__pe62__lane3_strm1_data          ( std__pe62__lane3_strm1_data       ),      
               .std__pe62__lane3_strm1_data_valid    ( std__pe62__lane3_strm1_data_valid ),      
               .std__pe62__lane3_strm1_data_mask     ( std__pe62__lane3_strm1_data_mask  ),      

               // PE 62, Lane 4                 
               .pe62__std__lane4_strm0_ready         ( pe62__std__lane4_strm0_ready      ),      
               .std__pe62__lane4_strm0_cntl          ( std__pe62__lane4_strm0_cntl       ),      
               .std__pe62__lane4_strm0_data          ( std__pe62__lane4_strm0_data       ),      
               .std__pe62__lane4_strm0_data_valid    ( std__pe62__lane4_strm0_data_valid ),      
               .std__pe62__lane4_strm0_data_mask     ( std__pe62__lane4_strm0_data_mask  ),      

               .pe62__std__lane4_strm1_ready         ( pe62__std__lane4_strm1_ready      ),      
               .std__pe62__lane4_strm1_cntl          ( std__pe62__lane4_strm1_cntl       ),      
               .std__pe62__lane4_strm1_data          ( std__pe62__lane4_strm1_data       ),      
               .std__pe62__lane4_strm1_data_valid    ( std__pe62__lane4_strm1_data_valid ),      
               .std__pe62__lane4_strm1_data_mask     ( std__pe62__lane4_strm1_data_mask  ),      

               // PE 62, Lane 5                 
               .pe62__std__lane5_strm0_ready         ( pe62__std__lane5_strm0_ready      ),      
               .std__pe62__lane5_strm0_cntl          ( std__pe62__lane5_strm0_cntl       ),      
               .std__pe62__lane5_strm0_data          ( std__pe62__lane5_strm0_data       ),      
               .std__pe62__lane5_strm0_data_valid    ( std__pe62__lane5_strm0_data_valid ),      
               .std__pe62__lane5_strm0_data_mask     ( std__pe62__lane5_strm0_data_mask  ),      

               .pe62__std__lane5_strm1_ready         ( pe62__std__lane5_strm1_ready      ),      
               .std__pe62__lane5_strm1_cntl          ( std__pe62__lane5_strm1_cntl       ),      
               .std__pe62__lane5_strm1_data          ( std__pe62__lane5_strm1_data       ),      
               .std__pe62__lane5_strm1_data_valid    ( std__pe62__lane5_strm1_data_valid ),      
               .std__pe62__lane5_strm1_data_mask     ( std__pe62__lane5_strm1_data_mask  ),      

               // PE 62, Lane 6                 
               .pe62__std__lane6_strm0_ready         ( pe62__std__lane6_strm0_ready      ),      
               .std__pe62__lane6_strm0_cntl          ( std__pe62__lane6_strm0_cntl       ),      
               .std__pe62__lane6_strm0_data          ( std__pe62__lane6_strm0_data       ),      
               .std__pe62__lane6_strm0_data_valid    ( std__pe62__lane6_strm0_data_valid ),      
               .std__pe62__lane6_strm0_data_mask     ( std__pe62__lane6_strm0_data_mask  ),      

               .pe62__std__lane6_strm1_ready         ( pe62__std__lane6_strm1_ready      ),      
               .std__pe62__lane6_strm1_cntl          ( std__pe62__lane6_strm1_cntl       ),      
               .std__pe62__lane6_strm1_data          ( std__pe62__lane6_strm1_data       ),      
               .std__pe62__lane6_strm1_data_valid    ( std__pe62__lane6_strm1_data_valid ),      
               .std__pe62__lane6_strm1_data_mask     ( std__pe62__lane6_strm1_data_mask  ),      

               // PE 62, Lane 7                 
               .pe62__std__lane7_strm0_ready         ( pe62__std__lane7_strm0_ready      ),      
               .std__pe62__lane7_strm0_cntl          ( std__pe62__lane7_strm0_cntl       ),      
               .std__pe62__lane7_strm0_data          ( std__pe62__lane7_strm0_data       ),      
               .std__pe62__lane7_strm0_data_valid    ( std__pe62__lane7_strm0_data_valid ),      
               .std__pe62__lane7_strm0_data_mask     ( std__pe62__lane7_strm0_data_mask  ),      

               .pe62__std__lane7_strm1_ready         ( pe62__std__lane7_strm1_ready      ),      
               .std__pe62__lane7_strm1_cntl          ( std__pe62__lane7_strm1_cntl       ),      
               .std__pe62__lane7_strm1_data          ( std__pe62__lane7_strm1_data       ),      
               .std__pe62__lane7_strm1_data_valid    ( std__pe62__lane7_strm1_data_valid ),      
               .std__pe62__lane7_strm1_data_mask     ( std__pe62__lane7_strm1_data_mask  ),      

               // PE 62, Lane 8                 
               .pe62__std__lane8_strm0_ready         ( pe62__std__lane8_strm0_ready      ),      
               .std__pe62__lane8_strm0_cntl          ( std__pe62__lane8_strm0_cntl       ),      
               .std__pe62__lane8_strm0_data          ( std__pe62__lane8_strm0_data       ),      
               .std__pe62__lane8_strm0_data_valid    ( std__pe62__lane8_strm0_data_valid ),      
               .std__pe62__lane8_strm0_data_mask     ( std__pe62__lane8_strm0_data_mask  ),      

               .pe62__std__lane8_strm1_ready         ( pe62__std__lane8_strm1_ready      ),      
               .std__pe62__lane8_strm1_cntl          ( std__pe62__lane8_strm1_cntl       ),      
               .std__pe62__lane8_strm1_data          ( std__pe62__lane8_strm1_data       ),      
               .std__pe62__lane8_strm1_data_valid    ( std__pe62__lane8_strm1_data_valid ),      
               .std__pe62__lane8_strm1_data_mask     ( std__pe62__lane8_strm1_data_mask  ),      

               // PE 62, Lane 9                 
               .pe62__std__lane9_strm0_ready         ( pe62__std__lane9_strm0_ready      ),      
               .std__pe62__lane9_strm0_cntl          ( std__pe62__lane9_strm0_cntl       ),      
               .std__pe62__lane9_strm0_data          ( std__pe62__lane9_strm0_data       ),      
               .std__pe62__lane9_strm0_data_valid    ( std__pe62__lane9_strm0_data_valid ),      
               .std__pe62__lane9_strm0_data_mask     ( std__pe62__lane9_strm0_data_mask  ),      

               .pe62__std__lane9_strm1_ready         ( pe62__std__lane9_strm1_ready      ),      
               .std__pe62__lane9_strm1_cntl          ( std__pe62__lane9_strm1_cntl       ),      
               .std__pe62__lane9_strm1_data          ( std__pe62__lane9_strm1_data       ),      
               .std__pe62__lane9_strm1_data_valid    ( std__pe62__lane9_strm1_data_valid ),      
               .std__pe62__lane9_strm1_data_mask     ( std__pe62__lane9_strm1_data_mask  ),      

               // PE 62, Lane 10                 
               .pe62__std__lane10_strm0_ready         ( pe62__std__lane10_strm0_ready      ),      
               .std__pe62__lane10_strm0_cntl          ( std__pe62__lane10_strm0_cntl       ),      
               .std__pe62__lane10_strm0_data          ( std__pe62__lane10_strm0_data       ),      
               .std__pe62__lane10_strm0_data_valid    ( std__pe62__lane10_strm0_data_valid ),      
               .std__pe62__lane10_strm0_data_mask     ( std__pe62__lane10_strm0_data_mask  ),      

               .pe62__std__lane10_strm1_ready         ( pe62__std__lane10_strm1_ready      ),      
               .std__pe62__lane10_strm1_cntl          ( std__pe62__lane10_strm1_cntl       ),      
               .std__pe62__lane10_strm1_data          ( std__pe62__lane10_strm1_data       ),      
               .std__pe62__lane10_strm1_data_valid    ( std__pe62__lane10_strm1_data_valid ),      
               .std__pe62__lane10_strm1_data_mask     ( std__pe62__lane10_strm1_data_mask  ),      

               // PE 62, Lane 11                 
               .pe62__std__lane11_strm0_ready         ( pe62__std__lane11_strm0_ready      ),      
               .std__pe62__lane11_strm0_cntl          ( std__pe62__lane11_strm0_cntl       ),      
               .std__pe62__lane11_strm0_data          ( std__pe62__lane11_strm0_data       ),      
               .std__pe62__lane11_strm0_data_valid    ( std__pe62__lane11_strm0_data_valid ),      
               .std__pe62__lane11_strm0_data_mask     ( std__pe62__lane11_strm0_data_mask  ),      

               .pe62__std__lane11_strm1_ready         ( pe62__std__lane11_strm1_ready      ),      
               .std__pe62__lane11_strm1_cntl          ( std__pe62__lane11_strm1_cntl       ),      
               .std__pe62__lane11_strm1_data          ( std__pe62__lane11_strm1_data       ),      
               .std__pe62__lane11_strm1_data_valid    ( std__pe62__lane11_strm1_data_valid ),      
               .std__pe62__lane11_strm1_data_mask     ( std__pe62__lane11_strm1_data_mask  ),      

               // PE 62, Lane 12                 
               .pe62__std__lane12_strm0_ready         ( pe62__std__lane12_strm0_ready      ),      
               .std__pe62__lane12_strm0_cntl          ( std__pe62__lane12_strm0_cntl       ),      
               .std__pe62__lane12_strm0_data          ( std__pe62__lane12_strm0_data       ),      
               .std__pe62__lane12_strm0_data_valid    ( std__pe62__lane12_strm0_data_valid ),      
               .std__pe62__lane12_strm0_data_mask     ( std__pe62__lane12_strm0_data_mask  ),      

               .pe62__std__lane12_strm1_ready         ( pe62__std__lane12_strm1_ready      ),      
               .std__pe62__lane12_strm1_cntl          ( std__pe62__lane12_strm1_cntl       ),      
               .std__pe62__lane12_strm1_data          ( std__pe62__lane12_strm1_data       ),      
               .std__pe62__lane12_strm1_data_valid    ( std__pe62__lane12_strm1_data_valid ),      
               .std__pe62__lane12_strm1_data_mask     ( std__pe62__lane12_strm1_data_mask  ),      

               // PE 62, Lane 13                 
               .pe62__std__lane13_strm0_ready         ( pe62__std__lane13_strm0_ready      ),      
               .std__pe62__lane13_strm0_cntl          ( std__pe62__lane13_strm0_cntl       ),      
               .std__pe62__lane13_strm0_data          ( std__pe62__lane13_strm0_data       ),      
               .std__pe62__lane13_strm0_data_valid    ( std__pe62__lane13_strm0_data_valid ),      
               .std__pe62__lane13_strm0_data_mask     ( std__pe62__lane13_strm0_data_mask  ),      

               .pe62__std__lane13_strm1_ready         ( pe62__std__lane13_strm1_ready      ),      
               .std__pe62__lane13_strm1_cntl          ( std__pe62__lane13_strm1_cntl       ),      
               .std__pe62__lane13_strm1_data          ( std__pe62__lane13_strm1_data       ),      
               .std__pe62__lane13_strm1_data_valid    ( std__pe62__lane13_strm1_data_valid ),      
               .std__pe62__lane13_strm1_data_mask     ( std__pe62__lane13_strm1_data_mask  ),      

               // PE 62, Lane 14                 
               .pe62__std__lane14_strm0_ready         ( pe62__std__lane14_strm0_ready      ),      
               .std__pe62__lane14_strm0_cntl          ( std__pe62__lane14_strm0_cntl       ),      
               .std__pe62__lane14_strm0_data          ( std__pe62__lane14_strm0_data       ),      
               .std__pe62__lane14_strm0_data_valid    ( std__pe62__lane14_strm0_data_valid ),      
               .std__pe62__lane14_strm0_data_mask     ( std__pe62__lane14_strm0_data_mask  ),      

               .pe62__std__lane14_strm1_ready         ( pe62__std__lane14_strm1_ready      ),      
               .std__pe62__lane14_strm1_cntl          ( std__pe62__lane14_strm1_cntl       ),      
               .std__pe62__lane14_strm1_data          ( std__pe62__lane14_strm1_data       ),      
               .std__pe62__lane14_strm1_data_valid    ( std__pe62__lane14_strm1_data_valid ),      
               .std__pe62__lane14_strm1_data_mask     ( std__pe62__lane14_strm1_data_mask  ),      

               // PE 62, Lane 15                 
               .pe62__std__lane15_strm0_ready         ( pe62__std__lane15_strm0_ready      ),      
               .std__pe62__lane15_strm0_cntl          ( std__pe62__lane15_strm0_cntl       ),      
               .std__pe62__lane15_strm0_data          ( std__pe62__lane15_strm0_data       ),      
               .std__pe62__lane15_strm0_data_valid    ( std__pe62__lane15_strm0_data_valid ),      
               .std__pe62__lane15_strm0_data_mask     ( std__pe62__lane15_strm0_data_mask  ),      

               .pe62__std__lane15_strm1_ready         ( pe62__std__lane15_strm1_ready      ),      
               .std__pe62__lane15_strm1_cntl          ( std__pe62__lane15_strm1_cntl       ),      
               .std__pe62__lane15_strm1_data          ( std__pe62__lane15_strm1_data       ),      
               .std__pe62__lane15_strm1_data_valid    ( std__pe62__lane15_strm1_data_valid ),      
               .std__pe62__lane15_strm1_data_mask     ( std__pe62__lane15_strm1_data_mask  ),      

               // PE 62, Lane 16                 
               .pe62__std__lane16_strm0_ready         ( pe62__std__lane16_strm0_ready      ),      
               .std__pe62__lane16_strm0_cntl          ( std__pe62__lane16_strm0_cntl       ),      
               .std__pe62__lane16_strm0_data          ( std__pe62__lane16_strm0_data       ),      
               .std__pe62__lane16_strm0_data_valid    ( std__pe62__lane16_strm0_data_valid ),      
               .std__pe62__lane16_strm0_data_mask     ( std__pe62__lane16_strm0_data_mask  ),      

               .pe62__std__lane16_strm1_ready         ( pe62__std__lane16_strm1_ready      ),      
               .std__pe62__lane16_strm1_cntl          ( std__pe62__lane16_strm1_cntl       ),      
               .std__pe62__lane16_strm1_data          ( std__pe62__lane16_strm1_data       ),      
               .std__pe62__lane16_strm1_data_valid    ( std__pe62__lane16_strm1_data_valid ),      
               .std__pe62__lane16_strm1_data_mask     ( std__pe62__lane16_strm1_data_mask  ),      

               // PE 62, Lane 17                 
               .pe62__std__lane17_strm0_ready         ( pe62__std__lane17_strm0_ready      ),      
               .std__pe62__lane17_strm0_cntl          ( std__pe62__lane17_strm0_cntl       ),      
               .std__pe62__lane17_strm0_data          ( std__pe62__lane17_strm0_data       ),      
               .std__pe62__lane17_strm0_data_valid    ( std__pe62__lane17_strm0_data_valid ),      
               .std__pe62__lane17_strm0_data_mask     ( std__pe62__lane17_strm0_data_mask  ),      

               .pe62__std__lane17_strm1_ready         ( pe62__std__lane17_strm1_ready      ),      
               .std__pe62__lane17_strm1_cntl          ( std__pe62__lane17_strm1_cntl       ),      
               .std__pe62__lane17_strm1_data          ( std__pe62__lane17_strm1_data       ),      
               .std__pe62__lane17_strm1_data_valid    ( std__pe62__lane17_strm1_data_valid ),      
               .std__pe62__lane17_strm1_data_mask     ( std__pe62__lane17_strm1_data_mask  ),      

               // PE 62, Lane 18                 
               .pe62__std__lane18_strm0_ready         ( pe62__std__lane18_strm0_ready      ),      
               .std__pe62__lane18_strm0_cntl          ( std__pe62__lane18_strm0_cntl       ),      
               .std__pe62__lane18_strm0_data          ( std__pe62__lane18_strm0_data       ),      
               .std__pe62__lane18_strm0_data_valid    ( std__pe62__lane18_strm0_data_valid ),      
               .std__pe62__lane18_strm0_data_mask     ( std__pe62__lane18_strm0_data_mask  ),      

               .pe62__std__lane18_strm1_ready         ( pe62__std__lane18_strm1_ready      ),      
               .std__pe62__lane18_strm1_cntl          ( std__pe62__lane18_strm1_cntl       ),      
               .std__pe62__lane18_strm1_data          ( std__pe62__lane18_strm1_data       ),      
               .std__pe62__lane18_strm1_data_valid    ( std__pe62__lane18_strm1_data_valid ),      
               .std__pe62__lane18_strm1_data_mask     ( std__pe62__lane18_strm1_data_mask  ),      

               // PE 62, Lane 19                 
               .pe62__std__lane19_strm0_ready         ( pe62__std__lane19_strm0_ready      ),      
               .std__pe62__lane19_strm0_cntl          ( std__pe62__lane19_strm0_cntl       ),      
               .std__pe62__lane19_strm0_data          ( std__pe62__lane19_strm0_data       ),      
               .std__pe62__lane19_strm0_data_valid    ( std__pe62__lane19_strm0_data_valid ),      
               .std__pe62__lane19_strm0_data_mask     ( std__pe62__lane19_strm0_data_mask  ),      

               .pe62__std__lane19_strm1_ready         ( pe62__std__lane19_strm1_ready      ),      
               .std__pe62__lane19_strm1_cntl          ( std__pe62__lane19_strm1_cntl       ),      
               .std__pe62__lane19_strm1_data          ( std__pe62__lane19_strm1_data       ),      
               .std__pe62__lane19_strm1_data_valid    ( std__pe62__lane19_strm1_data_valid ),      
               .std__pe62__lane19_strm1_data_mask     ( std__pe62__lane19_strm1_data_mask  ),      

               // PE 62, Lane 20                 
               .pe62__std__lane20_strm0_ready         ( pe62__std__lane20_strm0_ready      ),      
               .std__pe62__lane20_strm0_cntl          ( std__pe62__lane20_strm0_cntl       ),      
               .std__pe62__lane20_strm0_data          ( std__pe62__lane20_strm0_data       ),      
               .std__pe62__lane20_strm0_data_valid    ( std__pe62__lane20_strm0_data_valid ),      
               .std__pe62__lane20_strm0_data_mask     ( std__pe62__lane20_strm0_data_mask  ),      

               .pe62__std__lane20_strm1_ready         ( pe62__std__lane20_strm1_ready      ),      
               .std__pe62__lane20_strm1_cntl          ( std__pe62__lane20_strm1_cntl       ),      
               .std__pe62__lane20_strm1_data          ( std__pe62__lane20_strm1_data       ),      
               .std__pe62__lane20_strm1_data_valid    ( std__pe62__lane20_strm1_data_valid ),      
               .std__pe62__lane20_strm1_data_mask     ( std__pe62__lane20_strm1_data_mask  ),      

               // PE 62, Lane 21                 
               .pe62__std__lane21_strm0_ready         ( pe62__std__lane21_strm0_ready      ),      
               .std__pe62__lane21_strm0_cntl          ( std__pe62__lane21_strm0_cntl       ),      
               .std__pe62__lane21_strm0_data          ( std__pe62__lane21_strm0_data       ),      
               .std__pe62__lane21_strm0_data_valid    ( std__pe62__lane21_strm0_data_valid ),      
               .std__pe62__lane21_strm0_data_mask     ( std__pe62__lane21_strm0_data_mask  ),      

               .pe62__std__lane21_strm1_ready         ( pe62__std__lane21_strm1_ready      ),      
               .std__pe62__lane21_strm1_cntl          ( std__pe62__lane21_strm1_cntl       ),      
               .std__pe62__lane21_strm1_data          ( std__pe62__lane21_strm1_data       ),      
               .std__pe62__lane21_strm1_data_valid    ( std__pe62__lane21_strm1_data_valid ),      
               .std__pe62__lane21_strm1_data_mask     ( std__pe62__lane21_strm1_data_mask  ),      

               // PE 62, Lane 22                 
               .pe62__std__lane22_strm0_ready         ( pe62__std__lane22_strm0_ready      ),      
               .std__pe62__lane22_strm0_cntl          ( std__pe62__lane22_strm0_cntl       ),      
               .std__pe62__lane22_strm0_data          ( std__pe62__lane22_strm0_data       ),      
               .std__pe62__lane22_strm0_data_valid    ( std__pe62__lane22_strm0_data_valid ),      
               .std__pe62__lane22_strm0_data_mask     ( std__pe62__lane22_strm0_data_mask  ),      

               .pe62__std__lane22_strm1_ready         ( pe62__std__lane22_strm1_ready      ),      
               .std__pe62__lane22_strm1_cntl          ( std__pe62__lane22_strm1_cntl       ),      
               .std__pe62__lane22_strm1_data          ( std__pe62__lane22_strm1_data       ),      
               .std__pe62__lane22_strm1_data_valid    ( std__pe62__lane22_strm1_data_valid ),      
               .std__pe62__lane22_strm1_data_mask     ( std__pe62__lane22_strm1_data_mask  ),      

               // PE 62, Lane 23                 
               .pe62__std__lane23_strm0_ready         ( pe62__std__lane23_strm0_ready      ),      
               .std__pe62__lane23_strm0_cntl          ( std__pe62__lane23_strm0_cntl       ),      
               .std__pe62__lane23_strm0_data          ( std__pe62__lane23_strm0_data       ),      
               .std__pe62__lane23_strm0_data_valid    ( std__pe62__lane23_strm0_data_valid ),      
               .std__pe62__lane23_strm0_data_mask     ( std__pe62__lane23_strm0_data_mask  ),      

               .pe62__std__lane23_strm1_ready         ( pe62__std__lane23_strm1_ready      ),      
               .std__pe62__lane23_strm1_cntl          ( std__pe62__lane23_strm1_cntl       ),      
               .std__pe62__lane23_strm1_data          ( std__pe62__lane23_strm1_data       ),      
               .std__pe62__lane23_strm1_data_valid    ( std__pe62__lane23_strm1_data_valid ),      
               .std__pe62__lane23_strm1_data_mask     ( std__pe62__lane23_strm1_data_mask  ),      

               // PE 62, Lane 24                 
               .pe62__std__lane24_strm0_ready         ( pe62__std__lane24_strm0_ready      ),      
               .std__pe62__lane24_strm0_cntl          ( std__pe62__lane24_strm0_cntl       ),      
               .std__pe62__lane24_strm0_data          ( std__pe62__lane24_strm0_data       ),      
               .std__pe62__lane24_strm0_data_valid    ( std__pe62__lane24_strm0_data_valid ),      
               .std__pe62__lane24_strm0_data_mask     ( std__pe62__lane24_strm0_data_mask  ),      

               .pe62__std__lane24_strm1_ready         ( pe62__std__lane24_strm1_ready      ),      
               .std__pe62__lane24_strm1_cntl          ( std__pe62__lane24_strm1_cntl       ),      
               .std__pe62__lane24_strm1_data          ( std__pe62__lane24_strm1_data       ),      
               .std__pe62__lane24_strm1_data_valid    ( std__pe62__lane24_strm1_data_valid ),      
               .std__pe62__lane24_strm1_data_mask     ( std__pe62__lane24_strm1_data_mask  ),      

               // PE 62, Lane 25                 
               .pe62__std__lane25_strm0_ready         ( pe62__std__lane25_strm0_ready      ),      
               .std__pe62__lane25_strm0_cntl          ( std__pe62__lane25_strm0_cntl       ),      
               .std__pe62__lane25_strm0_data          ( std__pe62__lane25_strm0_data       ),      
               .std__pe62__lane25_strm0_data_valid    ( std__pe62__lane25_strm0_data_valid ),      
               .std__pe62__lane25_strm0_data_mask     ( std__pe62__lane25_strm0_data_mask  ),      

               .pe62__std__lane25_strm1_ready         ( pe62__std__lane25_strm1_ready      ),      
               .std__pe62__lane25_strm1_cntl          ( std__pe62__lane25_strm1_cntl       ),      
               .std__pe62__lane25_strm1_data          ( std__pe62__lane25_strm1_data       ),      
               .std__pe62__lane25_strm1_data_valid    ( std__pe62__lane25_strm1_data_valid ),      
               .std__pe62__lane25_strm1_data_mask     ( std__pe62__lane25_strm1_data_mask  ),      

               // PE 62, Lane 26                 
               .pe62__std__lane26_strm0_ready         ( pe62__std__lane26_strm0_ready      ),      
               .std__pe62__lane26_strm0_cntl          ( std__pe62__lane26_strm0_cntl       ),      
               .std__pe62__lane26_strm0_data          ( std__pe62__lane26_strm0_data       ),      
               .std__pe62__lane26_strm0_data_valid    ( std__pe62__lane26_strm0_data_valid ),      
               .std__pe62__lane26_strm0_data_mask     ( std__pe62__lane26_strm0_data_mask  ),      

               .pe62__std__lane26_strm1_ready         ( pe62__std__lane26_strm1_ready      ),      
               .std__pe62__lane26_strm1_cntl          ( std__pe62__lane26_strm1_cntl       ),      
               .std__pe62__lane26_strm1_data          ( std__pe62__lane26_strm1_data       ),      
               .std__pe62__lane26_strm1_data_valid    ( std__pe62__lane26_strm1_data_valid ),      
               .std__pe62__lane26_strm1_data_mask     ( std__pe62__lane26_strm1_data_mask  ),      

               // PE 62, Lane 27                 
               .pe62__std__lane27_strm0_ready         ( pe62__std__lane27_strm0_ready      ),      
               .std__pe62__lane27_strm0_cntl          ( std__pe62__lane27_strm0_cntl       ),      
               .std__pe62__lane27_strm0_data          ( std__pe62__lane27_strm0_data       ),      
               .std__pe62__lane27_strm0_data_valid    ( std__pe62__lane27_strm0_data_valid ),      
               .std__pe62__lane27_strm0_data_mask     ( std__pe62__lane27_strm0_data_mask  ),      

               .pe62__std__lane27_strm1_ready         ( pe62__std__lane27_strm1_ready      ),      
               .std__pe62__lane27_strm1_cntl          ( std__pe62__lane27_strm1_cntl       ),      
               .std__pe62__lane27_strm1_data          ( std__pe62__lane27_strm1_data       ),      
               .std__pe62__lane27_strm1_data_valid    ( std__pe62__lane27_strm1_data_valid ),      
               .std__pe62__lane27_strm1_data_mask     ( std__pe62__lane27_strm1_data_mask  ),      

               // PE 62, Lane 28                 
               .pe62__std__lane28_strm0_ready         ( pe62__std__lane28_strm0_ready      ),      
               .std__pe62__lane28_strm0_cntl          ( std__pe62__lane28_strm0_cntl       ),      
               .std__pe62__lane28_strm0_data          ( std__pe62__lane28_strm0_data       ),      
               .std__pe62__lane28_strm0_data_valid    ( std__pe62__lane28_strm0_data_valid ),      
               .std__pe62__lane28_strm0_data_mask     ( std__pe62__lane28_strm0_data_mask  ),      

               .pe62__std__lane28_strm1_ready         ( pe62__std__lane28_strm1_ready      ),      
               .std__pe62__lane28_strm1_cntl          ( std__pe62__lane28_strm1_cntl       ),      
               .std__pe62__lane28_strm1_data          ( std__pe62__lane28_strm1_data       ),      
               .std__pe62__lane28_strm1_data_valid    ( std__pe62__lane28_strm1_data_valid ),      
               .std__pe62__lane28_strm1_data_mask     ( std__pe62__lane28_strm1_data_mask  ),      

               // PE 62, Lane 29                 
               .pe62__std__lane29_strm0_ready         ( pe62__std__lane29_strm0_ready      ),      
               .std__pe62__lane29_strm0_cntl          ( std__pe62__lane29_strm0_cntl       ),      
               .std__pe62__lane29_strm0_data          ( std__pe62__lane29_strm0_data       ),      
               .std__pe62__lane29_strm0_data_valid    ( std__pe62__lane29_strm0_data_valid ),      
               .std__pe62__lane29_strm0_data_mask     ( std__pe62__lane29_strm0_data_mask  ),      

               .pe62__std__lane29_strm1_ready         ( pe62__std__lane29_strm1_ready      ),      
               .std__pe62__lane29_strm1_cntl          ( std__pe62__lane29_strm1_cntl       ),      
               .std__pe62__lane29_strm1_data          ( std__pe62__lane29_strm1_data       ),      
               .std__pe62__lane29_strm1_data_valid    ( std__pe62__lane29_strm1_data_valid ),      
               .std__pe62__lane29_strm1_data_mask     ( std__pe62__lane29_strm1_data_mask  ),      

               // PE 62, Lane 30                 
               .pe62__std__lane30_strm0_ready         ( pe62__std__lane30_strm0_ready      ),      
               .std__pe62__lane30_strm0_cntl          ( std__pe62__lane30_strm0_cntl       ),      
               .std__pe62__lane30_strm0_data          ( std__pe62__lane30_strm0_data       ),      
               .std__pe62__lane30_strm0_data_valid    ( std__pe62__lane30_strm0_data_valid ),      
               .std__pe62__lane30_strm0_data_mask     ( std__pe62__lane30_strm0_data_mask  ),      

               .pe62__std__lane30_strm1_ready         ( pe62__std__lane30_strm1_ready      ),      
               .std__pe62__lane30_strm1_cntl          ( std__pe62__lane30_strm1_cntl       ),      
               .std__pe62__lane30_strm1_data          ( std__pe62__lane30_strm1_data       ),      
               .std__pe62__lane30_strm1_data_valid    ( std__pe62__lane30_strm1_data_valid ),      
               .std__pe62__lane30_strm1_data_mask     ( std__pe62__lane30_strm1_data_mask  ),      

               // PE 62, Lane 31                 
               .pe62__std__lane31_strm0_ready         ( pe62__std__lane31_strm0_ready      ),      
               .std__pe62__lane31_strm0_cntl          ( std__pe62__lane31_strm0_cntl       ),      
               .std__pe62__lane31_strm0_data          ( std__pe62__lane31_strm0_data       ),      
               .std__pe62__lane31_strm0_data_valid    ( std__pe62__lane31_strm0_data_valid ),      
               .std__pe62__lane31_strm0_data_mask     ( std__pe62__lane31_strm0_data_mask  ),      

               .pe62__std__lane31_strm1_ready         ( pe62__std__lane31_strm1_ready      ),      
               .std__pe62__lane31_strm1_cntl          ( std__pe62__lane31_strm1_cntl       ),      
               .std__pe62__lane31_strm1_data          ( std__pe62__lane31_strm1_data       ),      
               .std__pe62__lane31_strm1_data_valid    ( std__pe62__lane31_strm1_data_valid ),      
               .std__pe62__lane31_strm1_data_mask     ( std__pe62__lane31_strm1_data_mask  ),      

               // PE 63, Lane 0                 
               .pe63__std__lane0_strm0_ready         ( pe63__std__lane0_strm0_ready      ),      
               .std__pe63__lane0_strm0_cntl          ( std__pe63__lane0_strm0_cntl       ),      
               .std__pe63__lane0_strm0_data          ( std__pe63__lane0_strm0_data       ),      
               .std__pe63__lane0_strm0_data_valid    ( std__pe63__lane0_strm0_data_valid ),      
               .std__pe63__lane0_strm0_data_mask     ( std__pe63__lane0_strm0_data_mask  ),      

               .pe63__std__lane0_strm1_ready         ( pe63__std__lane0_strm1_ready      ),      
               .std__pe63__lane0_strm1_cntl          ( std__pe63__lane0_strm1_cntl       ),      
               .std__pe63__lane0_strm1_data          ( std__pe63__lane0_strm1_data       ),      
               .std__pe63__lane0_strm1_data_valid    ( std__pe63__lane0_strm1_data_valid ),      
               .std__pe63__lane0_strm1_data_mask     ( std__pe63__lane0_strm1_data_mask  ),      

               // PE 63, Lane 1                 
               .pe63__std__lane1_strm0_ready         ( pe63__std__lane1_strm0_ready      ),      
               .std__pe63__lane1_strm0_cntl          ( std__pe63__lane1_strm0_cntl       ),      
               .std__pe63__lane1_strm0_data          ( std__pe63__lane1_strm0_data       ),      
               .std__pe63__lane1_strm0_data_valid    ( std__pe63__lane1_strm0_data_valid ),      
               .std__pe63__lane1_strm0_data_mask     ( std__pe63__lane1_strm0_data_mask  ),      

               .pe63__std__lane1_strm1_ready         ( pe63__std__lane1_strm1_ready      ),      
               .std__pe63__lane1_strm1_cntl          ( std__pe63__lane1_strm1_cntl       ),      
               .std__pe63__lane1_strm1_data          ( std__pe63__lane1_strm1_data       ),      
               .std__pe63__lane1_strm1_data_valid    ( std__pe63__lane1_strm1_data_valid ),      
               .std__pe63__lane1_strm1_data_mask     ( std__pe63__lane1_strm1_data_mask  ),      

               // PE 63, Lane 2                 
               .pe63__std__lane2_strm0_ready         ( pe63__std__lane2_strm0_ready      ),      
               .std__pe63__lane2_strm0_cntl          ( std__pe63__lane2_strm0_cntl       ),      
               .std__pe63__lane2_strm0_data          ( std__pe63__lane2_strm0_data       ),      
               .std__pe63__lane2_strm0_data_valid    ( std__pe63__lane2_strm0_data_valid ),      
               .std__pe63__lane2_strm0_data_mask     ( std__pe63__lane2_strm0_data_mask  ),      

               .pe63__std__lane2_strm1_ready         ( pe63__std__lane2_strm1_ready      ),      
               .std__pe63__lane2_strm1_cntl          ( std__pe63__lane2_strm1_cntl       ),      
               .std__pe63__lane2_strm1_data          ( std__pe63__lane2_strm1_data       ),      
               .std__pe63__lane2_strm1_data_valid    ( std__pe63__lane2_strm1_data_valid ),      
               .std__pe63__lane2_strm1_data_mask     ( std__pe63__lane2_strm1_data_mask  ),      

               // PE 63, Lane 3                 
               .pe63__std__lane3_strm0_ready         ( pe63__std__lane3_strm0_ready      ),      
               .std__pe63__lane3_strm0_cntl          ( std__pe63__lane3_strm0_cntl       ),      
               .std__pe63__lane3_strm0_data          ( std__pe63__lane3_strm0_data       ),      
               .std__pe63__lane3_strm0_data_valid    ( std__pe63__lane3_strm0_data_valid ),      
               .std__pe63__lane3_strm0_data_mask     ( std__pe63__lane3_strm0_data_mask  ),      

               .pe63__std__lane3_strm1_ready         ( pe63__std__lane3_strm1_ready      ),      
               .std__pe63__lane3_strm1_cntl          ( std__pe63__lane3_strm1_cntl       ),      
               .std__pe63__lane3_strm1_data          ( std__pe63__lane3_strm1_data       ),      
               .std__pe63__lane3_strm1_data_valid    ( std__pe63__lane3_strm1_data_valid ),      
               .std__pe63__lane3_strm1_data_mask     ( std__pe63__lane3_strm1_data_mask  ),      

               // PE 63, Lane 4                 
               .pe63__std__lane4_strm0_ready         ( pe63__std__lane4_strm0_ready      ),      
               .std__pe63__lane4_strm0_cntl          ( std__pe63__lane4_strm0_cntl       ),      
               .std__pe63__lane4_strm0_data          ( std__pe63__lane4_strm0_data       ),      
               .std__pe63__lane4_strm0_data_valid    ( std__pe63__lane4_strm0_data_valid ),      
               .std__pe63__lane4_strm0_data_mask     ( std__pe63__lane4_strm0_data_mask  ),      

               .pe63__std__lane4_strm1_ready         ( pe63__std__lane4_strm1_ready      ),      
               .std__pe63__lane4_strm1_cntl          ( std__pe63__lane4_strm1_cntl       ),      
               .std__pe63__lane4_strm1_data          ( std__pe63__lane4_strm1_data       ),      
               .std__pe63__lane4_strm1_data_valid    ( std__pe63__lane4_strm1_data_valid ),      
               .std__pe63__lane4_strm1_data_mask     ( std__pe63__lane4_strm1_data_mask  ),      

               // PE 63, Lane 5                 
               .pe63__std__lane5_strm0_ready         ( pe63__std__lane5_strm0_ready      ),      
               .std__pe63__lane5_strm0_cntl          ( std__pe63__lane5_strm0_cntl       ),      
               .std__pe63__lane5_strm0_data          ( std__pe63__lane5_strm0_data       ),      
               .std__pe63__lane5_strm0_data_valid    ( std__pe63__lane5_strm0_data_valid ),      
               .std__pe63__lane5_strm0_data_mask     ( std__pe63__lane5_strm0_data_mask  ),      

               .pe63__std__lane5_strm1_ready         ( pe63__std__lane5_strm1_ready      ),      
               .std__pe63__lane5_strm1_cntl          ( std__pe63__lane5_strm1_cntl       ),      
               .std__pe63__lane5_strm1_data          ( std__pe63__lane5_strm1_data       ),      
               .std__pe63__lane5_strm1_data_valid    ( std__pe63__lane5_strm1_data_valid ),      
               .std__pe63__lane5_strm1_data_mask     ( std__pe63__lane5_strm1_data_mask  ),      

               // PE 63, Lane 6                 
               .pe63__std__lane6_strm0_ready         ( pe63__std__lane6_strm0_ready      ),      
               .std__pe63__lane6_strm0_cntl          ( std__pe63__lane6_strm0_cntl       ),      
               .std__pe63__lane6_strm0_data          ( std__pe63__lane6_strm0_data       ),      
               .std__pe63__lane6_strm0_data_valid    ( std__pe63__lane6_strm0_data_valid ),      
               .std__pe63__lane6_strm0_data_mask     ( std__pe63__lane6_strm0_data_mask  ),      

               .pe63__std__lane6_strm1_ready         ( pe63__std__lane6_strm1_ready      ),      
               .std__pe63__lane6_strm1_cntl          ( std__pe63__lane6_strm1_cntl       ),      
               .std__pe63__lane6_strm1_data          ( std__pe63__lane6_strm1_data       ),      
               .std__pe63__lane6_strm1_data_valid    ( std__pe63__lane6_strm1_data_valid ),      
               .std__pe63__lane6_strm1_data_mask     ( std__pe63__lane6_strm1_data_mask  ),      

               // PE 63, Lane 7                 
               .pe63__std__lane7_strm0_ready         ( pe63__std__lane7_strm0_ready      ),      
               .std__pe63__lane7_strm0_cntl          ( std__pe63__lane7_strm0_cntl       ),      
               .std__pe63__lane7_strm0_data          ( std__pe63__lane7_strm0_data       ),      
               .std__pe63__lane7_strm0_data_valid    ( std__pe63__lane7_strm0_data_valid ),      
               .std__pe63__lane7_strm0_data_mask     ( std__pe63__lane7_strm0_data_mask  ),      

               .pe63__std__lane7_strm1_ready         ( pe63__std__lane7_strm1_ready      ),      
               .std__pe63__lane7_strm1_cntl          ( std__pe63__lane7_strm1_cntl       ),      
               .std__pe63__lane7_strm1_data          ( std__pe63__lane7_strm1_data       ),      
               .std__pe63__lane7_strm1_data_valid    ( std__pe63__lane7_strm1_data_valid ),      
               .std__pe63__lane7_strm1_data_mask     ( std__pe63__lane7_strm1_data_mask  ),      

               // PE 63, Lane 8                 
               .pe63__std__lane8_strm0_ready         ( pe63__std__lane8_strm0_ready      ),      
               .std__pe63__lane8_strm0_cntl          ( std__pe63__lane8_strm0_cntl       ),      
               .std__pe63__lane8_strm0_data          ( std__pe63__lane8_strm0_data       ),      
               .std__pe63__lane8_strm0_data_valid    ( std__pe63__lane8_strm0_data_valid ),      
               .std__pe63__lane8_strm0_data_mask     ( std__pe63__lane8_strm0_data_mask  ),      

               .pe63__std__lane8_strm1_ready         ( pe63__std__lane8_strm1_ready      ),      
               .std__pe63__lane8_strm1_cntl          ( std__pe63__lane8_strm1_cntl       ),      
               .std__pe63__lane8_strm1_data          ( std__pe63__lane8_strm1_data       ),      
               .std__pe63__lane8_strm1_data_valid    ( std__pe63__lane8_strm1_data_valid ),      
               .std__pe63__lane8_strm1_data_mask     ( std__pe63__lane8_strm1_data_mask  ),      

               // PE 63, Lane 9                 
               .pe63__std__lane9_strm0_ready         ( pe63__std__lane9_strm0_ready      ),      
               .std__pe63__lane9_strm0_cntl          ( std__pe63__lane9_strm0_cntl       ),      
               .std__pe63__lane9_strm0_data          ( std__pe63__lane9_strm0_data       ),      
               .std__pe63__lane9_strm0_data_valid    ( std__pe63__lane9_strm0_data_valid ),      
               .std__pe63__lane9_strm0_data_mask     ( std__pe63__lane9_strm0_data_mask  ),      

               .pe63__std__lane9_strm1_ready         ( pe63__std__lane9_strm1_ready      ),      
               .std__pe63__lane9_strm1_cntl          ( std__pe63__lane9_strm1_cntl       ),      
               .std__pe63__lane9_strm1_data          ( std__pe63__lane9_strm1_data       ),      
               .std__pe63__lane9_strm1_data_valid    ( std__pe63__lane9_strm1_data_valid ),      
               .std__pe63__lane9_strm1_data_mask     ( std__pe63__lane9_strm1_data_mask  ),      

               // PE 63, Lane 10                 
               .pe63__std__lane10_strm0_ready         ( pe63__std__lane10_strm0_ready      ),      
               .std__pe63__lane10_strm0_cntl          ( std__pe63__lane10_strm0_cntl       ),      
               .std__pe63__lane10_strm0_data          ( std__pe63__lane10_strm0_data       ),      
               .std__pe63__lane10_strm0_data_valid    ( std__pe63__lane10_strm0_data_valid ),      
               .std__pe63__lane10_strm0_data_mask     ( std__pe63__lane10_strm0_data_mask  ),      

               .pe63__std__lane10_strm1_ready         ( pe63__std__lane10_strm1_ready      ),      
               .std__pe63__lane10_strm1_cntl          ( std__pe63__lane10_strm1_cntl       ),      
               .std__pe63__lane10_strm1_data          ( std__pe63__lane10_strm1_data       ),      
               .std__pe63__lane10_strm1_data_valid    ( std__pe63__lane10_strm1_data_valid ),      
               .std__pe63__lane10_strm1_data_mask     ( std__pe63__lane10_strm1_data_mask  ),      

               // PE 63, Lane 11                 
               .pe63__std__lane11_strm0_ready         ( pe63__std__lane11_strm0_ready      ),      
               .std__pe63__lane11_strm0_cntl          ( std__pe63__lane11_strm0_cntl       ),      
               .std__pe63__lane11_strm0_data          ( std__pe63__lane11_strm0_data       ),      
               .std__pe63__lane11_strm0_data_valid    ( std__pe63__lane11_strm0_data_valid ),      
               .std__pe63__lane11_strm0_data_mask     ( std__pe63__lane11_strm0_data_mask  ),      

               .pe63__std__lane11_strm1_ready         ( pe63__std__lane11_strm1_ready      ),      
               .std__pe63__lane11_strm1_cntl          ( std__pe63__lane11_strm1_cntl       ),      
               .std__pe63__lane11_strm1_data          ( std__pe63__lane11_strm1_data       ),      
               .std__pe63__lane11_strm1_data_valid    ( std__pe63__lane11_strm1_data_valid ),      
               .std__pe63__lane11_strm1_data_mask     ( std__pe63__lane11_strm1_data_mask  ),      

               // PE 63, Lane 12                 
               .pe63__std__lane12_strm0_ready         ( pe63__std__lane12_strm0_ready      ),      
               .std__pe63__lane12_strm0_cntl          ( std__pe63__lane12_strm0_cntl       ),      
               .std__pe63__lane12_strm0_data          ( std__pe63__lane12_strm0_data       ),      
               .std__pe63__lane12_strm0_data_valid    ( std__pe63__lane12_strm0_data_valid ),      
               .std__pe63__lane12_strm0_data_mask     ( std__pe63__lane12_strm0_data_mask  ),      

               .pe63__std__lane12_strm1_ready         ( pe63__std__lane12_strm1_ready      ),      
               .std__pe63__lane12_strm1_cntl          ( std__pe63__lane12_strm1_cntl       ),      
               .std__pe63__lane12_strm1_data          ( std__pe63__lane12_strm1_data       ),      
               .std__pe63__lane12_strm1_data_valid    ( std__pe63__lane12_strm1_data_valid ),      
               .std__pe63__lane12_strm1_data_mask     ( std__pe63__lane12_strm1_data_mask  ),      

               // PE 63, Lane 13                 
               .pe63__std__lane13_strm0_ready         ( pe63__std__lane13_strm0_ready      ),      
               .std__pe63__lane13_strm0_cntl          ( std__pe63__lane13_strm0_cntl       ),      
               .std__pe63__lane13_strm0_data          ( std__pe63__lane13_strm0_data       ),      
               .std__pe63__lane13_strm0_data_valid    ( std__pe63__lane13_strm0_data_valid ),      
               .std__pe63__lane13_strm0_data_mask     ( std__pe63__lane13_strm0_data_mask  ),      

               .pe63__std__lane13_strm1_ready         ( pe63__std__lane13_strm1_ready      ),      
               .std__pe63__lane13_strm1_cntl          ( std__pe63__lane13_strm1_cntl       ),      
               .std__pe63__lane13_strm1_data          ( std__pe63__lane13_strm1_data       ),      
               .std__pe63__lane13_strm1_data_valid    ( std__pe63__lane13_strm1_data_valid ),      
               .std__pe63__lane13_strm1_data_mask     ( std__pe63__lane13_strm1_data_mask  ),      

               // PE 63, Lane 14                 
               .pe63__std__lane14_strm0_ready         ( pe63__std__lane14_strm0_ready      ),      
               .std__pe63__lane14_strm0_cntl          ( std__pe63__lane14_strm0_cntl       ),      
               .std__pe63__lane14_strm0_data          ( std__pe63__lane14_strm0_data       ),      
               .std__pe63__lane14_strm0_data_valid    ( std__pe63__lane14_strm0_data_valid ),      
               .std__pe63__lane14_strm0_data_mask     ( std__pe63__lane14_strm0_data_mask  ),      

               .pe63__std__lane14_strm1_ready         ( pe63__std__lane14_strm1_ready      ),      
               .std__pe63__lane14_strm1_cntl          ( std__pe63__lane14_strm1_cntl       ),      
               .std__pe63__lane14_strm1_data          ( std__pe63__lane14_strm1_data       ),      
               .std__pe63__lane14_strm1_data_valid    ( std__pe63__lane14_strm1_data_valid ),      
               .std__pe63__lane14_strm1_data_mask     ( std__pe63__lane14_strm1_data_mask  ),      

               // PE 63, Lane 15                 
               .pe63__std__lane15_strm0_ready         ( pe63__std__lane15_strm0_ready      ),      
               .std__pe63__lane15_strm0_cntl          ( std__pe63__lane15_strm0_cntl       ),      
               .std__pe63__lane15_strm0_data          ( std__pe63__lane15_strm0_data       ),      
               .std__pe63__lane15_strm0_data_valid    ( std__pe63__lane15_strm0_data_valid ),      
               .std__pe63__lane15_strm0_data_mask     ( std__pe63__lane15_strm0_data_mask  ),      

               .pe63__std__lane15_strm1_ready         ( pe63__std__lane15_strm1_ready      ),      
               .std__pe63__lane15_strm1_cntl          ( std__pe63__lane15_strm1_cntl       ),      
               .std__pe63__lane15_strm1_data          ( std__pe63__lane15_strm1_data       ),      
               .std__pe63__lane15_strm1_data_valid    ( std__pe63__lane15_strm1_data_valid ),      
               .std__pe63__lane15_strm1_data_mask     ( std__pe63__lane15_strm1_data_mask  ),      

               // PE 63, Lane 16                 
               .pe63__std__lane16_strm0_ready         ( pe63__std__lane16_strm0_ready      ),      
               .std__pe63__lane16_strm0_cntl          ( std__pe63__lane16_strm0_cntl       ),      
               .std__pe63__lane16_strm0_data          ( std__pe63__lane16_strm0_data       ),      
               .std__pe63__lane16_strm0_data_valid    ( std__pe63__lane16_strm0_data_valid ),      
               .std__pe63__lane16_strm0_data_mask     ( std__pe63__lane16_strm0_data_mask  ),      

               .pe63__std__lane16_strm1_ready         ( pe63__std__lane16_strm1_ready      ),      
               .std__pe63__lane16_strm1_cntl          ( std__pe63__lane16_strm1_cntl       ),      
               .std__pe63__lane16_strm1_data          ( std__pe63__lane16_strm1_data       ),      
               .std__pe63__lane16_strm1_data_valid    ( std__pe63__lane16_strm1_data_valid ),      
               .std__pe63__lane16_strm1_data_mask     ( std__pe63__lane16_strm1_data_mask  ),      

               // PE 63, Lane 17                 
               .pe63__std__lane17_strm0_ready         ( pe63__std__lane17_strm0_ready      ),      
               .std__pe63__lane17_strm0_cntl          ( std__pe63__lane17_strm0_cntl       ),      
               .std__pe63__lane17_strm0_data          ( std__pe63__lane17_strm0_data       ),      
               .std__pe63__lane17_strm0_data_valid    ( std__pe63__lane17_strm0_data_valid ),      
               .std__pe63__lane17_strm0_data_mask     ( std__pe63__lane17_strm0_data_mask  ),      

               .pe63__std__lane17_strm1_ready         ( pe63__std__lane17_strm1_ready      ),      
               .std__pe63__lane17_strm1_cntl          ( std__pe63__lane17_strm1_cntl       ),      
               .std__pe63__lane17_strm1_data          ( std__pe63__lane17_strm1_data       ),      
               .std__pe63__lane17_strm1_data_valid    ( std__pe63__lane17_strm1_data_valid ),      
               .std__pe63__lane17_strm1_data_mask     ( std__pe63__lane17_strm1_data_mask  ),      

               // PE 63, Lane 18                 
               .pe63__std__lane18_strm0_ready         ( pe63__std__lane18_strm0_ready      ),      
               .std__pe63__lane18_strm0_cntl          ( std__pe63__lane18_strm0_cntl       ),      
               .std__pe63__lane18_strm0_data          ( std__pe63__lane18_strm0_data       ),      
               .std__pe63__lane18_strm0_data_valid    ( std__pe63__lane18_strm0_data_valid ),      
               .std__pe63__lane18_strm0_data_mask     ( std__pe63__lane18_strm0_data_mask  ),      

               .pe63__std__lane18_strm1_ready         ( pe63__std__lane18_strm1_ready      ),      
               .std__pe63__lane18_strm1_cntl          ( std__pe63__lane18_strm1_cntl       ),      
               .std__pe63__lane18_strm1_data          ( std__pe63__lane18_strm1_data       ),      
               .std__pe63__lane18_strm1_data_valid    ( std__pe63__lane18_strm1_data_valid ),      
               .std__pe63__lane18_strm1_data_mask     ( std__pe63__lane18_strm1_data_mask  ),      

               // PE 63, Lane 19                 
               .pe63__std__lane19_strm0_ready         ( pe63__std__lane19_strm0_ready      ),      
               .std__pe63__lane19_strm0_cntl          ( std__pe63__lane19_strm0_cntl       ),      
               .std__pe63__lane19_strm0_data          ( std__pe63__lane19_strm0_data       ),      
               .std__pe63__lane19_strm0_data_valid    ( std__pe63__lane19_strm0_data_valid ),      
               .std__pe63__lane19_strm0_data_mask     ( std__pe63__lane19_strm0_data_mask  ),      

               .pe63__std__lane19_strm1_ready         ( pe63__std__lane19_strm1_ready      ),      
               .std__pe63__lane19_strm1_cntl          ( std__pe63__lane19_strm1_cntl       ),      
               .std__pe63__lane19_strm1_data          ( std__pe63__lane19_strm1_data       ),      
               .std__pe63__lane19_strm1_data_valid    ( std__pe63__lane19_strm1_data_valid ),      
               .std__pe63__lane19_strm1_data_mask     ( std__pe63__lane19_strm1_data_mask  ),      

               // PE 63, Lane 20                 
               .pe63__std__lane20_strm0_ready         ( pe63__std__lane20_strm0_ready      ),      
               .std__pe63__lane20_strm0_cntl          ( std__pe63__lane20_strm0_cntl       ),      
               .std__pe63__lane20_strm0_data          ( std__pe63__lane20_strm0_data       ),      
               .std__pe63__lane20_strm0_data_valid    ( std__pe63__lane20_strm0_data_valid ),      
               .std__pe63__lane20_strm0_data_mask     ( std__pe63__lane20_strm0_data_mask  ),      

               .pe63__std__lane20_strm1_ready         ( pe63__std__lane20_strm1_ready      ),      
               .std__pe63__lane20_strm1_cntl          ( std__pe63__lane20_strm1_cntl       ),      
               .std__pe63__lane20_strm1_data          ( std__pe63__lane20_strm1_data       ),      
               .std__pe63__lane20_strm1_data_valid    ( std__pe63__lane20_strm1_data_valid ),      
               .std__pe63__lane20_strm1_data_mask     ( std__pe63__lane20_strm1_data_mask  ),      

               // PE 63, Lane 21                 
               .pe63__std__lane21_strm0_ready         ( pe63__std__lane21_strm0_ready      ),      
               .std__pe63__lane21_strm0_cntl          ( std__pe63__lane21_strm0_cntl       ),      
               .std__pe63__lane21_strm0_data          ( std__pe63__lane21_strm0_data       ),      
               .std__pe63__lane21_strm0_data_valid    ( std__pe63__lane21_strm0_data_valid ),      
               .std__pe63__lane21_strm0_data_mask     ( std__pe63__lane21_strm0_data_mask  ),      

               .pe63__std__lane21_strm1_ready         ( pe63__std__lane21_strm1_ready      ),      
               .std__pe63__lane21_strm1_cntl          ( std__pe63__lane21_strm1_cntl       ),      
               .std__pe63__lane21_strm1_data          ( std__pe63__lane21_strm1_data       ),      
               .std__pe63__lane21_strm1_data_valid    ( std__pe63__lane21_strm1_data_valid ),      
               .std__pe63__lane21_strm1_data_mask     ( std__pe63__lane21_strm1_data_mask  ),      

               // PE 63, Lane 22                 
               .pe63__std__lane22_strm0_ready         ( pe63__std__lane22_strm0_ready      ),      
               .std__pe63__lane22_strm0_cntl          ( std__pe63__lane22_strm0_cntl       ),      
               .std__pe63__lane22_strm0_data          ( std__pe63__lane22_strm0_data       ),      
               .std__pe63__lane22_strm0_data_valid    ( std__pe63__lane22_strm0_data_valid ),      
               .std__pe63__lane22_strm0_data_mask     ( std__pe63__lane22_strm0_data_mask  ),      

               .pe63__std__lane22_strm1_ready         ( pe63__std__lane22_strm1_ready      ),      
               .std__pe63__lane22_strm1_cntl          ( std__pe63__lane22_strm1_cntl       ),      
               .std__pe63__lane22_strm1_data          ( std__pe63__lane22_strm1_data       ),      
               .std__pe63__lane22_strm1_data_valid    ( std__pe63__lane22_strm1_data_valid ),      
               .std__pe63__lane22_strm1_data_mask     ( std__pe63__lane22_strm1_data_mask  ),      

               // PE 63, Lane 23                 
               .pe63__std__lane23_strm0_ready         ( pe63__std__lane23_strm0_ready      ),      
               .std__pe63__lane23_strm0_cntl          ( std__pe63__lane23_strm0_cntl       ),      
               .std__pe63__lane23_strm0_data          ( std__pe63__lane23_strm0_data       ),      
               .std__pe63__lane23_strm0_data_valid    ( std__pe63__lane23_strm0_data_valid ),      
               .std__pe63__lane23_strm0_data_mask     ( std__pe63__lane23_strm0_data_mask  ),      

               .pe63__std__lane23_strm1_ready         ( pe63__std__lane23_strm1_ready      ),      
               .std__pe63__lane23_strm1_cntl          ( std__pe63__lane23_strm1_cntl       ),      
               .std__pe63__lane23_strm1_data          ( std__pe63__lane23_strm1_data       ),      
               .std__pe63__lane23_strm1_data_valid    ( std__pe63__lane23_strm1_data_valid ),      
               .std__pe63__lane23_strm1_data_mask     ( std__pe63__lane23_strm1_data_mask  ),      

               // PE 63, Lane 24                 
               .pe63__std__lane24_strm0_ready         ( pe63__std__lane24_strm0_ready      ),      
               .std__pe63__lane24_strm0_cntl          ( std__pe63__lane24_strm0_cntl       ),      
               .std__pe63__lane24_strm0_data          ( std__pe63__lane24_strm0_data       ),      
               .std__pe63__lane24_strm0_data_valid    ( std__pe63__lane24_strm0_data_valid ),      
               .std__pe63__lane24_strm0_data_mask     ( std__pe63__lane24_strm0_data_mask  ),      

               .pe63__std__lane24_strm1_ready         ( pe63__std__lane24_strm1_ready      ),      
               .std__pe63__lane24_strm1_cntl          ( std__pe63__lane24_strm1_cntl       ),      
               .std__pe63__lane24_strm1_data          ( std__pe63__lane24_strm1_data       ),      
               .std__pe63__lane24_strm1_data_valid    ( std__pe63__lane24_strm1_data_valid ),      
               .std__pe63__lane24_strm1_data_mask     ( std__pe63__lane24_strm1_data_mask  ),      

               // PE 63, Lane 25                 
               .pe63__std__lane25_strm0_ready         ( pe63__std__lane25_strm0_ready      ),      
               .std__pe63__lane25_strm0_cntl          ( std__pe63__lane25_strm0_cntl       ),      
               .std__pe63__lane25_strm0_data          ( std__pe63__lane25_strm0_data       ),      
               .std__pe63__lane25_strm0_data_valid    ( std__pe63__lane25_strm0_data_valid ),      
               .std__pe63__lane25_strm0_data_mask     ( std__pe63__lane25_strm0_data_mask  ),      

               .pe63__std__lane25_strm1_ready         ( pe63__std__lane25_strm1_ready      ),      
               .std__pe63__lane25_strm1_cntl          ( std__pe63__lane25_strm1_cntl       ),      
               .std__pe63__lane25_strm1_data          ( std__pe63__lane25_strm1_data       ),      
               .std__pe63__lane25_strm1_data_valid    ( std__pe63__lane25_strm1_data_valid ),      
               .std__pe63__lane25_strm1_data_mask     ( std__pe63__lane25_strm1_data_mask  ),      

               // PE 63, Lane 26                 
               .pe63__std__lane26_strm0_ready         ( pe63__std__lane26_strm0_ready      ),      
               .std__pe63__lane26_strm0_cntl          ( std__pe63__lane26_strm0_cntl       ),      
               .std__pe63__lane26_strm0_data          ( std__pe63__lane26_strm0_data       ),      
               .std__pe63__lane26_strm0_data_valid    ( std__pe63__lane26_strm0_data_valid ),      
               .std__pe63__lane26_strm0_data_mask     ( std__pe63__lane26_strm0_data_mask  ),      

               .pe63__std__lane26_strm1_ready         ( pe63__std__lane26_strm1_ready      ),      
               .std__pe63__lane26_strm1_cntl          ( std__pe63__lane26_strm1_cntl       ),      
               .std__pe63__lane26_strm1_data          ( std__pe63__lane26_strm1_data       ),      
               .std__pe63__lane26_strm1_data_valid    ( std__pe63__lane26_strm1_data_valid ),      
               .std__pe63__lane26_strm1_data_mask     ( std__pe63__lane26_strm1_data_mask  ),      

               // PE 63, Lane 27                 
               .pe63__std__lane27_strm0_ready         ( pe63__std__lane27_strm0_ready      ),      
               .std__pe63__lane27_strm0_cntl          ( std__pe63__lane27_strm0_cntl       ),      
               .std__pe63__lane27_strm0_data          ( std__pe63__lane27_strm0_data       ),      
               .std__pe63__lane27_strm0_data_valid    ( std__pe63__lane27_strm0_data_valid ),      
               .std__pe63__lane27_strm0_data_mask     ( std__pe63__lane27_strm0_data_mask  ),      

               .pe63__std__lane27_strm1_ready         ( pe63__std__lane27_strm1_ready      ),      
               .std__pe63__lane27_strm1_cntl          ( std__pe63__lane27_strm1_cntl       ),      
               .std__pe63__lane27_strm1_data          ( std__pe63__lane27_strm1_data       ),      
               .std__pe63__lane27_strm1_data_valid    ( std__pe63__lane27_strm1_data_valid ),      
               .std__pe63__lane27_strm1_data_mask     ( std__pe63__lane27_strm1_data_mask  ),      

               // PE 63, Lane 28                 
               .pe63__std__lane28_strm0_ready         ( pe63__std__lane28_strm0_ready      ),      
               .std__pe63__lane28_strm0_cntl          ( std__pe63__lane28_strm0_cntl       ),      
               .std__pe63__lane28_strm0_data          ( std__pe63__lane28_strm0_data       ),      
               .std__pe63__lane28_strm0_data_valid    ( std__pe63__lane28_strm0_data_valid ),      
               .std__pe63__lane28_strm0_data_mask     ( std__pe63__lane28_strm0_data_mask  ),      

               .pe63__std__lane28_strm1_ready         ( pe63__std__lane28_strm1_ready      ),      
               .std__pe63__lane28_strm1_cntl          ( std__pe63__lane28_strm1_cntl       ),      
               .std__pe63__lane28_strm1_data          ( std__pe63__lane28_strm1_data       ),      
               .std__pe63__lane28_strm1_data_valid    ( std__pe63__lane28_strm1_data_valid ),      
               .std__pe63__lane28_strm1_data_mask     ( std__pe63__lane28_strm1_data_mask  ),      

               // PE 63, Lane 29                 
               .pe63__std__lane29_strm0_ready         ( pe63__std__lane29_strm0_ready      ),      
               .std__pe63__lane29_strm0_cntl          ( std__pe63__lane29_strm0_cntl       ),      
               .std__pe63__lane29_strm0_data          ( std__pe63__lane29_strm0_data       ),      
               .std__pe63__lane29_strm0_data_valid    ( std__pe63__lane29_strm0_data_valid ),      
               .std__pe63__lane29_strm0_data_mask     ( std__pe63__lane29_strm0_data_mask  ),      

               .pe63__std__lane29_strm1_ready         ( pe63__std__lane29_strm1_ready      ),      
               .std__pe63__lane29_strm1_cntl          ( std__pe63__lane29_strm1_cntl       ),      
               .std__pe63__lane29_strm1_data          ( std__pe63__lane29_strm1_data       ),      
               .std__pe63__lane29_strm1_data_valid    ( std__pe63__lane29_strm1_data_valid ),      
               .std__pe63__lane29_strm1_data_mask     ( std__pe63__lane29_strm1_data_mask  ),      

               // PE 63, Lane 30                 
               .pe63__std__lane30_strm0_ready         ( pe63__std__lane30_strm0_ready      ),      
               .std__pe63__lane30_strm0_cntl          ( std__pe63__lane30_strm0_cntl       ),      
               .std__pe63__lane30_strm0_data          ( std__pe63__lane30_strm0_data       ),      
               .std__pe63__lane30_strm0_data_valid    ( std__pe63__lane30_strm0_data_valid ),      
               .std__pe63__lane30_strm0_data_mask     ( std__pe63__lane30_strm0_data_mask  ),      

               .pe63__std__lane30_strm1_ready         ( pe63__std__lane30_strm1_ready      ),      
               .std__pe63__lane30_strm1_cntl          ( std__pe63__lane30_strm1_cntl       ),      
               .std__pe63__lane30_strm1_data          ( std__pe63__lane30_strm1_data       ),      
               .std__pe63__lane30_strm1_data_valid    ( std__pe63__lane30_strm1_data_valid ),      
               .std__pe63__lane30_strm1_data_mask     ( std__pe63__lane30_strm1_data_mask  ),      

               // PE 63, Lane 31                 
               .pe63__std__lane31_strm0_ready         ( pe63__std__lane31_strm0_ready      ),      
               .std__pe63__lane31_strm0_cntl          ( std__pe63__lane31_strm0_cntl       ),      
               .std__pe63__lane31_strm0_data          ( std__pe63__lane31_strm0_data       ),      
               .std__pe63__lane31_strm0_data_valid    ( std__pe63__lane31_strm0_data_valid ),      
               .std__pe63__lane31_strm0_data_mask     ( std__pe63__lane31_strm0_data_mask  ),      

               .pe63__std__lane31_strm1_ready         ( pe63__std__lane31_strm1_ready      ),      
               .std__pe63__lane31_strm1_cntl          ( std__pe63__lane31_strm1_cntl       ),      
               .std__pe63__lane31_strm1_data          ( std__pe63__lane31_strm1_data       ),      
               .std__pe63__lane31_strm1_data_valid    ( std__pe63__lane31_strm1_data_valid ),      
               .std__pe63__lane31_strm1_data_mask     ( std__pe63__lane31_strm1_data_mask  ),      
