
`define NOC_CONT_MGR0_PORT0_DESTINATION_MGR_BITMASK  'b1111111011111110111111101111111011111110111111101111111011111110
`define NOC_CONT_MGR0_PORT1_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000001000000010000000100000000
`define NOC_CONT_MGR0_PORT2_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR0_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR1_PORT0_DESTINATION_MGR_BITMASK  'b1111110011111100111111001111110011111100111111001111110011111100
`define NOC_CONT_MGR1_PORT1_DESTINATION_MGR_BITMASK  'b0000001000000010000000100000001000000010000000100000001000000000
`define NOC_CONT_MGR1_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000001000000010000000100000001
`define NOC_CONT_MGR1_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR2_PORT0_DESTINATION_MGR_BITMASK  'b1111100011111000111110001111100011111000111110001111100011111000
`define NOC_CONT_MGR2_PORT1_DESTINATION_MGR_BITMASK  'b0000010000000100000001000000010000000100000001000000010000000000
`define NOC_CONT_MGR2_PORT2_DESTINATION_MGR_BITMASK  'b0000001100000011000000110000001100000011000000110000001100000011
`define NOC_CONT_MGR2_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR3_PORT0_DESTINATION_MGR_BITMASK  'b1111000011110000111100001111000011110000111100001111000011110000
`define NOC_CONT_MGR3_PORT1_DESTINATION_MGR_BITMASK  'b0000100000001000000010000000100000001000000010000000100000000000
`define NOC_CONT_MGR3_PORT2_DESTINATION_MGR_BITMASK  'b0000011100000111000001110000011100000111000001110000011100000111
`define NOC_CONT_MGR3_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR4_PORT0_DESTINATION_MGR_BITMASK  'b1110000011100000111000001110000011100000111000001110000011100000
`define NOC_CONT_MGR4_PORT1_DESTINATION_MGR_BITMASK  'b0001000000010000000100000001000000010000000100000001000000000000
`define NOC_CONT_MGR4_PORT2_DESTINATION_MGR_BITMASK  'b0000111100001111000011110000111100001111000011110000111100001111
`define NOC_CONT_MGR4_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR5_PORT0_DESTINATION_MGR_BITMASK  'b1100000011000000110000001100000011000000110000001100000011000000
`define NOC_CONT_MGR5_PORT1_DESTINATION_MGR_BITMASK  'b0010000000100000001000000010000000100000001000000010000000000000
`define NOC_CONT_MGR5_PORT2_DESTINATION_MGR_BITMASK  'b0001111100011111000111110001111100011111000111110001111100011111
`define NOC_CONT_MGR5_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR6_PORT0_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000010000000100000001000000010000000
`define NOC_CONT_MGR6_PORT1_DESTINATION_MGR_BITMASK  'b0100000001000000010000000100000001000000010000000100000000000000
`define NOC_CONT_MGR6_PORT2_DESTINATION_MGR_BITMASK  'b0011111100111111001111110011111100111111001111110011111100111111
`define NOC_CONT_MGR6_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR7_PORT0_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000010000000100000001000000000000000
`define NOC_CONT_MGR7_PORT1_DESTINATION_MGR_BITMASK  'b0111111101111111011111110111111101111111011111110111111101111111
`define NOC_CONT_MGR7_PORT2_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR7_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR8_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR8_PORT1_DESTINATION_MGR_BITMASK  'b1111111011111110111111101111111011111110111111101111111000000000
`define NOC_CONT_MGR8_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000001000000010000000000000000
`define NOC_CONT_MGR8_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR9_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR9_PORT1_DESTINATION_MGR_BITMASK  'b1111110011111100111111001111110011111100111111001111110000000000
`define NOC_CONT_MGR9_PORT2_DESTINATION_MGR_BITMASK  'b0000001000000010000000100000001000000010000000100000000000000000
`define NOC_CONT_MGR9_PORT3_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000001000000010000000100000000
`define NOC_CONT_MGR10_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR10_PORT1_DESTINATION_MGR_BITMASK  'b1111100011111000111110001111100011111000111110001111100000000000
`define NOC_CONT_MGR10_PORT2_DESTINATION_MGR_BITMASK  'b0000010000000100000001000000010000000100000001000000000000000000
`define NOC_CONT_MGR10_PORT3_DESTINATION_MGR_BITMASK  'b0000001100000011000000110000001100000011000000110000001100000000
`define NOC_CONT_MGR11_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR11_PORT1_DESTINATION_MGR_BITMASK  'b1111000011110000111100001111000011110000111100001111000000000000
`define NOC_CONT_MGR11_PORT2_DESTINATION_MGR_BITMASK  'b0000100000001000000010000000100000001000000010000000000000000000
`define NOC_CONT_MGR11_PORT3_DESTINATION_MGR_BITMASK  'b0000011100000111000001110000011100000111000001110000011100000000
`define NOC_CONT_MGR12_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR12_PORT1_DESTINATION_MGR_BITMASK  'b1110000011100000111000001110000011100000111000001110000000000000
`define NOC_CONT_MGR12_PORT2_DESTINATION_MGR_BITMASK  'b0001000000010000000100000001000000010000000100000000000000000000
`define NOC_CONT_MGR12_PORT3_DESTINATION_MGR_BITMASK  'b0000111100001111000011110000111100001111000011110000111100000000
`define NOC_CONT_MGR13_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR13_PORT1_DESTINATION_MGR_BITMASK  'b1100000011000000110000001100000011000000110000001100000000000000
`define NOC_CONT_MGR13_PORT2_DESTINATION_MGR_BITMASK  'b0010000000100000001000000010000000100000001000000000000000000000
`define NOC_CONT_MGR13_PORT3_DESTINATION_MGR_BITMASK  'b0001111100011111000111110001111100011111000111110001111100000000
`define NOC_CONT_MGR14_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR14_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000010000000100000001000000000000000
`define NOC_CONT_MGR14_PORT2_DESTINATION_MGR_BITMASK  'b0100000001000000010000000100000001000000010000000000000000000000
`define NOC_CONT_MGR14_PORT3_DESTINATION_MGR_BITMASK  'b0011111100111111001111110011111100111111001111110011111100000000
`define NOC_CONT_MGR15_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000000000000011111111
`define NOC_CONT_MGR15_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000010000000100000000000000000000000
`define NOC_CONT_MGR15_PORT2_DESTINATION_MGR_BITMASK  'b0111111101111111011111110111111101111111011111110111111100000000
`define NOC_CONT_MGR15_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR16_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR16_PORT1_DESTINATION_MGR_BITMASK  'b1111111011111110111111101111111011111110111111100000000000000000
`define NOC_CONT_MGR16_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000001000000000000000000000000
`define NOC_CONT_MGR16_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR17_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR17_PORT1_DESTINATION_MGR_BITMASK  'b1111110011111100111111001111110011111100111111000000000000000000
`define NOC_CONT_MGR17_PORT2_DESTINATION_MGR_BITMASK  'b0000001000000010000000100000001000000010000000000000000000000000
`define NOC_CONT_MGR17_PORT3_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000001000000010000000000000000
`define NOC_CONT_MGR18_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR18_PORT1_DESTINATION_MGR_BITMASK  'b1111100011111000111110001111100011111000111110000000000000000000
`define NOC_CONT_MGR18_PORT2_DESTINATION_MGR_BITMASK  'b0000010000000100000001000000010000000100000000000000000000000000
`define NOC_CONT_MGR18_PORT3_DESTINATION_MGR_BITMASK  'b0000001100000011000000110000001100000011000000110000000000000000
`define NOC_CONT_MGR19_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR19_PORT1_DESTINATION_MGR_BITMASK  'b1111000011110000111100001111000011110000111100000000000000000000
`define NOC_CONT_MGR19_PORT2_DESTINATION_MGR_BITMASK  'b0000100000001000000010000000100000001000000000000000000000000000
`define NOC_CONT_MGR19_PORT3_DESTINATION_MGR_BITMASK  'b0000011100000111000001110000011100000111000001110000000000000000
`define NOC_CONT_MGR20_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR20_PORT1_DESTINATION_MGR_BITMASK  'b1110000011100000111000001110000011100000111000000000000000000000
`define NOC_CONT_MGR20_PORT2_DESTINATION_MGR_BITMASK  'b0001000000010000000100000001000000010000000000000000000000000000
`define NOC_CONT_MGR20_PORT3_DESTINATION_MGR_BITMASK  'b0000111100001111000011110000111100001111000011110000000000000000
`define NOC_CONT_MGR21_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR21_PORT1_DESTINATION_MGR_BITMASK  'b1100000011000000110000001100000011000000110000000000000000000000
`define NOC_CONT_MGR21_PORT2_DESTINATION_MGR_BITMASK  'b0010000000100000001000000010000000100000000000000000000000000000
`define NOC_CONT_MGR21_PORT3_DESTINATION_MGR_BITMASK  'b0001111100011111000111110001111100011111000111110000000000000000
`define NOC_CONT_MGR22_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR22_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000010000000100000000000000000000000
`define NOC_CONT_MGR22_PORT2_DESTINATION_MGR_BITMASK  'b0100000001000000010000000100000001000000000000000000000000000000
`define NOC_CONT_MGR22_PORT3_DESTINATION_MGR_BITMASK  'b0011111100111111001111110011111100111111001111110000000000000000
`define NOC_CONT_MGR23_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000000000001111111111111111
`define NOC_CONT_MGR23_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000010000000000000000000000000000000
`define NOC_CONT_MGR23_PORT2_DESTINATION_MGR_BITMASK  'b0111111101111111011111110111111101111111011111110000000000000000
`define NOC_CONT_MGR23_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR24_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR24_PORT1_DESTINATION_MGR_BITMASK  'b1111111011111110111111101111111011111110000000000000000000000000
`define NOC_CONT_MGR24_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000000000000000000000000000000
`define NOC_CONT_MGR24_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR25_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR25_PORT1_DESTINATION_MGR_BITMASK  'b1111110011111100111111001111110011111100000000000000000000000000
`define NOC_CONT_MGR25_PORT2_DESTINATION_MGR_BITMASK  'b0000001000000010000000100000001000000000000000000000000000000000
`define NOC_CONT_MGR25_PORT3_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000001000000000000000000000000
`define NOC_CONT_MGR26_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR26_PORT1_DESTINATION_MGR_BITMASK  'b1111100011111000111110001111100011111000000000000000000000000000
`define NOC_CONT_MGR26_PORT2_DESTINATION_MGR_BITMASK  'b0000010000000100000001000000010000000000000000000000000000000000
`define NOC_CONT_MGR26_PORT3_DESTINATION_MGR_BITMASK  'b0000001100000011000000110000001100000011000000000000000000000000
`define NOC_CONT_MGR27_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR27_PORT1_DESTINATION_MGR_BITMASK  'b1111000011110000111100001111000011110000000000000000000000000000
`define NOC_CONT_MGR27_PORT2_DESTINATION_MGR_BITMASK  'b0000100000001000000010000000100000000000000000000000000000000000
`define NOC_CONT_MGR27_PORT3_DESTINATION_MGR_BITMASK  'b0000011100000111000001110000011100000111000000000000000000000000
`define NOC_CONT_MGR28_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR28_PORT1_DESTINATION_MGR_BITMASK  'b1110000011100000111000001110000011100000000000000000000000000000
`define NOC_CONT_MGR28_PORT2_DESTINATION_MGR_BITMASK  'b0001000000010000000100000001000000000000000000000000000000000000
`define NOC_CONT_MGR28_PORT3_DESTINATION_MGR_BITMASK  'b0000111100001111000011110000111100001111000000000000000000000000
`define NOC_CONT_MGR29_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR29_PORT1_DESTINATION_MGR_BITMASK  'b1100000011000000110000001100000011000000000000000000000000000000
`define NOC_CONT_MGR29_PORT2_DESTINATION_MGR_BITMASK  'b0010000000100000001000000010000000000000000000000000000000000000
`define NOC_CONT_MGR29_PORT3_DESTINATION_MGR_BITMASK  'b0001111100011111000111110001111100011111000000000000000000000000
`define NOC_CONT_MGR30_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR30_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000010000000000000000000000000000000
`define NOC_CONT_MGR30_PORT2_DESTINATION_MGR_BITMASK  'b0100000001000000010000000100000000000000000000000000000000000000
`define NOC_CONT_MGR30_PORT3_DESTINATION_MGR_BITMASK  'b0011111100111111001111110011111100111111000000000000000000000000
`define NOC_CONT_MGR31_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000000000000111111111111111111111111
`define NOC_CONT_MGR31_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000000000000000000000000000000000000
`define NOC_CONT_MGR31_PORT2_DESTINATION_MGR_BITMASK  'b0111111101111111011111110111111101111111000000000000000000000000
`define NOC_CONT_MGR31_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR32_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR32_PORT1_DESTINATION_MGR_BITMASK  'b1111111011111110111111101111111000000000000000000000000000000000
`define NOC_CONT_MGR32_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000000000000000000000000000000000000
`define NOC_CONT_MGR32_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR33_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR33_PORT1_DESTINATION_MGR_BITMASK  'b1111110011111100111111001111110000000000000000000000000000000000
`define NOC_CONT_MGR33_PORT2_DESTINATION_MGR_BITMASK  'b0000001000000010000000100000000000000000000000000000000000000000
`define NOC_CONT_MGR33_PORT3_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000100000000000000000000000000000000
`define NOC_CONT_MGR34_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR34_PORT1_DESTINATION_MGR_BITMASK  'b1111100011111000111110001111100000000000000000000000000000000000
`define NOC_CONT_MGR34_PORT2_DESTINATION_MGR_BITMASK  'b0000010000000100000001000000000000000000000000000000000000000000
`define NOC_CONT_MGR34_PORT3_DESTINATION_MGR_BITMASK  'b0000001100000011000000110000001100000000000000000000000000000000
`define NOC_CONT_MGR35_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR35_PORT1_DESTINATION_MGR_BITMASK  'b1111000011110000111100001111000000000000000000000000000000000000
`define NOC_CONT_MGR35_PORT2_DESTINATION_MGR_BITMASK  'b0000100000001000000010000000000000000000000000000000000000000000
`define NOC_CONT_MGR35_PORT3_DESTINATION_MGR_BITMASK  'b0000011100000111000001110000011100000000000000000000000000000000
`define NOC_CONT_MGR36_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR36_PORT1_DESTINATION_MGR_BITMASK  'b1110000011100000111000001110000000000000000000000000000000000000
`define NOC_CONT_MGR36_PORT2_DESTINATION_MGR_BITMASK  'b0001000000010000000100000000000000000000000000000000000000000000
`define NOC_CONT_MGR36_PORT3_DESTINATION_MGR_BITMASK  'b0000111100001111000011110000111100000000000000000000000000000000
`define NOC_CONT_MGR37_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR37_PORT1_DESTINATION_MGR_BITMASK  'b1100000011000000110000001100000000000000000000000000000000000000
`define NOC_CONT_MGR37_PORT2_DESTINATION_MGR_BITMASK  'b0010000000100000001000000000000000000000000000000000000000000000
`define NOC_CONT_MGR37_PORT3_DESTINATION_MGR_BITMASK  'b0001111100011111000111110001111100000000000000000000000000000000
`define NOC_CONT_MGR38_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR38_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000001000000000000000000000000000000000000000
`define NOC_CONT_MGR38_PORT2_DESTINATION_MGR_BITMASK  'b0100000001000000010000000000000000000000000000000000000000000000
`define NOC_CONT_MGR38_PORT3_DESTINATION_MGR_BITMASK  'b0011111100111111001111110011111100000000000000000000000000000000
`define NOC_CONT_MGR39_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000000000000011111111111111111111111111111111
`define NOC_CONT_MGR39_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000000000000000000000000000000000000000000000
`define NOC_CONT_MGR39_PORT2_DESTINATION_MGR_BITMASK  'b0111111101111111011111110111111100000000000000000000000000000000
`define NOC_CONT_MGR39_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR40_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR40_PORT1_DESTINATION_MGR_BITMASK  'b1111111011111110111111100000000000000000000000000000000000000000
`define NOC_CONT_MGR40_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000001000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR40_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR41_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR41_PORT1_DESTINATION_MGR_BITMASK  'b1111110011111100111111000000000000000000000000000000000000000000
`define NOC_CONT_MGR41_PORT2_DESTINATION_MGR_BITMASK  'b0000001000000010000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR41_PORT3_DESTINATION_MGR_BITMASK  'b0000000100000001000000010000000000000000000000000000000000000000
`define NOC_CONT_MGR42_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR42_PORT1_DESTINATION_MGR_BITMASK  'b1111100011111000111110000000000000000000000000000000000000000000
`define NOC_CONT_MGR42_PORT2_DESTINATION_MGR_BITMASK  'b0000010000000100000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR42_PORT3_DESTINATION_MGR_BITMASK  'b0000001100000011000000110000000000000000000000000000000000000000
`define NOC_CONT_MGR43_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR43_PORT1_DESTINATION_MGR_BITMASK  'b1111000011110000111100000000000000000000000000000000000000000000
`define NOC_CONT_MGR43_PORT2_DESTINATION_MGR_BITMASK  'b0000100000001000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR43_PORT3_DESTINATION_MGR_BITMASK  'b0000011100000111000001110000000000000000000000000000000000000000
`define NOC_CONT_MGR44_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR44_PORT1_DESTINATION_MGR_BITMASK  'b1110000011100000111000000000000000000000000000000000000000000000
`define NOC_CONT_MGR44_PORT2_DESTINATION_MGR_BITMASK  'b0001000000010000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR44_PORT3_DESTINATION_MGR_BITMASK  'b0000111100001111000011110000000000000000000000000000000000000000
`define NOC_CONT_MGR45_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR45_PORT1_DESTINATION_MGR_BITMASK  'b1100000011000000110000000000000000000000000000000000000000000000
`define NOC_CONT_MGR45_PORT2_DESTINATION_MGR_BITMASK  'b0010000000100000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR45_PORT3_DESTINATION_MGR_BITMASK  'b0001111100011111000111110000000000000000000000000000000000000000
`define NOC_CONT_MGR46_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR46_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000100000000000000000000000000000000000000000000000
`define NOC_CONT_MGR46_PORT2_DESTINATION_MGR_BITMASK  'b0100000001000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR46_PORT3_DESTINATION_MGR_BITMASK  'b0011111100111111001111110000000000000000000000000000000000000000
`define NOC_CONT_MGR47_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000000000001111111111111111111111111111111111111111
`define NOC_CONT_MGR47_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR47_PORT2_DESTINATION_MGR_BITMASK  'b0111111101111111011111110000000000000000000000000000000000000000
`define NOC_CONT_MGR47_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR48_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR48_PORT1_DESTINATION_MGR_BITMASK  'b1111111011111110000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR48_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR48_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR49_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR49_PORT1_DESTINATION_MGR_BITMASK  'b1111110011111100000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR49_PORT2_DESTINATION_MGR_BITMASK  'b0000001000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR49_PORT3_DESTINATION_MGR_BITMASK  'b0000000100000001000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR50_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR50_PORT1_DESTINATION_MGR_BITMASK  'b1111100011111000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR50_PORT2_DESTINATION_MGR_BITMASK  'b0000010000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR50_PORT3_DESTINATION_MGR_BITMASK  'b0000001100000011000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR51_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR51_PORT1_DESTINATION_MGR_BITMASK  'b1111000011110000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR51_PORT2_DESTINATION_MGR_BITMASK  'b0000100000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR51_PORT3_DESTINATION_MGR_BITMASK  'b0000011100000111000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR52_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR52_PORT1_DESTINATION_MGR_BITMASK  'b1110000011100000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR52_PORT2_DESTINATION_MGR_BITMASK  'b0001000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR52_PORT3_DESTINATION_MGR_BITMASK  'b0000111100001111000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR53_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR53_PORT1_DESTINATION_MGR_BITMASK  'b1100000011000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR53_PORT2_DESTINATION_MGR_BITMASK  'b0010000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR53_PORT3_DESTINATION_MGR_BITMASK  'b0001111100011111000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR54_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR54_PORT1_DESTINATION_MGR_BITMASK  'b1000000010000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR54_PORT2_DESTINATION_MGR_BITMASK  'b0100000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR54_PORT3_DESTINATION_MGR_BITMASK  'b0011111100111111000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR55_PORT0_DESTINATION_MGR_BITMASK  'b0000000000000000111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR55_PORT1_DESTINATION_MGR_BITMASK  'b1000000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR55_PORT2_DESTINATION_MGR_BITMASK  'b0111111101111111000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR55_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR56_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR56_PORT1_DESTINATION_MGR_BITMASK  'b1111111000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR56_PORT2_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR56_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR57_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR57_PORT1_DESTINATION_MGR_BITMASK  'b1111110000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR57_PORT2_DESTINATION_MGR_BITMASK  'b0000000100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR57_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR58_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR58_PORT1_DESTINATION_MGR_BITMASK  'b1111100000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR58_PORT2_DESTINATION_MGR_BITMASK  'b0000001100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR58_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR59_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR59_PORT1_DESTINATION_MGR_BITMASK  'b1111000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR59_PORT2_DESTINATION_MGR_BITMASK  'b0000011100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR59_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR60_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR60_PORT1_DESTINATION_MGR_BITMASK  'b1110000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR60_PORT2_DESTINATION_MGR_BITMASK  'b0000111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR60_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR61_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR61_PORT1_DESTINATION_MGR_BITMASK  'b1100000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR61_PORT2_DESTINATION_MGR_BITMASK  'b0001111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR61_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR62_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR62_PORT1_DESTINATION_MGR_BITMASK  'b1000000000000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR62_PORT2_DESTINATION_MGR_BITMASK  'b0011111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR62_PORT3_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR63_PORT0_DESTINATION_MGR_BITMASK  'b0000000011111111111111111111111111111111111111111111111111111111
`define NOC_CONT_MGR63_PORT1_DESTINATION_MGR_BITMASK  'b0111111100000000000000000000000000000000000000000000000000000000
`define NOC_CONT_MGR63_PORT2_DESTINATION_MGR_BITMASK  'd0
`define NOC_CONT_MGR63_PORT3_DESTINATION_MGR_BITMASK  'd0
