
      scntl__sdp__lane0_stOp_operation, 
      scntl__sdp__lane1_stOp_operation, 
      scntl__sdp__lane2_stOp_operation, 
      scntl__sdp__lane3_stOp_operation, 
      scntl__sdp__lane4_stOp_operation, 
      scntl__sdp__lane5_stOp_operation, 
      scntl__sdp__lane6_stOp_operation, 
      scntl__sdp__lane7_stOp_operation, 
      scntl__sdp__lane8_stOp_operation, 
      scntl__sdp__lane9_stOp_operation, 
      scntl__sdp__lane10_stOp_operation, 
      scntl__sdp__lane11_stOp_operation, 
      scntl__sdp__lane12_stOp_operation, 
      scntl__sdp__lane13_stOp_operation, 
      scntl__sdp__lane14_stOp_operation, 
      scntl__sdp__lane15_stOp_operation, 
      scntl__sdp__lane16_stOp_operation, 
      scntl__sdp__lane17_stOp_operation, 
      scntl__sdp__lane18_stOp_operation, 
      scntl__sdp__lane19_stOp_operation, 
      scntl__sdp__lane20_stOp_operation, 
      scntl__sdp__lane21_stOp_operation, 
      scntl__sdp__lane22_stOp_operation, 
      scntl__sdp__lane23_stOp_operation, 
      scntl__sdp__lane24_stOp_operation, 
      scntl__sdp__lane25_stOp_operation, 
      scntl__sdp__lane26_stOp_operation, 
      scntl__sdp__lane27_stOp_operation, 
      scntl__sdp__lane28_stOp_operation, 
      scntl__sdp__lane29_stOp_operation, 
      scntl__sdp__lane30_stOp_operation, 
      scntl__sdp__lane31_stOp_operation, 

      scntl__sdp__lane0_dma_operation, 
      scntl__sdp__lane1_dma_operation, 
      scntl__sdp__lane2_dma_operation, 
      scntl__sdp__lane3_dma_operation, 
      scntl__sdp__lane4_dma_operation, 
      scntl__sdp__lane5_dma_operation, 
      scntl__sdp__lane6_dma_operation, 
      scntl__sdp__lane7_dma_operation, 
      scntl__sdp__lane8_dma_operation, 
      scntl__sdp__lane9_dma_operation, 
      scntl__sdp__lane10_dma_operation, 
      scntl__sdp__lane11_dma_operation, 
      scntl__sdp__lane12_dma_operation, 
      scntl__sdp__lane13_dma_operation, 
      scntl__sdp__lane14_dma_operation, 
      scntl__sdp__lane15_dma_operation, 
      scntl__sdp__lane16_dma_operation, 
      scntl__sdp__lane17_dma_operation, 
      scntl__sdp__lane18_dma_operation, 
      scntl__sdp__lane19_dma_operation, 
      scntl__sdp__lane20_dma_operation, 
      scntl__sdp__lane21_dma_operation, 
      scntl__sdp__lane22_dma_operation, 
      scntl__sdp__lane23_dma_operation, 
      scntl__sdp__lane24_dma_operation, 
      scntl__sdp__lane25_dma_operation, 
      scntl__sdp__lane26_dma_operation, 
      scntl__sdp__lane27_dma_operation, 
      scntl__sdp__lane28_dma_operation, 
      scntl__sdp__lane29_dma_operation, 
      scntl__sdp__lane30_dma_operation, 
      scntl__sdp__lane31_dma_operation, 

      scntl__sdp__lane0_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane0_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane0_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane0_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane0_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane0_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane0_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane0_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane0_type0                      ,                                       
      scntl__sdp__lane0_num_of_types0              ,                                       
      scntl__sdp__lane1_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane1_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane1_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane1_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane1_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane1_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane1_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane1_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane1_type0                      ,                                       
      scntl__sdp__lane1_num_of_types0              ,                                       
      scntl__sdp__lane2_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane2_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane2_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane2_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane2_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane2_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane2_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane2_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane2_type0                      ,                                       
      scntl__sdp__lane2_num_of_types0              ,                                       
      scntl__sdp__lane3_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane3_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane3_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane3_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane3_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane3_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane3_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane3_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane3_type0                      ,                                       
      scntl__sdp__lane3_num_of_types0              ,                                       
      scntl__sdp__lane4_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane4_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane4_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane4_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane4_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane4_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane4_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane4_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane4_type0                      ,                                       
      scntl__sdp__lane4_num_of_types0              ,                                       
      scntl__sdp__lane5_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane5_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane5_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane5_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane5_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane5_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane5_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane5_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane5_type0                      ,                                       
      scntl__sdp__lane5_num_of_types0              ,                                       
      scntl__sdp__lane6_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane6_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane6_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane6_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane6_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane6_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane6_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane6_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane6_type0                      ,                                       
      scntl__sdp__lane6_num_of_types0              ,                                       
      scntl__sdp__lane7_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane7_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane7_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane7_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane7_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane7_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane7_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane7_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane7_type0                      ,                                       
      scntl__sdp__lane7_num_of_types0              ,                                       
      scntl__sdp__lane8_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane8_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane8_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane8_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane8_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane8_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane8_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane8_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane8_type0                      ,                                       
      scntl__sdp__lane8_num_of_types0              ,                                       
      scntl__sdp__lane9_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane9_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane9_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane9_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane9_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane9_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane9_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane9_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane9_type0                      ,                                       
      scntl__sdp__lane9_num_of_types0              ,                                       
      scntl__sdp__lane10_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane10_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane10_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane10_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane10_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane10_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane10_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane10_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane10_type0                      ,                                       
      scntl__sdp__lane10_num_of_types0              ,                                       
      scntl__sdp__lane11_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane11_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane11_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane11_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane11_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane11_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane11_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane11_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane11_type0                      ,                                       
      scntl__sdp__lane11_num_of_types0              ,                                       
      scntl__sdp__lane12_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane12_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane12_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane12_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane12_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane12_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane12_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane12_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane12_type0                      ,                                       
      scntl__sdp__lane12_num_of_types0              ,                                       
      scntl__sdp__lane13_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane13_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane13_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane13_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane13_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane13_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane13_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane13_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane13_type0                      ,                                       
      scntl__sdp__lane13_num_of_types0              ,                                       
      scntl__sdp__lane14_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane14_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane14_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane14_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane14_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane14_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane14_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane14_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane14_type0                      ,                                       
      scntl__sdp__lane14_num_of_types0              ,                                       
      scntl__sdp__lane15_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane15_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane15_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane15_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane15_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane15_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane15_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane15_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane15_type0                      ,                                       
      scntl__sdp__lane15_num_of_types0              ,                                       
      scntl__sdp__lane16_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane16_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane16_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane16_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane16_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane16_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane16_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane16_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane16_type0                      ,                                       
      scntl__sdp__lane16_num_of_types0              ,                                       
      scntl__sdp__lane17_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane17_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane17_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane17_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane17_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane17_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane17_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane17_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane17_type0                      ,                                       
      scntl__sdp__lane17_num_of_types0              ,                                       
      scntl__sdp__lane18_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane18_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane18_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane18_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane18_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane18_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane18_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane18_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane18_type0                      ,                                       
      scntl__sdp__lane18_num_of_types0              ,                                       
      scntl__sdp__lane19_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane19_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane19_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane19_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane19_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane19_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane19_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane19_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane19_type0                      ,                                       
      scntl__sdp__lane19_num_of_types0              ,                                       
      scntl__sdp__lane20_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane20_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane20_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane20_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane20_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane20_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane20_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane20_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane20_type0                      ,                                       
      scntl__sdp__lane20_num_of_types0              ,                                       
      scntl__sdp__lane21_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane21_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane21_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane21_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane21_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane21_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane21_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane21_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane21_type0                      ,                                       
      scntl__sdp__lane21_num_of_types0              ,                                       
      scntl__sdp__lane22_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane22_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane22_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane22_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane22_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane22_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane22_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane22_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane22_type0                      ,                                       
      scntl__sdp__lane22_num_of_types0              ,                                       
      scntl__sdp__lane23_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane23_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane23_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane23_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane23_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane23_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane23_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane23_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane23_type0                      ,                                       
      scntl__sdp__lane23_num_of_types0              ,                                       
      scntl__sdp__lane24_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane24_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane24_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane24_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane24_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane24_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane24_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane24_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane24_type0                      ,                                       
      scntl__sdp__lane24_num_of_types0              ,                                       
      scntl__sdp__lane25_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane25_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane25_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane25_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane25_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane25_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane25_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane25_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane25_type0                      ,                                       
      scntl__sdp__lane25_num_of_types0              ,                                       
      scntl__sdp__lane26_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane26_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane26_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane26_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane26_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane26_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane26_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane26_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane26_type0                      ,                                       
      scntl__sdp__lane26_num_of_types0              ,                                       
      scntl__sdp__lane27_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane27_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane27_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane27_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane27_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane27_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane27_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane27_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane27_type0                      ,                                       
      scntl__sdp__lane27_num_of_types0              ,                                       
      scntl__sdp__lane28_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane28_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane28_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane28_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane28_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane28_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane28_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane28_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane28_type0                      ,                                       
      scntl__sdp__lane28_num_of_types0              ,                                       
      scntl__sdp__lane29_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane29_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane29_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane29_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane29_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane29_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane29_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane29_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane29_type0                      ,                                       
      scntl__sdp__lane29_num_of_types0              ,                                       
      scntl__sdp__lane30_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane30_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane30_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane30_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane30_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane30_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane30_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane30_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane30_type0                      ,                                       
      scntl__sdp__lane30_num_of_types0              ,                                       
      scntl__sdp__lane31_strm0_read_enable          ,  // enable the stream read mode       
      scntl__sdp__lane31_strm0_write_enable         ,  // enable the stream write mode      
      sdp__scntl__lane31_strm0_read_ready           ,  // stream read mode ready            
      sdp__scntl__lane31_strm0_write_ready          ,  // stream write mode ready           
      sdp__scntl__lane31_strm0_read_complete        ,  // stream read mode complete         
      sdp__scntl__lane31_strm0_write_complete       ,  // stream write mode complete        
      scntl__sdp__lane31_strm0_read_start_address   ,  // streaming op arg0               
      scntl__sdp__lane31_strm0_write_start_address  ,  // streaming op result start address 
      scntl__sdp__lane31_type0                      ,                                       
      scntl__sdp__lane31_num_of_types0              ,                                       

      scntl__sdp__lane0_strm0_stOp_source          ,                                       
      scntl__sdp__lane0_strm0_stOp_destination     ,                                       
      scntl__sdp__lane0_strm0_stOp_enable          ,                                       
      sdp__scntl__lane0_strm0_stOp_ready           ,                                       
      sdp__scntl__lane0_strm0_stOp_complete        ,                                       
      scntl__sdp__lane0_strm1_stOp_source          ,                                       
      scntl__sdp__lane0_strm1_stOp_destination     ,                                       
      scntl__sdp__lane0_strm1_stOp_enable          ,                                       
      sdp__scntl__lane0_strm1_stOp_ready           ,                                       
      sdp__scntl__lane0_strm1_stOp_complete        ,                                       
      scntl__sdp__lane1_strm0_stOp_source          ,                                       
      scntl__sdp__lane1_strm0_stOp_destination     ,                                       
      scntl__sdp__lane1_strm0_stOp_enable          ,                                       
      sdp__scntl__lane1_strm0_stOp_ready           ,                                       
      sdp__scntl__lane1_strm0_stOp_complete        ,                                       
      scntl__sdp__lane1_strm1_stOp_source          ,                                       
      scntl__sdp__lane1_strm1_stOp_destination     ,                                       
      scntl__sdp__lane1_strm1_stOp_enable          ,                                       
      sdp__scntl__lane1_strm1_stOp_ready           ,                                       
      sdp__scntl__lane1_strm1_stOp_complete        ,                                       
      scntl__sdp__lane2_strm0_stOp_source          ,                                       
      scntl__sdp__lane2_strm0_stOp_destination     ,                                       
      scntl__sdp__lane2_strm0_stOp_enable          ,                                       
      sdp__scntl__lane2_strm0_stOp_ready           ,                                       
      sdp__scntl__lane2_strm0_stOp_complete        ,                                       
      scntl__sdp__lane2_strm1_stOp_source          ,                                       
      scntl__sdp__lane2_strm1_stOp_destination     ,                                       
      scntl__sdp__lane2_strm1_stOp_enable          ,                                       
      sdp__scntl__lane2_strm1_stOp_ready           ,                                       
      sdp__scntl__lane2_strm1_stOp_complete        ,                                       
      scntl__sdp__lane3_strm0_stOp_source          ,                                       
      scntl__sdp__lane3_strm0_stOp_destination     ,                                       
      scntl__sdp__lane3_strm0_stOp_enable          ,                                       
      sdp__scntl__lane3_strm0_stOp_ready           ,                                       
      sdp__scntl__lane3_strm0_stOp_complete        ,                                       
      scntl__sdp__lane3_strm1_stOp_source          ,                                       
      scntl__sdp__lane3_strm1_stOp_destination     ,                                       
      scntl__sdp__lane3_strm1_stOp_enable          ,                                       
      sdp__scntl__lane3_strm1_stOp_ready           ,                                       
      sdp__scntl__lane3_strm1_stOp_complete        ,                                       
      scntl__sdp__lane4_strm0_stOp_source          ,                                       
      scntl__sdp__lane4_strm0_stOp_destination     ,                                       
      scntl__sdp__lane4_strm0_stOp_enable          ,                                       
      sdp__scntl__lane4_strm0_stOp_ready           ,                                       
      sdp__scntl__lane4_strm0_stOp_complete        ,                                       
      scntl__sdp__lane4_strm1_stOp_source          ,                                       
      scntl__sdp__lane4_strm1_stOp_destination     ,                                       
      scntl__sdp__lane4_strm1_stOp_enable          ,                                       
      sdp__scntl__lane4_strm1_stOp_ready           ,                                       
      sdp__scntl__lane4_strm1_stOp_complete        ,                                       
      scntl__sdp__lane5_strm0_stOp_source          ,                                       
      scntl__sdp__lane5_strm0_stOp_destination     ,                                       
      scntl__sdp__lane5_strm0_stOp_enable          ,                                       
      sdp__scntl__lane5_strm0_stOp_ready           ,                                       
      sdp__scntl__lane5_strm0_stOp_complete        ,                                       
      scntl__sdp__lane5_strm1_stOp_source          ,                                       
      scntl__sdp__lane5_strm1_stOp_destination     ,                                       
      scntl__sdp__lane5_strm1_stOp_enable          ,                                       
      sdp__scntl__lane5_strm1_stOp_ready           ,                                       
      sdp__scntl__lane5_strm1_stOp_complete        ,                                       
      scntl__sdp__lane6_strm0_stOp_source          ,                                       
      scntl__sdp__lane6_strm0_stOp_destination     ,                                       
      scntl__sdp__lane6_strm0_stOp_enable          ,                                       
      sdp__scntl__lane6_strm0_stOp_ready           ,                                       
      sdp__scntl__lane6_strm0_stOp_complete        ,                                       
      scntl__sdp__lane6_strm1_stOp_source          ,                                       
      scntl__sdp__lane6_strm1_stOp_destination     ,                                       
      scntl__sdp__lane6_strm1_stOp_enable          ,                                       
      sdp__scntl__lane6_strm1_stOp_ready           ,                                       
      sdp__scntl__lane6_strm1_stOp_complete        ,                                       
      scntl__sdp__lane7_strm0_stOp_source          ,                                       
      scntl__sdp__lane7_strm0_stOp_destination     ,                                       
      scntl__sdp__lane7_strm0_stOp_enable          ,                                       
      sdp__scntl__lane7_strm0_stOp_ready           ,                                       
      sdp__scntl__lane7_strm0_stOp_complete        ,                                       
      scntl__sdp__lane7_strm1_stOp_source          ,                                       
      scntl__sdp__lane7_strm1_stOp_destination     ,                                       
      scntl__sdp__lane7_strm1_stOp_enable          ,                                       
      sdp__scntl__lane7_strm1_stOp_ready           ,                                       
      sdp__scntl__lane7_strm1_stOp_complete        ,                                       
      scntl__sdp__lane8_strm0_stOp_source          ,                                       
      scntl__sdp__lane8_strm0_stOp_destination     ,                                       
      scntl__sdp__lane8_strm0_stOp_enable          ,                                       
      sdp__scntl__lane8_strm0_stOp_ready           ,                                       
      sdp__scntl__lane8_strm0_stOp_complete        ,                                       
      scntl__sdp__lane8_strm1_stOp_source          ,                                       
      scntl__sdp__lane8_strm1_stOp_destination     ,                                       
      scntl__sdp__lane8_strm1_stOp_enable          ,                                       
      sdp__scntl__lane8_strm1_stOp_ready           ,                                       
      sdp__scntl__lane8_strm1_stOp_complete        ,                                       
      scntl__sdp__lane9_strm0_stOp_source          ,                                       
      scntl__sdp__lane9_strm0_stOp_destination     ,                                       
      scntl__sdp__lane9_strm0_stOp_enable          ,                                       
      sdp__scntl__lane9_strm0_stOp_ready           ,                                       
      sdp__scntl__lane9_strm0_stOp_complete        ,                                       
      scntl__sdp__lane9_strm1_stOp_source          ,                                       
      scntl__sdp__lane9_strm1_stOp_destination     ,                                       
      scntl__sdp__lane9_strm1_stOp_enable          ,                                       
      sdp__scntl__lane9_strm1_stOp_ready           ,                                       
      sdp__scntl__lane9_strm1_stOp_complete        ,                                       
      scntl__sdp__lane10_strm0_stOp_source          ,                                       
      scntl__sdp__lane10_strm0_stOp_destination     ,                                       
      scntl__sdp__lane10_strm0_stOp_enable          ,                                       
      sdp__scntl__lane10_strm0_stOp_ready           ,                                       
      sdp__scntl__lane10_strm0_stOp_complete        ,                                       
      scntl__sdp__lane10_strm1_stOp_source          ,                                       
      scntl__sdp__lane10_strm1_stOp_destination     ,                                       
      scntl__sdp__lane10_strm1_stOp_enable          ,                                       
      sdp__scntl__lane10_strm1_stOp_ready           ,                                       
      sdp__scntl__lane10_strm1_stOp_complete        ,                                       
      scntl__sdp__lane11_strm0_stOp_source          ,                                       
      scntl__sdp__lane11_strm0_stOp_destination     ,                                       
      scntl__sdp__lane11_strm0_stOp_enable          ,                                       
      sdp__scntl__lane11_strm0_stOp_ready           ,                                       
      sdp__scntl__lane11_strm0_stOp_complete        ,                                       
      scntl__sdp__lane11_strm1_stOp_source          ,                                       
      scntl__sdp__lane11_strm1_stOp_destination     ,                                       
      scntl__sdp__lane11_strm1_stOp_enable          ,                                       
      sdp__scntl__lane11_strm1_stOp_ready           ,                                       
      sdp__scntl__lane11_strm1_stOp_complete        ,                                       
      scntl__sdp__lane12_strm0_stOp_source          ,                                       
      scntl__sdp__lane12_strm0_stOp_destination     ,                                       
      scntl__sdp__lane12_strm0_stOp_enable          ,                                       
      sdp__scntl__lane12_strm0_stOp_ready           ,                                       
      sdp__scntl__lane12_strm0_stOp_complete        ,                                       
      scntl__sdp__lane12_strm1_stOp_source          ,                                       
      scntl__sdp__lane12_strm1_stOp_destination     ,                                       
      scntl__sdp__lane12_strm1_stOp_enable          ,                                       
      sdp__scntl__lane12_strm1_stOp_ready           ,                                       
      sdp__scntl__lane12_strm1_stOp_complete        ,                                       
      scntl__sdp__lane13_strm0_stOp_source          ,                                       
      scntl__sdp__lane13_strm0_stOp_destination     ,                                       
      scntl__sdp__lane13_strm0_stOp_enable          ,                                       
      sdp__scntl__lane13_strm0_stOp_ready           ,                                       
      sdp__scntl__lane13_strm0_stOp_complete        ,                                       
      scntl__sdp__lane13_strm1_stOp_source          ,                                       
      scntl__sdp__lane13_strm1_stOp_destination     ,                                       
      scntl__sdp__lane13_strm1_stOp_enable          ,                                       
      sdp__scntl__lane13_strm1_stOp_ready           ,                                       
      sdp__scntl__lane13_strm1_stOp_complete        ,                                       
      scntl__sdp__lane14_strm0_stOp_source          ,                                       
      scntl__sdp__lane14_strm0_stOp_destination     ,                                       
      scntl__sdp__lane14_strm0_stOp_enable          ,                                       
      sdp__scntl__lane14_strm0_stOp_ready           ,                                       
      sdp__scntl__lane14_strm0_stOp_complete        ,                                       
      scntl__sdp__lane14_strm1_stOp_source          ,                                       
      scntl__sdp__lane14_strm1_stOp_destination     ,                                       
      scntl__sdp__lane14_strm1_stOp_enable          ,                                       
      sdp__scntl__lane14_strm1_stOp_ready           ,                                       
      sdp__scntl__lane14_strm1_stOp_complete        ,                                       
      scntl__sdp__lane15_strm0_stOp_source          ,                                       
      scntl__sdp__lane15_strm0_stOp_destination     ,                                       
      scntl__sdp__lane15_strm0_stOp_enable          ,                                       
      sdp__scntl__lane15_strm0_stOp_ready           ,                                       
      sdp__scntl__lane15_strm0_stOp_complete        ,                                       
      scntl__sdp__lane15_strm1_stOp_source          ,                                       
      scntl__sdp__lane15_strm1_stOp_destination     ,                                       
      scntl__sdp__lane15_strm1_stOp_enable          ,                                       
      sdp__scntl__lane15_strm1_stOp_ready           ,                                       
      sdp__scntl__lane15_strm1_stOp_complete        ,                                       
      scntl__sdp__lane16_strm0_stOp_source          ,                                       
      scntl__sdp__lane16_strm0_stOp_destination     ,                                       
      scntl__sdp__lane16_strm0_stOp_enable          ,                                       
      sdp__scntl__lane16_strm0_stOp_ready           ,                                       
      sdp__scntl__lane16_strm0_stOp_complete        ,                                       
      scntl__sdp__lane16_strm1_stOp_source          ,                                       
      scntl__sdp__lane16_strm1_stOp_destination     ,                                       
      scntl__sdp__lane16_strm1_stOp_enable          ,                                       
      sdp__scntl__lane16_strm1_stOp_ready           ,                                       
      sdp__scntl__lane16_strm1_stOp_complete        ,                                       
      scntl__sdp__lane17_strm0_stOp_source          ,                                       
      scntl__sdp__lane17_strm0_stOp_destination     ,                                       
      scntl__sdp__lane17_strm0_stOp_enable          ,                                       
      sdp__scntl__lane17_strm0_stOp_ready           ,                                       
      sdp__scntl__lane17_strm0_stOp_complete        ,                                       
      scntl__sdp__lane17_strm1_stOp_source          ,                                       
      scntl__sdp__lane17_strm1_stOp_destination     ,                                       
      scntl__sdp__lane17_strm1_stOp_enable          ,                                       
      sdp__scntl__lane17_strm1_stOp_ready           ,                                       
      sdp__scntl__lane17_strm1_stOp_complete        ,                                       
      scntl__sdp__lane18_strm0_stOp_source          ,                                       
      scntl__sdp__lane18_strm0_stOp_destination     ,                                       
      scntl__sdp__lane18_strm0_stOp_enable          ,                                       
      sdp__scntl__lane18_strm0_stOp_ready           ,                                       
      sdp__scntl__lane18_strm0_stOp_complete        ,                                       
      scntl__sdp__lane18_strm1_stOp_source          ,                                       
      scntl__sdp__lane18_strm1_stOp_destination     ,                                       
      scntl__sdp__lane18_strm1_stOp_enable          ,                                       
      sdp__scntl__lane18_strm1_stOp_ready           ,                                       
      sdp__scntl__lane18_strm1_stOp_complete        ,                                       
      scntl__sdp__lane19_strm0_stOp_source          ,                                       
      scntl__sdp__lane19_strm0_stOp_destination     ,                                       
      scntl__sdp__lane19_strm0_stOp_enable          ,                                       
      sdp__scntl__lane19_strm0_stOp_ready           ,                                       
      sdp__scntl__lane19_strm0_stOp_complete        ,                                       
      scntl__sdp__lane19_strm1_stOp_source          ,                                       
      scntl__sdp__lane19_strm1_stOp_destination     ,                                       
      scntl__sdp__lane19_strm1_stOp_enable          ,                                       
      sdp__scntl__lane19_strm1_stOp_ready           ,                                       
      sdp__scntl__lane19_strm1_stOp_complete        ,                                       
      scntl__sdp__lane20_strm0_stOp_source          ,                                       
      scntl__sdp__lane20_strm0_stOp_destination     ,                                       
      scntl__sdp__lane20_strm0_stOp_enable          ,                                       
      sdp__scntl__lane20_strm0_stOp_ready           ,                                       
      sdp__scntl__lane20_strm0_stOp_complete        ,                                       
      scntl__sdp__lane20_strm1_stOp_source          ,                                       
      scntl__sdp__lane20_strm1_stOp_destination     ,                                       
      scntl__sdp__lane20_strm1_stOp_enable          ,                                       
      sdp__scntl__lane20_strm1_stOp_ready           ,                                       
      sdp__scntl__lane20_strm1_stOp_complete        ,                                       
      scntl__sdp__lane21_strm0_stOp_source          ,                                       
      scntl__sdp__lane21_strm0_stOp_destination     ,                                       
      scntl__sdp__lane21_strm0_stOp_enable          ,                                       
      sdp__scntl__lane21_strm0_stOp_ready           ,                                       
      sdp__scntl__lane21_strm0_stOp_complete        ,                                       
      scntl__sdp__lane21_strm1_stOp_source          ,                                       
      scntl__sdp__lane21_strm1_stOp_destination     ,                                       
      scntl__sdp__lane21_strm1_stOp_enable          ,                                       
      sdp__scntl__lane21_strm1_stOp_ready           ,                                       
      sdp__scntl__lane21_strm1_stOp_complete        ,                                       
      scntl__sdp__lane22_strm0_stOp_source          ,                                       
      scntl__sdp__lane22_strm0_stOp_destination     ,                                       
      scntl__sdp__lane22_strm0_stOp_enable          ,                                       
      sdp__scntl__lane22_strm0_stOp_ready           ,                                       
      sdp__scntl__lane22_strm0_stOp_complete        ,                                       
      scntl__sdp__lane22_strm1_stOp_source          ,                                       
      scntl__sdp__lane22_strm1_stOp_destination     ,                                       
      scntl__sdp__lane22_strm1_stOp_enable          ,                                       
      sdp__scntl__lane22_strm1_stOp_ready           ,                                       
      sdp__scntl__lane22_strm1_stOp_complete        ,                                       
      scntl__sdp__lane23_strm0_stOp_source          ,                                       
      scntl__sdp__lane23_strm0_stOp_destination     ,                                       
      scntl__sdp__lane23_strm0_stOp_enable          ,                                       
      sdp__scntl__lane23_strm0_stOp_ready           ,                                       
      sdp__scntl__lane23_strm0_stOp_complete        ,                                       
      scntl__sdp__lane23_strm1_stOp_source          ,                                       
      scntl__sdp__lane23_strm1_stOp_destination     ,                                       
      scntl__sdp__lane23_strm1_stOp_enable          ,                                       
      sdp__scntl__lane23_strm1_stOp_ready           ,                                       
      sdp__scntl__lane23_strm1_stOp_complete        ,                                       
      scntl__sdp__lane24_strm0_stOp_source          ,                                       
      scntl__sdp__lane24_strm0_stOp_destination     ,                                       
      scntl__sdp__lane24_strm0_stOp_enable          ,                                       
      sdp__scntl__lane24_strm0_stOp_ready           ,                                       
      sdp__scntl__lane24_strm0_stOp_complete        ,                                       
      scntl__sdp__lane24_strm1_stOp_source          ,                                       
      scntl__sdp__lane24_strm1_stOp_destination     ,                                       
      scntl__sdp__lane24_strm1_stOp_enable          ,                                       
      sdp__scntl__lane24_strm1_stOp_ready           ,                                       
      sdp__scntl__lane24_strm1_stOp_complete        ,                                       
      scntl__sdp__lane25_strm0_stOp_source          ,                                       
      scntl__sdp__lane25_strm0_stOp_destination     ,                                       
      scntl__sdp__lane25_strm0_stOp_enable          ,                                       
      sdp__scntl__lane25_strm0_stOp_ready           ,                                       
      sdp__scntl__lane25_strm0_stOp_complete        ,                                       
      scntl__sdp__lane25_strm1_stOp_source          ,                                       
      scntl__sdp__lane25_strm1_stOp_destination     ,                                       
      scntl__sdp__lane25_strm1_stOp_enable          ,                                       
      sdp__scntl__lane25_strm1_stOp_ready           ,                                       
      sdp__scntl__lane25_strm1_stOp_complete        ,                                       
      scntl__sdp__lane26_strm0_stOp_source          ,                                       
      scntl__sdp__lane26_strm0_stOp_destination     ,                                       
      scntl__sdp__lane26_strm0_stOp_enable          ,                                       
      sdp__scntl__lane26_strm0_stOp_ready           ,                                       
      sdp__scntl__lane26_strm0_stOp_complete        ,                                       
      scntl__sdp__lane26_strm1_stOp_source          ,                                       
      scntl__sdp__lane26_strm1_stOp_destination     ,                                       
      scntl__sdp__lane26_strm1_stOp_enable          ,                                       
      sdp__scntl__lane26_strm1_stOp_ready           ,                                       
      sdp__scntl__lane26_strm1_stOp_complete        ,                                       
      scntl__sdp__lane27_strm0_stOp_source          ,                                       
      scntl__sdp__lane27_strm0_stOp_destination     ,                                       
      scntl__sdp__lane27_strm0_stOp_enable          ,                                       
      sdp__scntl__lane27_strm0_stOp_ready           ,                                       
      sdp__scntl__lane27_strm0_stOp_complete        ,                                       
      scntl__sdp__lane27_strm1_stOp_source          ,                                       
      scntl__sdp__lane27_strm1_stOp_destination     ,                                       
      scntl__sdp__lane27_strm1_stOp_enable          ,                                       
      sdp__scntl__lane27_strm1_stOp_ready           ,                                       
      sdp__scntl__lane27_strm1_stOp_complete        ,                                       
      scntl__sdp__lane28_strm0_stOp_source          ,                                       
      scntl__sdp__lane28_strm0_stOp_destination     ,                                       
      scntl__sdp__lane28_strm0_stOp_enable          ,                                       
      sdp__scntl__lane28_strm0_stOp_ready           ,                                       
      sdp__scntl__lane28_strm0_stOp_complete        ,                                       
      scntl__sdp__lane28_strm1_stOp_source          ,                                       
      scntl__sdp__lane28_strm1_stOp_destination     ,                                       
      scntl__sdp__lane28_strm1_stOp_enable          ,                                       
      sdp__scntl__lane28_strm1_stOp_ready           ,                                       
      sdp__scntl__lane28_strm1_stOp_complete        ,                                       
      scntl__sdp__lane29_strm0_stOp_source          ,                                       
      scntl__sdp__lane29_strm0_stOp_destination     ,                                       
      scntl__sdp__lane29_strm0_stOp_enable          ,                                       
      sdp__scntl__lane29_strm0_stOp_ready           ,                                       
      sdp__scntl__lane29_strm0_stOp_complete        ,                                       
      scntl__sdp__lane29_strm1_stOp_source          ,                                       
      scntl__sdp__lane29_strm1_stOp_destination     ,                                       
      scntl__sdp__lane29_strm1_stOp_enable          ,                                       
      sdp__scntl__lane29_strm1_stOp_ready           ,                                       
      sdp__scntl__lane29_strm1_stOp_complete        ,                                       
      scntl__sdp__lane30_strm0_stOp_source          ,                                       
      scntl__sdp__lane30_strm0_stOp_destination     ,                                       
      scntl__sdp__lane30_strm0_stOp_enable          ,                                       
      sdp__scntl__lane30_strm0_stOp_ready           ,                                       
      sdp__scntl__lane30_strm0_stOp_complete        ,                                       
      scntl__sdp__lane30_strm1_stOp_source          ,                                       
      scntl__sdp__lane30_strm1_stOp_destination     ,                                       
      scntl__sdp__lane30_strm1_stOp_enable          ,                                       
      sdp__scntl__lane30_strm1_stOp_ready           ,                                       
      sdp__scntl__lane30_strm1_stOp_complete        ,                                       
      scntl__sdp__lane31_strm0_stOp_source          ,                                       
      scntl__sdp__lane31_strm0_stOp_destination     ,                                       
      scntl__sdp__lane31_strm0_stOp_enable          ,                                       
      sdp__scntl__lane31_strm0_stOp_ready           ,                                       
      sdp__scntl__lane31_strm0_stOp_complete        ,                                       
      scntl__sdp__lane31_strm1_stOp_source          ,                                       
      scntl__sdp__lane31_strm1_stOp_destination     ,                                       
      scntl__sdp__lane31_strm1_stOp_enable          ,                                       
      sdp__scntl__lane31_strm1_stOp_ready           ,                                       
      sdp__scntl__lane31_strm1_stOp_complete        ,                                       
