
    // Common (Scalar) Register(s)                
            rs0                  ,
            rs1                  ,

    // Lane 0                 
            lane0_r128                  ,
            lane0_r129                  ,
            lane0_r130                  ,
            lane0_r131                  ,
            lane0_r132                  ,
            lane0_r133                  ,
            lane0_r134                  ,
            lane0_r135                  ,

    // Lane 1                 
            lane1_r128                  ,
            lane1_r129                  ,
            lane1_r130                  ,
            lane1_r131                  ,
            lane1_r132                  ,
            lane1_r133                  ,
            lane1_r134                  ,
            lane1_r135                  ,

    // Lane 2                 
            lane2_r128                  ,
            lane2_r129                  ,
            lane2_r130                  ,
            lane2_r131                  ,
            lane2_r132                  ,
            lane2_r133                  ,
            lane2_r134                  ,
            lane2_r135                  ,

    // Lane 3                 
            lane3_r128                  ,
            lane3_r129                  ,
            lane3_r130                  ,
            lane3_r131                  ,
            lane3_r132                  ,
            lane3_r133                  ,
            lane3_r134                  ,
            lane3_r135                  ,

    // Lane 4                 
            lane4_r128                  ,
            lane4_r129                  ,
            lane4_r130                  ,
            lane4_r131                  ,
            lane4_r132                  ,
            lane4_r133                  ,
            lane4_r134                  ,
            lane4_r135                  ,

    // Lane 5                 
            lane5_r128                  ,
            lane5_r129                  ,
            lane5_r130                  ,
            lane5_r131                  ,
            lane5_r132                  ,
            lane5_r133                  ,
            lane5_r134                  ,
            lane5_r135                  ,

    // Lane 6                 
            lane6_r128                  ,
            lane6_r129                  ,
            lane6_r130                  ,
            lane6_r131                  ,
            lane6_r132                  ,
            lane6_r133                  ,
            lane6_r134                  ,
            lane6_r135                  ,

    // Lane 7                 
            lane7_r128                  ,
            lane7_r129                  ,
            lane7_r130                  ,
            lane7_r131                  ,
            lane7_r132                  ,
            lane7_r133                  ,
            lane7_r134                  ,
            lane7_r135                  ,

    // Lane 8                 
            lane8_r128                  ,
            lane8_r129                  ,
            lane8_r130                  ,
            lane8_r131                  ,
            lane8_r132                  ,
            lane8_r133                  ,
            lane8_r134                  ,
            lane8_r135                  ,

    // Lane 9                 
            lane9_r128                  ,
            lane9_r129                  ,
            lane9_r130                  ,
            lane9_r131                  ,
            lane9_r132                  ,
            lane9_r133                  ,
            lane9_r134                  ,
            lane9_r135                  ,

    // Lane 10                 
            lane10_r128                  ,
            lane10_r129                  ,
            lane10_r130                  ,
            lane10_r131                  ,
            lane10_r132                  ,
            lane10_r133                  ,
            lane10_r134                  ,
            lane10_r135                  ,

    // Lane 11                 
            lane11_r128                  ,
            lane11_r129                  ,
            lane11_r130                  ,
            lane11_r131                  ,
            lane11_r132                  ,
            lane11_r133                  ,
            lane11_r134                  ,
            lane11_r135                  ,

    // Lane 12                 
            lane12_r128                  ,
            lane12_r129                  ,
            lane12_r130                  ,
            lane12_r131                  ,
            lane12_r132                  ,
            lane12_r133                  ,
            lane12_r134                  ,
            lane12_r135                  ,

    // Lane 13                 
            lane13_r128                  ,
            lane13_r129                  ,
            lane13_r130                  ,
            lane13_r131                  ,
            lane13_r132                  ,
            lane13_r133                  ,
            lane13_r134                  ,
            lane13_r135                  ,

    // Lane 14                 
            lane14_r128                  ,
            lane14_r129                  ,
            lane14_r130                  ,
            lane14_r131                  ,
            lane14_r132                  ,
            lane14_r133                  ,
            lane14_r134                  ,
            lane14_r135                  ,

    // Lane 15                 
            lane15_r128                  ,
            lane15_r129                  ,
            lane15_r130                  ,
            lane15_r131                  ,
            lane15_r132                  ,
            lane15_r133                  ,
            lane15_r134                  ,
            lane15_r135                  ,

    // Lane 16                 
            lane16_r128                  ,
            lane16_r129                  ,
            lane16_r130                  ,
            lane16_r131                  ,
            lane16_r132                  ,
            lane16_r133                  ,
            lane16_r134                  ,
            lane16_r135                  ,

    // Lane 17                 
            lane17_r128                  ,
            lane17_r129                  ,
            lane17_r130                  ,
            lane17_r131                  ,
            lane17_r132                  ,
            lane17_r133                  ,
            lane17_r134                  ,
            lane17_r135                  ,

    // Lane 18                 
            lane18_r128                  ,
            lane18_r129                  ,
            lane18_r130                  ,
            lane18_r131                  ,
            lane18_r132                  ,
            lane18_r133                  ,
            lane18_r134                  ,
            lane18_r135                  ,

    // Lane 19                 
            lane19_r128                  ,
            lane19_r129                  ,
            lane19_r130                  ,
            lane19_r131                  ,
            lane19_r132                  ,
            lane19_r133                  ,
            lane19_r134                  ,
            lane19_r135                  ,

    // Lane 20                 
            lane20_r128                  ,
            lane20_r129                  ,
            lane20_r130                  ,
            lane20_r131                  ,
            lane20_r132                  ,
            lane20_r133                  ,
            lane20_r134                  ,
            lane20_r135                  ,

    // Lane 21                 
            lane21_r128                  ,
            lane21_r129                  ,
            lane21_r130                  ,
            lane21_r131                  ,
            lane21_r132                  ,
            lane21_r133                  ,
            lane21_r134                  ,
            lane21_r135                  ,

    // Lane 22                 
            lane22_r128                  ,
            lane22_r129                  ,
            lane22_r130                  ,
            lane22_r131                  ,
            lane22_r132                  ,
            lane22_r133                  ,
            lane22_r134                  ,
            lane22_r135                  ,

    // Lane 23                 
            lane23_r128                  ,
            lane23_r129                  ,
            lane23_r130                  ,
            lane23_r131                  ,
            lane23_r132                  ,
            lane23_r133                  ,
            lane23_r134                  ,
            lane23_r135                  ,

    // Lane 24                 
            lane24_r128                  ,
            lane24_r129                  ,
            lane24_r130                  ,
            lane24_r131                  ,
            lane24_r132                  ,
            lane24_r133                  ,
            lane24_r134                  ,
            lane24_r135                  ,

    // Lane 25                 
            lane25_r128                  ,
            lane25_r129                  ,
            lane25_r130                  ,
            lane25_r131                  ,
            lane25_r132                  ,
            lane25_r133                  ,
            lane25_r134                  ,
            lane25_r135                  ,

    // Lane 26                 
            lane26_r128                  ,
            lane26_r129                  ,
            lane26_r130                  ,
            lane26_r131                  ,
            lane26_r132                  ,
            lane26_r133                  ,
            lane26_r134                  ,
            lane26_r135                  ,

    // Lane 27                 
            lane27_r128                  ,
            lane27_r129                  ,
            lane27_r130                  ,
            lane27_r131                  ,
            lane27_r132                  ,
            lane27_r133                  ,
            lane27_r134                  ,
            lane27_r135                  ,

    // Lane 28                 
            lane28_r128                  ,
            lane28_r129                  ,
            lane28_r130                  ,
            lane28_r131                  ,
            lane28_r132                  ,
            lane28_r133                  ,
            lane28_r134                  ,
            lane28_r135                  ,

    // Lane 29                 
            lane29_r128                  ,
            lane29_r129                  ,
            lane29_r130                  ,
            lane29_r131                  ,
            lane29_r132                  ,
            lane29_r133                  ,
            lane29_r134                  ,
            lane29_r135                  ,

    // Lane 30                 
            lane30_r128                  ,
            lane30_r129                  ,
            lane30_r130                  ,
            lane30_r131                  ,
            lane30_r132                  ,
            lane30_r133                  ,
            lane30_r134                  ,
            lane30_r135                  ,

    // Lane 31                 
            lane31_r128                  ,
            lane31_r129                  ,
            lane31_r130                  ,
            lane31_r131                  ,
            lane31_r132                  ,
            lane31_r133                  ,
            lane31_r134                  ,
            lane31_r135                  ,
