
            begin
              @(final_operation[0][0]) ;
              //$display("@%0t LEE: Received final operation event for 0,0\n", $time);
            end
            begin
              @(final_operation[0][1]) ;
              //$display("@%0t LEE: Received final operation event for 0,1\n", $time);
            end
            begin
              @(final_operation[0][2]) ;
              //$display("@%0t LEE: Received final operation event for 0,2\n", $time);
            end
            begin
              @(final_operation[0][3]) ;
              //$display("@%0t LEE: Received final operation event for 0,3\n", $time);
            end
            begin
              @(final_operation[0][4]) ;
              //$display("@%0t LEE: Received final operation event for 0,4\n", $time);
            end
            begin
              @(final_operation[0][5]) ;
              //$display("@%0t LEE: Received final operation event for 0,5\n", $time);
            end
            begin
              @(final_operation[0][6]) ;
              //$display("@%0t LEE: Received final operation event for 0,6\n", $time);
            end
            begin
              @(final_operation[0][7]) ;
              //$display("@%0t LEE: Received final operation event for 0,7\n", $time);
            end
            begin
              @(final_operation[0][8]) ;
              //$display("@%0t LEE: Received final operation event for 0,8\n", $time);
            end
            begin
              @(final_operation[0][9]) ;
              //$display("@%0t LEE: Received final operation event for 0,9\n", $time);
            end
            begin
              @(final_operation[0][10]) ;
              //$display("@%0t LEE: Received final operation event for 0,10\n", $time);
            end
            begin
              @(final_operation[0][11]) ;
              //$display("@%0t LEE: Received final operation event for 0,11\n", $time);
            end
            begin
              @(final_operation[0][12]) ;
              //$display("@%0t LEE: Received final operation event for 0,12\n", $time);
            end
            begin
              @(final_operation[0][13]) ;
              //$display("@%0t LEE: Received final operation event for 0,13\n", $time);
            end
            begin
              @(final_operation[0][14]) ;
              //$display("@%0t LEE: Received final operation event for 0,14\n", $time);
            end
            begin
              @(final_operation[0][15]) ;
              //$display("@%0t LEE: Received final operation event for 0,15\n", $time);
            end
            begin
              @(final_operation[0][16]) ;
              //$display("@%0t LEE: Received final operation event for 0,16\n", $time);
            end
            begin
              @(final_operation[0][17]) ;
              //$display("@%0t LEE: Received final operation event for 0,17\n", $time);
            end
            begin
              @(final_operation[0][18]) ;
              //$display("@%0t LEE: Received final operation event for 0,18\n", $time);
            end
            begin
              @(final_operation[0][19]) ;
              //$display("@%0t LEE: Received final operation event for 0,19\n", $time);
            end
            begin
              @(final_operation[0][20]) ;
              //$display("@%0t LEE: Received final operation event for 0,20\n", $time);
            end
            begin
              @(final_operation[0][21]) ;
              //$display("@%0t LEE: Received final operation event for 0,21\n", $time);
            end
            begin
              @(final_operation[0][22]) ;
              //$display("@%0t LEE: Received final operation event for 0,22\n", $time);
            end
            begin
              @(final_operation[0][23]) ;
              //$display("@%0t LEE: Received final operation event for 0,23\n", $time);
            end
            begin
              @(final_operation[0][24]) ;
              //$display("@%0t LEE: Received final operation event for 0,24\n", $time);
            end
            begin
              @(final_operation[0][25]) ;
              //$display("@%0t LEE: Received final operation event for 0,25\n", $time);
            end
            begin
              @(final_operation[0][26]) ;
              //$display("@%0t LEE: Received final operation event for 0,26\n", $time);
            end
            begin
              @(final_operation[0][27]) ;
              //$display("@%0t LEE: Received final operation event for 0,27\n", $time);
            end
            begin
              @(final_operation[0][28]) ;
              //$display("@%0t LEE: Received final operation event for 0,28\n", $time);
            end
            begin
              @(final_operation[0][29]) ;
              //$display("@%0t LEE: Received final operation event for 0,29\n", $time);
            end
            begin
              @(final_operation[0][30]) ;
              //$display("@%0t LEE: Received final operation event for 0,30\n", $time);
            end
            begin
              @(final_operation[0][31]) ;
              //$display("@%0t LEE: Received final operation event for 0,31\n", $time);
            end

            begin
              @(final_operation[1][0]) ;
              //$display("@%0t LEE: Received final operation event for 1,0\n", $time);
            end
            begin
              @(final_operation[1][1]) ;
              //$display("@%0t LEE: Received final operation event for 1,1\n", $time);
            end
            begin
              @(final_operation[1][2]) ;
              //$display("@%0t LEE: Received final operation event for 1,2\n", $time);
            end
            begin
              @(final_operation[1][3]) ;
              //$display("@%0t LEE: Received final operation event for 1,3\n", $time);
            end
            begin
              @(final_operation[1][4]) ;
              //$display("@%0t LEE: Received final operation event for 1,4\n", $time);
            end
            begin
              @(final_operation[1][5]) ;
              //$display("@%0t LEE: Received final operation event for 1,5\n", $time);
            end
            begin
              @(final_operation[1][6]) ;
              //$display("@%0t LEE: Received final operation event for 1,6\n", $time);
            end
            begin
              @(final_operation[1][7]) ;
              //$display("@%0t LEE: Received final operation event for 1,7\n", $time);
            end
            begin
              @(final_operation[1][8]) ;
              //$display("@%0t LEE: Received final operation event for 1,8\n", $time);
            end
            begin
              @(final_operation[1][9]) ;
              //$display("@%0t LEE: Received final operation event for 1,9\n", $time);
            end
            begin
              @(final_operation[1][10]) ;
              //$display("@%0t LEE: Received final operation event for 1,10\n", $time);
            end
            begin
              @(final_operation[1][11]) ;
              //$display("@%0t LEE: Received final operation event for 1,11\n", $time);
            end
            begin
              @(final_operation[1][12]) ;
              //$display("@%0t LEE: Received final operation event for 1,12\n", $time);
            end
            begin
              @(final_operation[1][13]) ;
              //$display("@%0t LEE: Received final operation event for 1,13\n", $time);
            end
            begin
              @(final_operation[1][14]) ;
              //$display("@%0t LEE: Received final operation event for 1,14\n", $time);
            end
            begin
              @(final_operation[1][15]) ;
              //$display("@%0t LEE: Received final operation event for 1,15\n", $time);
            end
            begin
              @(final_operation[1][16]) ;
              //$display("@%0t LEE: Received final operation event for 1,16\n", $time);
            end
            begin
              @(final_operation[1][17]) ;
              //$display("@%0t LEE: Received final operation event for 1,17\n", $time);
            end
            begin
              @(final_operation[1][18]) ;
              //$display("@%0t LEE: Received final operation event for 1,18\n", $time);
            end
            begin
              @(final_operation[1][19]) ;
              //$display("@%0t LEE: Received final operation event for 1,19\n", $time);
            end
            begin
              @(final_operation[1][20]) ;
              //$display("@%0t LEE: Received final operation event for 1,20\n", $time);
            end
            begin
              @(final_operation[1][21]) ;
              //$display("@%0t LEE: Received final operation event for 1,21\n", $time);
            end
            begin
              @(final_operation[1][22]) ;
              //$display("@%0t LEE: Received final operation event for 1,22\n", $time);
            end
            begin
              @(final_operation[1][23]) ;
              //$display("@%0t LEE: Received final operation event for 1,23\n", $time);
            end
            begin
              @(final_operation[1][24]) ;
              //$display("@%0t LEE: Received final operation event for 1,24\n", $time);
            end
            begin
              @(final_operation[1][25]) ;
              //$display("@%0t LEE: Received final operation event for 1,25\n", $time);
            end
            begin
              @(final_operation[1][26]) ;
              //$display("@%0t LEE: Received final operation event for 1,26\n", $time);
            end
            begin
              @(final_operation[1][27]) ;
              //$display("@%0t LEE: Received final operation event for 1,27\n", $time);
            end
            begin
              @(final_operation[1][28]) ;
              //$display("@%0t LEE: Received final operation event for 1,28\n", $time);
            end
            begin
              @(final_operation[1][29]) ;
              //$display("@%0t LEE: Received final operation event for 1,29\n", $time);
            end
            begin
              @(final_operation[1][30]) ;
              //$display("@%0t LEE: Received final operation event for 1,30\n", $time);
            end
            begin
              @(final_operation[1][31]) ;
              //$display("@%0t LEE: Received final operation event for 1,31\n", $time);
            end

            begin
              @(final_operation[2][0]) ;
              //$display("@%0t LEE: Received final operation event for 2,0\n", $time);
            end
            begin
              @(final_operation[2][1]) ;
              //$display("@%0t LEE: Received final operation event for 2,1\n", $time);
            end
            begin
              @(final_operation[2][2]) ;
              //$display("@%0t LEE: Received final operation event for 2,2\n", $time);
            end
            begin
              @(final_operation[2][3]) ;
              //$display("@%0t LEE: Received final operation event for 2,3\n", $time);
            end
            begin
              @(final_operation[2][4]) ;
              //$display("@%0t LEE: Received final operation event for 2,4\n", $time);
            end
            begin
              @(final_operation[2][5]) ;
              //$display("@%0t LEE: Received final operation event for 2,5\n", $time);
            end
            begin
              @(final_operation[2][6]) ;
              //$display("@%0t LEE: Received final operation event for 2,6\n", $time);
            end
            begin
              @(final_operation[2][7]) ;
              //$display("@%0t LEE: Received final operation event for 2,7\n", $time);
            end
            begin
              @(final_operation[2][8]) ;
              //$display("@%0t LEE: Received final operation event for 2,8\n", $time);
            end
            begin
              @(final_operation[2][9]) ;
              //$display("@%0t LEE: Received final operation event for 2,9\n", $time);
            end
            begin
              @(final_operation[2][10]) ;
              //$display("@%0t LEE: Received final operation event for 2,10\n", $time);
            end
            begin
              @(final_operation[2][11]) ;
              //$display("@%0t LEE: Received final operation event for 2,11\n", $time);
            end
            begin
              @(final_operation[2][12]) ;
              //$display("@%0t LEE: Received final operation event for 2,12\n", $time);
            end
            begin
              @(final_operation[2][13]) ;
              //$display("@%0t LEE: Received final operation event for 2,13\n", $time);
            end
            begin
              @(final_operation[2][14]) ;
              //$display("@%0t LEE: Received final operation event for 2,14\n", $time);
            end
            begin
              @(final_operation[2][15]) ;
              //$display("@%0t LEE: Received final operation event for 2,15\n", $time);
            end
            begin
              @(final_operation[2][16]) ;
              //$display("@%0t LEE: Received final operation event for 2,16\n", $time);
            end
            begin
              @(final_operation[2][17]) ;
              //$display("@%0t LEE: Received final operation event for 2,17\n", $time);
            end
            begin
              @(final_operation[2][18]) ;
              //$display("@%0t LEE: Received final operation event for 2,18\n", $time);
            end
            begin
              @(final_operation[2][19]) ;
              //$display("@%0t LEE: Received final operation event for 2,19\n", $time);
            end
            begin
              @(final_operation[2][20]) ;
              //$display("@%0t LEE: Received final operation event for 2,20\n", $time);
            end
            begin
              @(final_operation[2][21]) ;
              //$display("@%0t LEE: Received final operation event for 2,21\n", $time);
            end
            begin
              @(final_operation[2][22]) ;
              //$display("@%0t LEE: Received final operation event for 2,22\n", $time);
            end
            begin
              @(final_operation[2][23]) ;
              //$display("@%0t LEE: Received final operation event for 2,23\n", $time);
            end
            begin
              @(final_operation[2][24]) ;
              //$display("@%0t LEE: Received final operation event for 2,24\n", $time);
            end
            begin
              @(final_operation[2][25]) ;
              //$display("@%0t LEE: Received final operation event for 2,25\n", $time);
            end
            begin
              @(final_operation[2][26]) ;
              //$display("@%0t LEE: Received final operation event for 2,26\n", $time);
            end
            begin
              @(final_operation[2][27]) ;
              //$display("@%0t LEE: Received final operation event for 2,27\n", $time);
            end
            begin
              @(final_operation[2][28]) ;
              //$display("@%0t LEE: Received final operation event for 2,28\n", $time);
            end
            begin
              @(final_operation[2][29]) ;
              //$display("@%0t LEE: Received final operation event for 2,29\n", $time);
            end
            begin
              @(final_operation[2][30]) ;
              //$display("@%0t LEE: Received final operation event for 2,30\n", $time);
            end
            begin
              @(final_operation[2][31]) ;
              //$display("@%0t LEE: Received final operation event for 2,31\n", $time);
            end

            begin
              @(final_operation[3][0]) ;
              //$display("@%0t LEE: Received final operation event for 3,0\n", $time);
            end
            begin
              @(final_operation[3][1]) ;
              //$display("@%0t LEE: Received final operation event for 3,1\n", $time);
            end
            begin
              @(final_operation[3][2]) ;
              //$display("@%0t LEE: Received final operation event for 3,2\n", $time);
            end
            begin
              @(final_operation[3][3]) ;
              //$display("@%0t LEE: Received final operation event for 3,3\n", $time);
            end
            begin
              @(final_operation[3][4]) ;
              //$display("@%0t LEE: Received final operation event for 3,4\n", $time);
            end
            begin
              @(final_operation[3][5]) ;
              //$display("@%0t LEE: Received final operation event for 3,5\n", $time);
            end
            begin
              @(final_operation[3][6]) ;
              //$display("@%0t LEE: Received final operation event for 3,6\n", $time);
            end
            begin
              @(final_operation[3][7]) ;
              //$display("@%0t LEE: Received final operation event for 3,7\n", $time);
            end
            begin
              @(final_operation[3][8]) ;
              //$display("@%0t LEE: Received final operation event for 3,8\n", $time);
            end
            begin
              @(final_operation[3][9]) ;
              //$display("@%0t LEE: Received final operation event for 3,9\n", $time);
            end
            begin
              @(final_operation[3][10]) ;
              //$display("@%0t LEE: Received final operation event for 3,10\n", $time);
            end
            begin
              @(final_operation[3][11]) ;
              //$display("@%0t LEE: Received final operation event for 3,11\n", $time);
            end
            begin
              @(final_operation[3][12]) ;
              //$display("@%0t LEE: Received final operation event for 3,12\n", $time);
            end
            begin
              @(final_operation[3][13]) ;
              //$display("@%0t LEE: Received final operation event for 3,13\n", $time);
            end
            begin
              @(final_operation[3][14]) ;
              //$display("@%0t LEE: Received final operation event for 3,14\n", $time);
            end
            begin
              @(final_operation[3][15]) ;
              //$display("@%0t LEE: Received final operation event for 3,15\n", $time);
            end
            begin
              @(final_operation[3][16]) ;
              //$display("@%0t LEE: Received final operation event for 3,16\n", $time);
            end
            begin
              @(final_operation[3][17]) ;
              //$display("@%0t LEE: Received final operation event for 3,17\n", $time);
            end
            begin
              @(final_operation[3][18]) ;
              //$display("@%0t LEE: Received final operation event for 3,18\n", $time);
            end
            begin
              @(final_operation[3][19]) ;
              //$display("@%0t LEE: Received final operation event for 3,19\n", $time);
            end
            begin
              @(final_operation[3][20]) ;
              //$display("@%0t LEE: Received final operation event for 3,20\n", $time);
            end
            begin
              @(final_operation[3][21]) ;
              //$display("@%0t LEE: Received final operation event for 3,21\n", $time);
            end
            begin
              @(final_operation[3][22]) ;
              //$display("@%0t LEE: Received final operation event for 3,22\n", $time);
            end
            begin
              @(final_operation[3][23]) ;
              //$display("@%0t LEE: Received final operation event for 3,23\n", $time);
            end
            begin
              @(final_operation[3][24]) ;
              //$display("@%0t LEE: Received final operation event for 3,24\n", $time);
            end
            begin
              @(final_operation[3][25]) ;
              //$display("@%0t LEE: Received final operation event for 3,25\n", $time);
            end
            begin
              @(final_operation[3][26]) ;
              //$display("@%0t LEE: Received final operation event for 3,26\n", $time);
            end
            begin
              @(final_operation[3][27]) ;
              //$display("@%0t LEE: Received final operation event for 3,27\n", $time);
            end
            begin
              @(final_operation[3][28]) ;
              //$display("@%0t LEE: Received final operation event for 3,28\n", $time);
            end
            begin
              @(final_operation[3][29]) ;
              //$display("@%0t LEE: Received final operation event for 3,29\n", $time);
            end
            begin
              @(final_operation[3][30]) ;
              //$display("@%0t LEE: Received final operation event for 3,30\n", $time);
            end
            begin
              @(final_operation[3][31]) ;
              //$display("@%0t LEE: Received final operation event for 3,31\n", $time);
            end

            begin
              @(final_operation[4][0]) ;
              //$display("@%0t LEE: Received final operation event for 4,0\n", $time);
            end
            begin
              @(final_operation[4][1]) ;
              //$display("@%0t LEE: Received final operation event for 4,1\n", $time);
            end
            begin
              @(final_operation[4][2]) ;
              //$display("@%0t LEE: Received final operation event for 4,2\n", $time);
            end
            begin
              @(final_operation[4][3]) ;
              //$display("@%0t LEE: Received final operation event for 4,3\n", $time);
            end
            begin
              @(final_operation[4][4]) ;
              //$display("@%0t LEE: Received final operation event for 4,4\n", $time);
            end
            begin
              @(final_operation[4][5]) ;
              //$display("@%0t LEE: Received final operation event for 4,5\n", $time);
            end
            begin
              @(final_operation[4][6]) ;
              //$display("@%0t LEE: Received final operation event for 4,6\n", $time);
            end
            begin
              @(final_operation[4][7]) ;
              //$display("@%0t LEE: Received final operation event for 4,7\n", $time);
            end
            begin
              @(final_operation[4][8]) ;
              //$display("@%0t LEE: Received final operation event for 4,8\n", $time);
            end
            begin
              @(final_operation[4][9]) ;
              //$display("@%0t LEE: Received final operation event for 4,9\n", $time);
            end
            begin
              @(final_operation[4][10]) ;
              //$display("@%0t LEE: Received final operation event for 4,10\n", $time);
            end
            begin
              @(final_operation[4][11]) ;
              //$display("@%0t LEE: Received final operation event for 4,11\n", $time);
            end
            begin
              @(final_operation[4][12]) ;
              //$display("@%0t LEE: Received final operation event for 4,12\n", $time);
            end
            begin
              @(final_operation[4][13]) ;
              //$display("@%0t LEE: Received final operation event for 4,13\n", $time);
            end
            begin
              @(final_operation[4][14]) ;
              //$display("@%0t LEE: Received final operation event for 4,14\n", $time);
            end
            begin
              @(final_operation[4][15]) ;
              //$display("@%0t LEE: Received final operation event for 4,15\n", $time);
            end
            begin
              @(final_operation[4][16]) ;
              //$display("@%0t LEE: Received final operation event for 4,16\n", $time);
            end
            begin
              @(final_operation[4][17]) ;
              //$display("@%0t LEE: Received final operation event for 4,17\n", $time);
            end
            begin
              @(final_operation[4][18]) ;
              //$display("@%0t LEE: Received final operation event for 4,18\n", $time);
            end
            begin
              @(final_operation[4][19]) ;
              //$display("@%0t LEE: Received final operation event for 4,19\n", $time);
            end
            begin
              @(final_operation[4][20]) ;
              //$display("@%0t LEE: Received final operation event for 4,20\n", $time);
            end
            begin
              @(final_operation[4][21]) ;
              //$display("@%0t LEE: Received final operation event for 4,21\n", $time);
            end
            begin
              @(final_operation[4][22]) ;
              //$display("@%0t LEE: Received final operation event for 4,22\n", $time);
            end
            begin
              @(final_operation[4][23]) ;
              //$display("@%0t LEE: Received final operation event for 4,23\n", $time);
            end
            begin
              @(final_operation[4][24]) ;
              //$display("@%0t LEE: Received final operation event for 4,24\n", $time);
            end
            begin
              @(final_operation[4][25]) ;
              //$display("@%0t LEE: Received final operation event for 4,25\n", $time);
            end
            begin
              @(final_operation[4][26]) ;
              //$display("@%0t LEE: Received final operation event for 4,26\n", $time);
            end
            begin
              @(final_operation[4][27]) ;
              //$display("@%0t LEE: Received final operation event for 4,27\n", $time);
            end
            begin
              @(final_operation[4][28]) ;
              //$display("@%0t LEE: Received final operation event for 4,28\n", $time);
            end
            begin
              @(final_operation[4][29]) ;
              //$display("@%0t LEE: Received final operation event for 4,29\n", $time);
            end
            begin
              @(final_operation[4][30]) ;
              //$display("@%0t LEE: Received final operation event for 4,30\n", $time);
            end
            begin
              @(final_operation[4][31]) ;
              //$display("@%0t LEE: Received final operation event for 4,31\n", $time);
            end

            begin
              @(final_operation[5][0]) ;
              //$display("@%0t LEE: Received final operation event for 5,0\n", $time);
            end
            begin
              @(final_operation[5][1]) ;
              //$display("@%0t LEE: Received final operation event for 5,1\n", $time);
            end
            begin
              @(final_operation[5][2]) ;
              //$display("@%0t LEE: Received final operation event for 5,2\n", $time);
            end
            begin
              @(final_operation[5][3]) ;
              //$display("@%0t LEE: Received final operation event for 5,3\n", $time);
            end
            begin
              @(final_operation[5][4]) ;
              //$display("@%0t LEE: Received final operation event for 5,4\n", $time);
            end
            begin
              @(final_operation[5][5]) ;
              //$display("@%0t LEE: Received final operation event for 5,5\n", $time);
            end
            begin
              @(final_operation[5][6]) ;
              //$display("@%0t LEE: Received final operation event for 5,6\n", $time);
            end
            begin
              @(final_operation[5][7]) ;
              //$display("@%0t LEE: Received final operation event for 5,7\n", $time);
            end
            begin
              @(final_operation[5][8]) ;
              //$display("@%0t LEE: Received final operation event for 5,8\n", $time);
            end
            begin
              @(final_operation[5][9]) ;
              //$display("@%0t LEE: Received final operation event for 5,9\n", $time);
            end
            begin
              @(final_operation[5][10]) ;
              //$display("@%0t LEE: Received final operation event for 5,10\n", $time);
            end
            begin
              @(final_operation[5][11]) ;
              //$display("@%0t LEE: Received final operation event for 5,11\n", $time);
            end
            begin
              @(final_operation[5][12]) ;
              //$display("@%0t LEE: Received final operation event for 5,12\n", $time);
            end
            begin
              @(final_operation[5][13]) ;
              //$display("@%0t LEE: Received final operation event for 5,13\n", $time);
            end
            begin
              @(final_operation[5][14]) ;
              //$display("@%0t LEE: Received final operation event for 5,14\n", $time);
            end
            begin
              @(final_operation[5][15]) ;
              //$display("@%0t LEE: Received final operation event for 5,15\n", $time);
            end
            begin
              @(final_operation[5][16]) ;
              //$display("@%0t LEE: Received final operation event for 5,16\n", $time);
            end
            begin
              @(final_operation[5][17]) ;
              //$display("@%0t LEE: Received final operation event for 5,17\n", $time);
            end
            begin
              @(final_operation[5][18]) ;
              //$display("@%0t LEE: Received final operation event for 5,18\n", $time);
            end
            begin
              @(final_operation[5][19]) ;
              //$display("@%0t LEE: Received final operation event for 5,19\n", $time);
            end
            begin
              @(final_operation[5][20]) ;
              //$display("@%0t LEE: Received final operation event for 5,20\n", $time);
            end
            begin
              @(final_operation[5][21]) ;
              //$display("@%0t LEE: Received final operation event for 5,21\n", $time);
            end
            begin
              @(final_operation[5][22]) ;
              //$display("@%0t LEE: Received final operation event for 5,22\n", $time);
            end
            begin
              @(final_operation[5][23]) ;
              //$display("@%0t LEE: Received final operation event for 5,23\n", $time);
            end
            begin
              @(final_operation[5][24]) ;
              //$display("@%0t LEE: Received final operation event for 5,24\n", $time);
            end
            begin
              @(final_operation[5][25]) ;
              //$display("@%0t LEE: Received final operation event for 5,25\n", $time);
            end
            begin
              @(final_operation[5][26]) ;
              //$display("@%0t LEE: Received final operation event for 5,26\n", $time);
            end
            begin
              @(final_operation[5][27]) ;
              //$display("@%0t LEE: Received final operation event for 5,27\n", $time);
            end
            begin
              @(final_operation[5][28]) ;
              //$display("@%0t LEE: Received final operation event for 5,28\n", $time);
            end
            begin
              @(final_operation[5][29]) ;
              //$display("@%0t LEE: Received final operation event for 5,29\n", $time);
            end
            begin
              @(final_operation[5][30]) ;
              //$display("@%0t LEE: Received final operation event for 5,30\n", $time);
            end
            begin
              @(final_operation[5][31]) ;
              //$display("@%0t LEE: Received final operation event for 5,31\n", $time);
            end

            begin
              @(final_operation[6][0]) ;
              //$display("@%0t LEE: Received final operation event for 6,0\n", $time);
            end
            begin
              @(final_operation[6][1]) ;
              //$display("@%0t LEE: Received final operation event for 6,1\n", $time);
            end
            begin
              @(final_operation[6][2]) ;
              //$display("@%0t LEE: Received final operation event for 6,2\n", $time);
            end
            begin
              @(final_operation[6][3]) ;
              //$display("@%0t LEE: Received final operation event for 6,3\n", $time);
            end
            begin
              @(final_operation[6][4]) ;
              //$display("@%0t LEE: Received final operation event for 6,4\n", $time);
            end
            begin
              @(final_operation[6][5]) ;
              //$display("@%0t LEE: Received final operation event for 6,5\n", $time);
            end
            begin
              @(final_operation[6][6]) ;
              //$display("@%0t LEE: Received final operation event for 6,6\n", $time);
            end
            begin
              @(final_operation[6][7]) ;
              //$display("@%0t LEE: Received final operation event for 6,7\n", $time);
            end
            begin
              @(final_operation[6][8]) ;
              //$display("@%0t LEE: Received final operation event for 6,8\n", $time);
            end
            begin
              @(final_operation[6][9]) ;
              //$display("@%0t LEE: Received final operation event for 6,9\n", $time);
            end
            begin
              @(final_operation[6][10]) ;
              //$display("@%0t LEE: Received final operation event for 6,10\n", $time);
            end
            begin
              @(final_operation[6][11]) ;
              //$display("@%0t LEE: Received final operation event for 6,11\n", $time);
            end
            begin
              @(final_operation[6][12]) ;
              //$display("@%0t LEE: Received final operation event for 6,12\n", $time);
            end
            begin
              @(final_operation[6][13]) ;
              //$display("@%0t LEE: Received final operation event for 6,13\n", $time);
            end
            begin
              @(final_operation[6][14]) ;
              //$display("@%0t LEE: Received final operation event for 6,14\n", $time);
            end
            begin
              @(final_operation[6][15]) ;
              //$display("@%0t LEE: Received final operation event for 6,15\n", $time);
            end
            begin
              @(final_operation[6][16]) ;
              //$display("@%0t LEE: Received final operation event for 6,16\n", $time);
            end
            begin
              @(final_operation[6][17]) ;
              //$display("@%0t LEE: Received final operation event for 6,17\n", $time);
            end
            begin
              @(final_operation[6][18]) ;
              //$display("@%0t LEE: Received final operation event for 6,18\n", $time);
            end
            begin
              @(final_operation[6][19]) ;
              //$display("@%0t LEE: Received final operation event for 6,19\n", $time);
            end
            begin
              @(final_operation[6][20]) ;
              //$display("@%0t LEE: Received final operation event for 6,20\n", $time);
            end
            begin
              @(final_operation[6][21]) ;
              //$display("@%0t LEE: Received final operation event for 6,21\n", $time);
            end
            begin
              @(final_operation[6][22]) ;
              //$display("@%0t LEE: Received final operation event for 6,22\n", $time);
            end
            begin
              @(final_operation[6][23]) ;
              //$display("@%0t LEE: Received final operation event for 6,23\n", $time);
            end
            begin
              @(final_operation[6][24]) ;
              //$display("@%0t LEE: Received final operation event for 6,24\n", $time);
            end
            begin
              @(final_operation[6][25]) ;
              //$display("@%0t LEE: Received final operation event for 6,25\n", $time);
            end
            begin
              @(final_operation[6][26]) ;
              //$display("@%0t LEE: Received final operation event for 6,26\n", $time);
            end
            begin
              @(final_operation[6][27]) ;
              //$display("@%0t LEE: Received final operation event for 6,27\n", $time);
            end
            begin
              @(final_operation[6][28]) ;
              //$display("@%0t LEE: Received final operation event for 6,28\n", $time);
            end
            begin
              @(final_operation[6][29]) ;
              //$display("@%0t LEE: Received final operation event for 6,29\n", $time);
            end
            begin
              @(final_operation[6][30]) ;
              //$display("@%0t LEE: Received final operation event for 6,30\n", $time);
            end
            begin
              @(final_operation[6][31]) ;
              //$display("@%0t LEE: Received final operation event for 6,31\n", $time);
            end

            begin
              @(final_operation[7][0]) ;
              //$display("@%0t LEE: Received final operation event for 7,0\n", $time);
            end
            begin
              @(final_operation[7][1]) ;
              //$display("@%0t LEE: Received final operation event for 7,1\n", $time);
            end
            begin
              @(final_operation[7][2]) ;
              //$display("@%0t LEE: Received final operation event for 7,2\n", $time);
            end
            begin
              @(final_operation[7][3]) ;
              //$display("@%0t LEE: Received final operation event for 7,3\n", $time);
            end
            begin
              @(final_operation[7][4]) ;
              //$display("@%0t LEE: Received final operation event for 7,4\n", $time);
            end
            begin
              @(final_operation[7][5]) ;
              //$display("@%0t LEE: Received final operation event for 7,5\n", $time);
            end
            begin
              @(final_operation[7][6]) ;
              //$display("@%0t LEE: Received final operation event for 7,6\n", $time);
            end
            begin
              @(final_operation[7][7]) ;
              //$display("@%0t LEE: Received final operation event for 7,7\n", $time);
            end
            begin
              @(final_operation[7][8]) ;
              //$display("@%0t LEE: Received final operation event for 7,8\n", $time);
            end
            begin
              @(final_operation[7][9]) ;
              //$display("@%0t LEE: Received final operation event for 7,9\n", $time);
            end
            begin
              @(final_operation[7][10]) ;
              //$display("@%0t LEE: Received final operation event for 7,10\n", $time);
            end
            begin
              @(final_operation[7][11]) ;
              //$display("@%0t LEE: Received final operation event for 7,11\n", $time);
            end
            begin
              @(final_operation[7][12]) ;
              //$display("@%0t LEE: Received final operation event for 7,12\n", $time);
            end
            begin
              @(final_operation[7][13]) ;
              //$display("@%0t LEE: Received final operation event for 7,13\n", $time);
            end
            begin
              @(final_operation[7][14]) ;
              //$display("@%0t LEE: Received final operation event for 7,14\n", $time);
            end
            begin
              @(final_operation[7][15]) ;
              //$display("@%0t LEE: Received final operation event for 7,15\n", $time);
            end
            begin
              @(final_operation[7][16]) ;
              //$display("@%0t LEE: Received final operation event for 7,16\n", $time);
            end
            begin
              @(final_operation[7][17]) ;
              //$display("@%0t LEE: Received final operation event for 7,17\n", $time);
            end
            begin
              @(final_operation[7][18]) ;
              //$display("@%0t LEE: Received final operation event for 7,18\n", $time);
            end
            begin
              @(final_operation[7][19]) ;
              //$display("@%0t LEE: Received final operation event for 7,19\n", $time);
            end
            begin
              @(final_operation[7][20]) ;
              //$display("@%0t LEE: Received final operation event for 7,20\n", $time);
            end
            begin
              @(final_operation[7][21]) ;
              //$display("@%0t LEE: Received final operation event for 7,21\n", $time);
            end
            begin
              @(final_operation[7][22]) ;
              //$display("@%0t LEE: Received final operation event for 7,22\n", $time);
            end
            begin
              @(final_operation[7][23]) ;
              //$display("@%0t LEE: Received final operation event for 7,23\n", $time);
            end
            begin
              @(final_operation[7][24]) ;
              //$display("@%0t LEE: Received final operation event for 7,24\n", $time);
            end
            begin
              @(final_operation[7][25]) ;
              //$display("@%0t LEE: Received final operation event for 7,25\n", $time);
            end
            begin
              @(final_operation[7][26]) ;
              //$display("@%0t LEE: Received final operation event for 7,26\n", $time);
            end
            begin
              @(final_operation[7][27]) ;
              //$display("@%0t LEE: Received final operation event for 7,27\n", $time);
            end
            begin
              @(final_operation[7][28]) ;
              //$display("@%0t LEE: Received final operation event for 7,28\n", $time);
            end
            begin
              @(final_operation[7][29]) ;
              //$display("@%0t LEE: Received final operation event for 7,29\n", $time);
            end
            begin
              @(final_operation[7][30]) ;
              //$display("@%0t LEE: Received final operation event for 7,30\n", $time);
            end
            begin
              @(final_operation[7][31]) ;
              //$display("@%0t LEE: Received final operation event for 7,31\n", $time);
            end

            begin
              @(final_operation[8][0]) ;
              //$display("@%0t LEE: Received final operation event for 8,0\n", $time);
            end
            begin
              @(final_operation[8][1]) ;
              //$display("@%0t LEE: Received final operation event for 8,1\n", $time);
            end
            begin
              @(final_operation[8][2]) ;
              //$display("@%0t LEE: Received final operation event for 8,2\n", $time);
            end
            begin
              @(final_operation[8][3]) ;
              //$display("@%0t LEE: Received final operation event for 8,3\n", $time);
            end
            begin
              @(final_operation[8][4]) ;
              //$display("@%0t LEE: Received final operation event for 8,4\n", $time);
            end
            begin
              @(final_operation[8][5]) ;
              //$display("@%0t LEE: Received final operation event for 8,5\n", $time);
            end
            begin
              @(final_operation[8][6]) ;
              //$display("@%0t LEE: Received final operation event for 8,6\n", $time);
            end
            begin
              @(final_operation[8][7]) ;
              //$display("@%0t LEE: Received final operation event for 8,7\n", $time);
            end
            begin
              @(final_operation[8][8]) ;
              //$display("@%0t LEE: Received final operation event for 8,8\n", $time);
            end
            begin
              @(final_operation[8][9]) ;
              //$display("@%0t LEE: Received final operation event for 8,9\n", $time);
            end
            begin
              @(final_operation[8][10]) ;
              //$display("@%0t LEE: Received final operation event for 8,10\n", $time);
            end
            begin
              @(final_operation[8][11]) ;
              //$display("@%0t LEE: Received final operation event for 8,11\n", $time);
            end
            begin
              @(final_operation[8][12]) ;
              //$display("@%0t LEE: Received final operation event for 8,12\n", $time);
            end
            begin
              @(final_operation[8][13]) ;
              //$display("@%0t LEE: Received final operation event for 8,13\n", $time);
            end
            begin
              @(final_operation[8][14]) ;
              //$display("@%0t LEE: Received final operation event for 8,14\n", $time);
            end
            begin
              @(final_operation[8][15]) ;
              //$display("@%0t LEE: Received final operation event for 8,15\n", $time);
            end
            begin
              @(final_operation[8][16]) ;
              //$display("@%0t LEE: Received final operation event for 8,16\n", $time);
            end
            begin
              @(final_operation[8][17]) ;
              //$display("@%0t LEE: Received final operation event for 8,17\n", $time);
            end
            begin
              @(final_operation[8][18]) ;
              //$display("@%0t LEE: Received final operation event for 8,18\n", $time);
            end
            begin
              @(final_operation[8][19]) ;
              //$display("@%0t LEE: Received final operation event for 8,19\n", $time);
            end
            begin
              @(final_operation[8][20]) ;
              //$display("@%0t LEE: Received final operation event for 8,20\n", $time);
            end
            begin
              @(final_operation[8][21]) ;
              //$display("@%0t LEE: Received final operation event for 8,21\n", $time);
            end
            begin
              @(final_operation[8][22]) ;
              //$display("@%0t LEE: Received final operation event for 8,22\n", $time);
            end
            begin
              @(final_operation[8][23]) ;
              //$display("@%0t LEE: Received final operation event for 8,23\n", $time);
            end
            begin
              @(final_operation[8][24]) ;
              //$display("@%0t LEE: Received final operation event for 8,24\n", $time);
            end
            begin
              @(final_operation[8][25]) ;
              //$display("@%0t LEE: Received final operation event for 8,25\n", $time);
            end
            begin
              @(final_operation[8][26]) ;
              //$display("@%0t LEE: Received final operation event for 8,26\n", $time);
            end
            begin
              @(final_operation[8][27]) ;
              //$display("@%0t LEE: Received final operation event for 8,27\n", $time);
            end
            begin
              @(final_operation[8][28]) ;
              //$display("@%0t LEE: Received final operation event for 8,28\n", $time);
            end
            begin
              @(final_operation[8][29]) ;
              //$display("@%0t LEE: Received final operation event for 8,29\n", $time);
            end
            begin
              @(final_operation[8][30]) ;
              //$display("@%0t LEE: Received final operation event for 8,30\n", $time);
            end
            begin
              @(final_operation[8][31]) ;
              //$display("@%0t LEE: Received final operation event for 8,31\n", $time);
            end

            begin
              @(final_operation[9][0]) ;
              //$display("@%0t LEE: Received final operation event for 9,0\n", $time);
            end
            begin
              @(final_operation[9][1]) ;
              //$display("@%0t LEE: Received final operation event for 9,1\n", $time);
            end
            begin
              @(final_operation[9][2]) ;
              //$display("@%0t LEE: Received final operation event for 9,2\n", $time);
            end
            begin
              @(final_operation[9][3]) ;
              //$display("@%0t LEE: Received final operation event for 9,3\n", $time);
            end
            begin
              @(final_operation[9][4]) ;
              //$display("@%0t LEE: Received final operation event for 9,4\n", $time);
            end
            begin
              @(final_operation[9][5]) ;
              //$display("@%0t LEE: Received final operation event for 9,5\n", $time);
            end
            begin
              @(final_operation[9][6]) ;
              //$display("@%0t LEE: Received final operation event for 9,6\n", $time);
            end
            begin
              @(final_operation[9][7]) ;
              //$display("@%0t LEE: Received final operation event for 9,7\n", $time);
            end
            begin
              @(final_operation[9][8]) ;
              //$display("@%0t LEE: Received final operation event for 9,8\n", $time);
            end
            begin
              @(final_operation[9][9]) ;
              //$display("@%0t LEE: Received final operation event for 9,9\n", $time);
            end
            begin
              @(final_operation[9][10]) ;
              //$display("@%0t LEE: Received final operation event for 9,10\n", $time);
            end
            begin
              @(final_operation[9][11]) ;
              //$display("@%0t LEE: Received final operation event for 9,11\n", $time);
            end
            begin
              @(final_operation[9][12]) ;
              //$display("@%0t LEE: Received final operation event for 9,12\n", $time);
            end
            begin
              @(final_operation[9][13]) ;
              //$display("@%0t LEE: Received final operation event for 9,13\n", $time);
            end
            begin
              @(final_operation[9][14]) ;
              //$display("@%0t LEE: Received final operation event for 9,14\n", $time);
            end
            begin
              @(final_operation[9][15]) ;
              //$display("@%0t LEE: Received final operation event for 9,15\n", $time);
            end
            begin
              @(final_operation[9][16]) ;
              //$display("@%0t LEE: Received final operation event for 9,16\n", $time);
            end
            begin
              @(final_operation[9][17]) ;
              //$display("@%0t LEE: Received final operation event for 9,17\n", $time);
            end
            begin
              @(final_operation[9][18]) ;
              //$display("@%0t LEE: Received final operation event for 9,18\n", $time);
            end
            begin
              @(final_operation[9][19]) ;
              //$display("@%0t LEE: Received final operation event for 9,19\n", $time);
            end
            begin
              @(final_operation[9][20]) ;
              //$display("@%0t LEE: Received final operation event for 9,20\n", $time);
            end
            begin
              @(final_operation[9][21]) ;
              //$display("@%0t LEE: Received final operation event for 9,21\n", $time);
            end
            begin
              @(final_operation[9][22]) ;
              //$display("@%0t LEE: Received final operation event for 9,22\n", $time);
            end
            begin
              @(final_operation[9][23]) ;
              //$display("@%0t LEE: Received final operation event for 9,23\n", $time);
            end
            begin
              @(final_operation[9][24]) ;
              //$display("@%0t LEE: Received final operation event for 9,24\n", $time);
            end
            begin
              @(final_operation[9][25]) ;
              //$display("@%0t LEE: Received final operation event for 9,25\n", $time);
            end
            begin
              @(final_operation[9][26]) ;
              //$display("@%0t LEE: Received final operation event for 9,26\n", $time);
            end
            begin
              @(final_operation[9][27]) ;
              //$display("@%0t LEE: Received final operation event for 9,27\n", $time);
            end
            begin
              @(final_operation[9][28]) ;
              //$display("@%0t LEE: Received final operation event for 9,28\n", $time);
            end
            begin
              @(final_operation[9][29]) ;
              //$display("@%0t LEE: Received final operation event for 9,29\n", $time);
            end
            begin
              @(final_operation[9][30]) ;
              //$display("@%0t LEE: Received final operation event for 9,30\n", $time);
            end
            begin
              @(final_operation[9][31]) ;
              //$display("@%0t LEE: Received final operation event for 9,31\n", $time);
            end

            begin
              @(final_operation[10][0]) ;
              //$display("@%0t LEE: Received final operation event for 10,0\n", $time);
            end
            begin
              @(final_operation[10][1]) ;
              //$display("@%0t LEE: Received final operation event for 10,1\n", $time);
            end
            begin
              @(final_operation[10][2]) ;
              //$display("@%0t LEE: Received final operation event for 10,2\n", $time);
            end
            begin
              @(final_operation[10][3]) ;
              //$display("@%0t LEE: Received final operation event for 10,3\n", $time);
            end
            begin
              @(final_operation[10][4]) ;
              //$display("@%0t LEE: Received final operation event for 10,4\n", $time);
            end
            begin
              @(final_operation[10][5]) ;
              //$display("@%0t LEE: Received final operation event for 10,5\n", $time);
            end
            begin
              @(final_operation[10][6]) ;
              //$display("@%0t LEE: Received final operation event for 10,6\n", $time);
            end
            begin
              @(final_operation[10][7]) ;
              //$display("@%0t LEE: Received final operation event for 10,7\n", $time);
            end
            begin
              @(final_operation[10][8]) ;
              //$display("@%0t LEE: Received final operation event for 10,8\n", $time);
            end
            begin
              @(final_operation[10][9]) ;
              //$display("@%0t LEE: Received final operation event for 10,9\n", $time);
            end
            begin
              @(final_operation[10][10]) ;
              //$display("@%0t LEE: Received final operation event for 10,10\n", $time);
            end
            begin
              @(final_operation[10][11]) ;
              //$display("@%0t LEE: Received final operation event for 10,11\n", $time);
            end
            begin
              @(final_operation[10][12]) ;
              //$display("@%0t LEE: Received final operation event for 10,12\n", $time);
            end
            begin
              @(final_operation[10][13]) ;
              //$display("@%0t LEE: Received final operation event for 10,13\n", $time);
            end
            begin
              @(final_operation[10][14]) ;
              //$display("@%0t LEE: Received final operation event for 10,14\n", $time);
            end
            begin
              @(final_operation[10][15]) ;
              //$display("@%0t LEE: Received final operation event for 10,15\n", $time);
            end
            begin
              @(final_operation[10][16]) ;
              //$display("@%0t LEE: Received final operation event for 10,16\n", $time);
            end
            begin
              @(final_operation[10][17]) ;
              //$display("@%0t LEE: Received final operation event for 10,17\n", $time);
            end
            begin
              @(final_operation[10][18]) ;
              //$display("@%0t LEE: Received final operation event for 10,18\n", $time);
            end
            begin
              @(final_operation[10][19]) ;
              //$display("@%0t LEE: Received final operation event for 10,19\n", $time);
            end
            begin
              @(final_operation[10][20]) ;
              //$display("@%0t LEE: Received final operation event for 10,20\n", $time);
            end
            begin
              @(final_operation[10][21]) ;
              //$display("@%0t LEE: Received final operation event for 10,21\n", $time);
            end
            begin
              @(final_operation[10][22]) ;
              //$display("@%0t LEE: Received final operation event for 10,22\n", $time);
            end
            begin
              @(final_operation[10][23]) ;
              //$display("@%0t LEE: Received final operation event for 10,23\n", $time);
            end
            begin
              @(final_operation[10][24]) ;
              //$display("@%0t LEE: Received final operation event for 10,24\n", $time);
            end
            begin
              @(final_operation[10][25]) ;
              //$display("@%0t LEE: Received final operation event for 10,25\n", $time);
            end
            begin
              @(final_operation[10][26]) ;
              //$display("@%0t LEE: Received final operation event for 10,26\n", $time);
            end
            begin
              @(final_operation[10][27]) ;
              //$display("@%0t LEE: Received final operation event for 10,27\n", $time);
            end
            begin
              @(final_operation[10][28]) ;
              //$display("@%0t LEE: Received final operation event for 10,28\n", $time);
            end
            begin
              @(final_operation[10][29]) ;
              //$display("@%0t LEE: Received final operation event for 10,29\n", $time);
            end
            begin
              @(final_operation[10][30]) ;
              //$display("@%0t LEE: Received final operation event for 10,30\n", $time);
            end
            begin
              @(final_operation[10][31]) ;
              //$display("@%0t LEE: Received final operation event for 10,31\n", $time);
            end

            begin
              @(final_operation[11][0]) ;
              //$display("@%0t LEE: Received final operation event for 11,0\n", $time);
            end
            begin
              @(final_operation[11][1]) ;
              //$display("@%0t LEE: Received final operation event for 11,1\n", $time);
            end
            begin
              @(final_operation[11][2]) ;
              //$display("@%0t LEE: Received final operation event for 11,2\n", $time);
            end
            begin
              @(final_operation[11][3]) ;
              //$display("@%0t LEE: Received final operation event for 11,3\n", $time);
            end
            begin
              @(final_operation[11][4]) ;
              //$display("@%0t LEE: Received final operation event for 11,4\n", $time);
            end
            begin
              @(final_operation[11][5]) ;
              //$display("@%0t LEE: Received final operation event for 11,5\n", $time);
            end
            begin
              @(final_operation[11][6]) ;
              //$display("@%0t LEE: Received final operation event for 11,6\n", $time);
            end
            begin
              @(final_operation[11][7]) ;
              //$display("@%0t LEE: Received final operation event for 11,7\n", $time);
            end
            begin
              @(final_operation[11][8]) ;
              //$display("@%0t LEE: Received final operation event for 11,8\n", $time);
            end
            begin
              @(final_operation[11][9]) ;
              //$display("@%0t LEE: Received final operation event for 11,9\n", $time);
            end
            begin
              @(final_operation[11][10]) ;
              //$display("@%0t LEE: Received final operation event for 11,10\n", $time);
            end
            begin
              @(final_operation[11][11]) ;
              //$display("@%0t LEE: Received final operation event for 11,11\n", $time);
            end
            begin
              @(final_operation[11][12]) ;
              //$display("@%0t LEE: Received final operation event for 11,12\n", $time);
            end
            begin
              @(final_operation[11][13]) ;
              //$display("@%0t LEE: Received final operation event for 11,13\n", $time);
            end
            begin
              @(final_operation[11][14]) ;
              //$display("@%0t LEE: Received final operation event for 11,14\n", $time);
            end
            begin
              @(final_operation[11][15]) ;
              //$display("@%0t LEE: Received final operation event for 11,15\n", $time);
            end
            begin
              @(final_operation[11][16]) ;
              //$display("@%0t LEE: Received final operation event for 11,16\n", $time);
            end
            begin
              @(final_operation[11][17]) ;
              //$display("@%0t LEE: Received final operation event for 11,17\n", $time);
            end
            begin
              @(final_operation[11][18]) ;
              //$display("@%0t LEE: Received final operation event for 11,18\n", $time);
            end
            begin
              @(final_operation[11][19]) ;
              //$display("@%0t LEE: Received final operation event for 11,19\n", $time);
            end
            begin
              @(final_operation[11][20]) ;
              //$display("@%0t LEE: Received final operation event for 11,20\n", $time);
            end
            begin
              @(final_operation[11][21]) ;
              //$display("@%0t LEE: Received final operation event for 11,21\n", $time);
            end
            begin
              @(final_operation[11][22]) ;
              //$display("@%0t LEE: Received final operation event for 11,22\n", $time);
            end
            begin
              @(final_operation[11][23]) ;
              //$display("@%0t LEE: Received final operation event for 11,23\n", $time);
            end
            begin
              @(final_operation[11][24]) ;
              //$display("@%0t LEE: Received final operation event for 11,24\n", $time);
            end
            begin
              @(final_operation[11][25]) ;
              //$display("@%0t LEE: Received final operation event for 11,25\n", $time);
            end
            begin
              @(final_operation[11][26]) ;
              //$display("@%0t LEE: Received final operation event for 11,26\n", $time);
            end
            begin
              @(final_operation[11][27]) ;
              //$display("@%0t LEE: Received final operation event for 11,27\n", $time);
            end
            begin
              @(final_operation[11][28]) ;
              //$display("@%0t LEE: Received final operation event for 11,28\n", $time);
            end
            begin
              @(final_operation[11][29]) ;
              //$display("@%0t LEE: Received final operation event for 11,29\n", $time);
            end
            begin
              @(final_operation[11][30]) ;
              //$display("@%0t LEE: Received final operation event for 11,30\n", $time);
            end
            begin
              @(final_operation[11][31]) ;
              //$display("@%0t LEE: Received final operation event for 11,31\n", $time);
            end

            begin
              @(final_operation[12][0]) ;
              //$display("@%0t LEE: Received final operation event for 12,0\n", $time);
            end
            begin
              @(final_operation[12][1]) ;
              //$display("@%0t LEE: Received final operation event for 12,1\n", $time);
            end
            begin
              @(final_operation[12][2]) ;
              //$display("@%0t LEE: Received final operation event for 12,2\n", $time);
            end
            begin
              @(final_operation[12][3]) ;
              //$display("@%0t LEE: Received final operation event for 12,3\n", $time);
            end
            begin
              @(final_operation[12][4]) ;
              //$display("@%0t LEE: Received final operation event for 12,4\n", $time);
            end
            begin
              @(final_operation[12][5]) ;
              //$display("@%0t LEE: Received final operation event for 12,5\n", $time);
            end
            begin
              @(final_operation[12][6]) ;
              //$display("@%0t LEE: Received final operation event for 12,6\n", $time);
            end
            begin
              @(final_operation[12][7]) ;
              //$display("@%0t LEE: Received final operation event for 12,7\n", $time);
            end
            begin
              @(final_operation[12][8]) ;
              //$display("@%0t LEE: Received final operation event for 12,8\n", $time);
            end
            begin
              @(final_operation[12][9]) ;
              //$display("@%0t LEE: Received final operation event for 12,9\n", $time);
            end
            begin
              @(final_operation[12][10]) ;
              //$display("@%0t LEE: Received final operation event for 12,10\n", $time);
            end
            begin
              @(final_operation[12][11]) ;
              //$display("@%0t LEE: Received final operation event for 12,11\n", $time);
            end
            begin
              @(final_operation[12][12]) ;
              //$display("@%0t LEE: Received final operation event for 12,12\n", $time);
            end
            begin
              @(final_operation[12][13]) ;
              //$display("@%0t LEE: Received final operation event for 12,13\n", $time);
            end
            begin
              @(final_operation[12][14]) ;
              //$display("@%0t LEE: Received final operation event for 12,14\n", $time);
            end
            begin
              @(final_operation[12][15]) ;
              //$display("@%0t LEE: Received final operation event for 12,15\n", $time);
            end
            begin
              @(final_operation[12][16]) ;
              //$display("@%0t LEE: Received final operation event for 12,16\n", $time);
            end
            begin
              @(final_operation[12][17]) ;
              //$display("@%0t LEE: Received final operation event for 12,17\n", $time);
            end
            begin
              @(final_operation[12][18]) ;
              //$display("@%0t LEE: Received final operation event for 12,18\n", $time);
            end
            begin
              @(final_operation[12][19]) ;
              //$display("@%0t LEE: Received final operation event for 12,19\n", $time);
            end
            begin
              @(final_operation[12][20]) ;
              //$display("@%0t LEE: Received final operation event for 12,20\n", $time);
            end
            begin
              @(final_operation[12][21]) ;
              //$display("@%0t LEE: Received final operation event for 12,21\n", $time);
            end
            begin
              @(final_operation[12][22]) ;
              //$display("@%0t LEE: Received final operation event for 12,22\n", $time);
            end
            begin
              @(final_operation[12][23]) ;
              //$display("@%0t LEE: Received final operation event for 12,23\n", $time);
            end
            begin
              @(final_operation[12][24]) ;
              //$display("@%0t LEE: Received final operation event for 12,24\n", $time);
            end
            begin
              @(final_operation[12][25]) ;
              //$display("@%0t LEE: Received final operation event for 12,25\n", $time);
            end
            begin
              @(final_operation[12][26]) ;
              //$display("@%0t LEE: Received final operation event for 12,26\n", $time);
            end
            begin
              @(final_operation[12][27]) ;
              //$display("@%0t LEE: Received final operation event for 12,27\n", $time);
            end
            begin
              @(final_operation[12][28]) ;
              //$display("@%0t LEE: Received final operation event for 12,28\n", $time);
            end
            begin
              @(final_operation[12][29]) ;
              //$display("@%0t LEE: Received final operation event for 12,29\n", $time);
            end
            begin
              @(final_operation[12][30]) ;
              //$display("@%0t LEE: Received final operation event for 12,30\n", $time);
            end
            begin
              @(final_operation[12][31]) ;
              //$display("@%0t LEE: Received final operation event for 12,31\n", $time);
            end

            begin
              @(final_operation[13][0]) ;
              //$display("@%0t LEE: Received final operation event for 13,0\n", $time);
            end
            begin
              @(final_operation[13][1]) ;
              //$display("@%0t LEE: Received final operation event for 13,1\n", $time);
            end
            begin
              @(final_operation[13][2]) ;
              //$display("@%0t LEE: Received final operation event for 13,2\n", $time);
            end
            begin
              @(final_operation[13][3]) ;
              //$display("@%0t LEE: Received final operation event for 13,3\n", $time);
            end
            begin
              @(final_operation[13][4]) ;
              //$display("@%0t LEE: Received final operation event for 13,4\n", $time);
            end
            begin
              @(final_operation[13][5]) ;
              //$display("@%0t LEE: Received final operation event for 13,5\n", $time);
            end
            begin
              @(final_operation[13][6]) ;
              //$display("@%0t LEE: Received final operation event for 13,6\n", $time);
            end
            begin
              @(final_operation[13][7]) ;
              //$display("@%0t LEE: Received final operation event for 13,7\n", $time);
            end
            begin
              @(final_operation[13][8]) ;
              //$display("@%0t LEE: Received final operation event for 13,8\n", $time);
            end
            begin
              @(final_operation[13][9]) ;
              //$display("@%0t LEE: Received final operation event for 13,9\n", $time);
            end
            begin
              @(final_operation[13][10]) ;
              //$display("@%0t LEE: Received final operation event for 13,10\n", $time);
            end
            begin
              @(final_operation[13][11]) ;
              //$display("@%0t LEE: Received final operation event for 13,11\n", $time);
            end
            begin
              @(final_operation[13][12]) ;
              //$display("@%0t LEE: Received final operation event for 13,12\n", $time);
            end
            begin
              @(final_operation[13][13]) ;
              //$display("@%0t LEE: Received final operation event for 13,13\n", $time);
            end
            begin
              @(final_operation[13][14]) ;
              //$display("@%0t LEE: Received final operation event for 13,14\n", $time);
            end
            begin
              @(final_operation[13][15]) ;
              //$display("@%0t LEE: Received final operation event for 13,15\n", $time);
            end
            begin
              @(final_operation[13][16]) ;
              //$display("@%0t LEE: Received final operation event for 13,16\n", $time);
            end
            begin
              @(final_operation[13][17]) ;
              //$display("@%0t LEE: Received final operation event for 13,17\n", $time);
            end
            begin
              @(final_operation[13][18]) ;
              //$display("@%0t LEE: Received final operation event for 13,18\n", $time);
            end
            begin
              @(final_operation[13][19]) ;
              //$display("@%0t LEE: Received final operation event for 13,19\n", $time);
            end
            begin
              @(final_operation[13][20]) ;
              //$display("@%0t LEE: Received final operation event for 13,20\n", $time);
            end
            begin
              @(final_operation[13][21]) ;
              //$display("@%0t LEE: Received final operation event for 13,21\n", $time);
            end
            begin
              @(final_operation[13][22]) ;
              //$display("@%0t LEE: Received final operation event for 13,22\n", $time);
            end
            begin
              @(final_operation[13][23]) ;
              //$display("@%0t LEE: Received final operation event for 13,23\n", $time);
            end
            begin
              @(final_operation[13][24]) ;
              //$display("@%0t LEE: Received final operation event for 13,24\n", $time);
            end
            begin
              @(final_operation[13][25]) ;
              //$display("@%0t LEE: Received final operation event for 13,25\n", $time);
            end
            begin
              @(final_operation[13][26]) ;
              //$display("@%0t LEE: Received final operation event for 13,26\n", $time);
            end
            begin
              @(final_operation[13][27]) ;
              //$display("@%0t LEE: Received final operation event for 13,27\n", $time);
            end
            begin
              @(final_operation[13][28]) ;
              //$display("@%0t LEE: Received final operation event for 13,28\n", $time);
            end
            begin
              @(final_operation[13][29]) ;
              //$display("@%0t LEE: Received final operation event for 13,29\n", $time);
            end
            begin
              @(final_operation[13][30]) ;
              //$display("@%0t LEE: Received final operation event for 13,30\n", $time);
            end
            begin
              @(final_operation[13][31]) ;
              //$display("@%0t LEE: Received final operation event for 13,31\n", $time);
            end

            begin
              @(final_operation[14][0]) ;
              //$display("@%0t LEE: Received final operation event for 14,0\n", $time);
            end
            begin
              @(final_operation[14][1]) ;
              //$display("@%0t LEE: Received final operation event for 14,1\n", $time);
            end
            begin
              @(final_operation[14][2]) ;
              //$display("@%0t LEE: Received final operation event for 14,2\n", $time);
            end
            begin
              @(final_operation[14][3]) ;
              //$display("@%0t LEE: Received final operation event for 14,3\n", $time);
            end
            begin
              @(final_operation[14][4]) ;
              //$display("@%0t LEE: Received final operation event for 14,4\n", $time);
            end
            begin
              @(final_operation[14][5]) ;
              //$display("@%0t LEE: Received final operation event for 14,5\n", $time);
            end
            begin
              @(final_operation[14][6]) ;
              //$display("@%0t LEE: Received final operation event for 14,6\n", $time);
            end
            begin
              @(final_operation[14][7]) ;
              //$display("@%0t LEE: Received final operation event for 14,7\n", $time);
            end
            begin
              @(final_operation[14][8]) ;
              //$display("@%0t LEE: Received final operation event for 14,8\n", $time);
            end
            begin
              @(final_operation[14][9]) ;
              //$display("@%0t LEE: Received final operation event for 14,9\n", $time);
            end
            begin
              @(final_operation[14][10]) ;
              //$display("@%0t LEE: Received final operation event for 14,10\n", $time);
            end
            begin
              @(final_operation[14][11]) ;
              //$display("@%0t LEE: Received final operation event for 14,11\n", $time);
            end
            begin
              @(final_operation[14][12]) ;
              //$display("@%0t LEE: Received final operation event for 14,12\n", $time);
            end
            begin
              @(final_operation[14][13]) ;
              //$display("@%0t LEE: Received final operation event for 14,13\n", $time);
            end
            begin
              @(final_operation[14][14]) ;
              //$display("@%0t LEE: Received final operation event for 14,14\n", $time);
            end
            begin
              @(final_operation[14][15]) ;
              //$display("@%0t LEE: Received final operation event for 14,15\n", $time);
            end
            begin
              @(final_operation[14][16]) ;
              //$display("@%0t LEE: Received final operation event for 14,16\n", $time);
            end
            begin
              @(final_operation[14][17]) ;
              //$display("@%0t LEE: Received final operation event for 14,17\n", $time);
            end
            begin
              @(final_operation[14][18]) ;
              //$display("@%0t LEE: Received final operation event for 14,18\n", $time);
            end
            begin
              @(final_operation[14][19]) ;
              //$display("@%0t LEE: Received final operation event for 14,19\n", $time);
            end
            begin
              @(final_operation[14][20]) ;
              //$display("@%0t LEE: Received final operation event for 14,20\n", $time);
            end
            begin
              @(final_operation[14][21]) ;
              //$display("@%0t LEE: Received final operation event for 14,21\n", $time);
            end
            begin
              @(final_operation[14][22]) ;
              //$display("@%0t LEE: Received final operation event for 14,22\n", $time);
            end
            begin
              @(final_operation[14][23]) ;
              //$display("@%0t LEE: Received final operation event for 14,23\n", $time);
            end
            begin
              @(final_operation[14][24]) ;
              //$display("@%0t LEE: Received final operation event for 14,24\n", $time);
            end
            begin
              @(final_operation[14][25]) ;
              //$display("@%0t LEE: Received final operation event for 14,25\n", $time);
            end
            begin
              @(final_operation[14][26]) ;
              //$display("@%0t LEE: Received final operation event for 14,26\n", $time);
            end
            begin
              @(final_operation[14][27]) ;
              //$display("@%0t LEE: Received final operation event for 14,27\n", $time);
            end
            begin
              @(final_operation[14][28]) ;
              //$display("@%0t LEE: Received final operation event for 14,28\n", $time);
            end
            begin
              @(final_operation[14][29]) ;
              //$display("@%0t LEE: Received final operation event for 14,29\n", $time);
            end
            begin
              @(final_operation[14][30]) ;
              //$display("@%0t LEE: Received final operation event for 14,30\n", $time);
            end
            begin
              @(final_operation[14][31]) ;
              //$display("@%0t LEE: Received final operation event for 14,31\n", $time);
            end

            begin
              @(final_operation[15][0]) ;
              //$display("@%0t LEE: Received final operation event for 15,0\n", $time);
            end
            begin
              @(final_operation[15][1]) ;
              //$display("@%0t LEE: Received final operation event for 15,1\n", $time);
            end
            begin
              @(final_operation[15][2]) ;
              //$display("@%0t LEE: Received final operation event for 15,2\n", $time);
            end
            begin
              @(final_operation[15][3]) ;
              //$display("@%0t LEE: Received final operation event for 15,3\n", $time);
            end
            begin
              @(final_operation[15][4]) ;
              //$display("@%0t LEE: Received final operation event for 15,4\n", $time);
            end
            begin
              @(final_operation[15][5]) ;
              //$display("@%0t LEE: Received final operation event for 15,5\n", $time);
            end
            begin
              @(final_operation[15][6]) ;
              //$display("@%0t LEE: Received final operation event for 15,6\n", $time);
            end
            begin
              @(final_operation[15][7]) ;
              //$display("@%0t LEE: Received final operation event for 15,7\n", $time);
            end
            begin
              @(final_operation[15][8]) ;
              //$display("@%0t LEE: Received final operation event for 15,8\n", $time);
            end
            begin
              @(final_operation[15][9]) ;
              //$display("@%0t LEE: Received final operation event for 15,9\n", $time);
            end
            begin
              @(final_operation[15][10]) ;
              //$display("@%0t LEE: Received final operation event for 15,10\n", $time);
            end
            begin
              @(final_operation[15][11]) ;
              //$display("@%0t LEE: Received final operation event for 15,11\n", $time);
            end
            begin
              @(final_operation[15][12]) ;
              //$display("@%0t LEE: Received final operation event for 15,12\n", $time);
            end
            begin
              @(final_operation[15][13]) ;
              //$display("@%0t LEE: Received final operation event for 15,13\n", $time);
            end
            begin
              @(final_operation[15][14]) ;
              //$display("@%0t LEE: Received final operation event for 15,14\n", $time);
            end
            begin
              @(final_operation[15][15]) ;
              //$display("@%0t LEE: Received final operation event for 15,15\n", $time);
            end
            begin
              @(final_operation[15][16]) ;
              //$display("@%0t LEE: Received final operation event for 15,16\n", $time);
            end
            begin
              @(final_operation[15][17]) ;
              //$display("@%0t LEE: Received final operation event for 15,17\n", $time);
            end
            begin
              @(final_operation[15][18]) ;
              //$display("@%0t LEE: Received final operation event for 15,18\n", $time);
            end
            begin
              @(final_operation[15][19]) ;
              //$display("@%0t LEE: Received final operation event for 15,19\n", $time);
            end
            begin
              @(final_operation[15][20]) ;
              //$display("@%0t LEE: Received final operation event for 15,20\n", $time);
            end
            begin
              @(final_operation[15][21]) ;
              //$display("@%0t LEE: Received final operation event for 15,21\n", $time);
            end
            begin
              @(final_operation[15][22]) ;
              //$display("@%0t LEE: Received final operation event for 15,22\n", $time);
            end
            begin
              @(final_operation[15][23]) ;
              //$display("@%0t LEE: Received final operation event for 15,23\n", $time);
            end
            begin
              @(final_operation[15][24]) ;
              //$display("@%0t LEE: Received final operation event for 15,24\n", $time);
            end
            begin
              @(final_operation[15][25]) ;
              //$display("@%0t LEE: Received final operation event for 15,25\n", $time);
            end
            begin
              @(final_operation[15][26]) ;
              //$display("@%0t LEE: Received final operation event for 15,26\n", $time);
            end
            begin
              @(final_operation[15][27]) ;
              //$display("@%0t LEE: Received final operation event for 15,27\n", $time);
            end
            begin
              @(final_operation[15][28]) ;
              //$display("@%0t LEE: Received final operation event for 15,28\n", $time);
            end
            begin
              @(final_operation[15][29]) ;
              //$display("@%0t LEE: Received final operation event for 15,29\n", $time);
            end
            begin
              @(final_operation[15][30]) ;
              //$display("@%0t LEE: Received final operation event for 15,30\n", $time);
            end
            begin
              @(final_operation[15][31]) ;
              //$display("@%0t LEE: Received final operation event for 15,31\n", $time);
            end

            begin
              @(final_operation[16][0]) ;
              //$display("@%0t LEE: Received final operation event for 16,0\n", $time);
            end
            begin
              @(final_operation[16][1]) ;
              //$display("@%0t LEE: Received final operation event for 16,1\n", $time);
            end
            begin
              @(final_operation[16][2]) ;
              //$display("@%0t LEE: Received final operation event for 16,2\n", $time);
            end
            begin
              @(final_operation[16][3]) ;
              //$display("@%0t LEE: Received final operation event for 16,3\n", $time);
            end
            begin
              @(final_operation[16][4]) ;
              //$display("@%0t LEE: Received final operation event for 16,4\n", $time);
            end
            begin
              @(final_operation[16][5]) ;
              //$display("@%0t LEE: Received final operation event for 16,5\n", $time);
            end
            begin
              @(final_operation[16][6]) ;
              //$display("@%0t LEE: Received final operation event for 16,6\n", $time);
            end
            begin
              @(final_operation[16][7]) ;
              //$display("@%0t LEE: Received final operation event for 16,7\n", $time);
            end
            begin
              @(final_operation[16][8]) ;
              //$display("@%0t LEE: Received final operation event for 16,8\n", $time);
            end
            begin
              @(final_operation[16][9]) ;
              //$display("@%0t LEE: Received final operation event for 16,9\n", $time);
            end
            begin
              @(final_operation[16][10]) ;
              //$display("@%0t LEE: Received final operation event for 16,10\n", $time);
            end
            begin
              @(final_operation[16][11]) ;
              //$display("@%0t LEE: Received final operation event for 16,11\n", $time);
            end
            begin
              @(final_operation[16][12]) ;
              //$display("@%0t LEE: Received final operation event for 16,12\n", $time);
            end
            begin
              @(final_operation[16][13]) ;
              //$display("@%0t LEE: Received final operation event for 16,13\n", $time);
            end
            begin
              @(final_operation[16][14]) ;
              //$display("@%0t LEE: Received final operation event for 16,14\n", $time);
            end
            begin
              @(final_operation[16][15]) ;
              //$display("@%0t LEE: Received final operation event for 16,15\n", $time);
            end
            begin
              @(final_operation[16][16]) ;
              //$display("@%0t LEE: Received final operation event for 16,16\n", $time);
            end
            begin
              @(final_operation[16][17]) ;
              //$display("@%0t LEE: Received final operation event for 16,17\n", $time);
            end
            begin
              @(final_operation[16][18]) ;
              //$display("@%0t LEE: Received final operation event for 16,18\n", $time);
            end
            begin
              @(final_operation[16][19]) ;
              //$display("@%0t LEE: Received final operation event for 16,19\n", $time);
            end
            begin
              @(final_operation[16][20]) ;
              //$display("@%0t LEE: Received final operation event for 16,20\n", $time);
            end
            begin
              @(final_operation[16][21]) ;
              //$display("@%0t LEE: Received final operation event for 16,21\n", $time);
            end
            begin
              @(final_operation[16][22]) ;
              //$display("@%0t LEE: Received final operation event for 16,22\n", $time);
            end
            begin
              @(final_operation[16][23]) ;
              //$display("@%0t LEE: Received final operation event for 16,23\n", $time);
            end
            begin
              @(final_operation[16][24]) ;
              //$display("@%0t LEE: Received final operation event for 16,24\n", $time);
            end
            begin
              @(final_operation[16][25]) ;
              //$display("@%0t LEE: Received final operation event for 16,25\n", $time);
            end
            begin
              @(final_operation[16][26]) ;
              //$display("@%0t LEE: Received final operation event for 16,26\n", $time);
            end
            begin
              @(final_operation[16][27]) ;
              //$display("@%0t LEE: Received final operation event for 16,27\n", $time);
            end
            begin
              @(final_operation[16][28]) ;
              //$display("@%0t LEE: Received final operation event for 16,28\n", $time);
            end
            begin
              @(final_operation[16][29]) ;
              //$display("@%0t LEE: Received final operation event for 16,29\n", $time);
            end
            begin
              @(final_operation[16][30]) ;
              //$display("@%0t LEE: Received final operation event for 16,30\n", $time);
            end
            begin
              @(final_operation[16][31]) ;
              //$display("@%0t LEE: Received final operation event for 16,31\n", $time);
            end

            begin
              @(final_operation[17][0]) ;
              //$display("@%0t LEE: Received final operation event for 17,0\n", $time);
            end
            begin
              @(final_operation[17][1]) ;
              //$display("@%0t LEE: Received final operation event for 17,1\n", $time);
            end
            begin
              @(final_operation[17][2]) ;
              //$display("@%0t LEE: Received final operation event for 17,2\n", $time);
            end
            begin
              @(final_operation[17][3]) ;
              //$display("@%0t LEE: Received final operation event for 17,3\n", $time);
            end
            begin
              @(final_operation[17][4]) ;
              //$display("@%0t LEE: Received final operation event for 17,4\n", $time);
            end
            begin
              @(final_operation[17][5]) ;
              //$display("@%0t LEE: Received final operation event for 17,5\n", $time);
            end
            begin
              @(final_operation[17][6]) ;
              //$display("@%0t LEE: Received final operation event for 17,6\n", $time);
            end
            begin
              @(final_operation[17][7]) ;
              //$display("@%0t LEE: Received final operation event for 17,7\n", $time);
            end
            begin
              @(final_operation[17][8]) ;
              //$display("@%0t LEE: Received final operation event for 17,8\n", $time);
            end
            begin
              @(final_operation[17][9]) ;
              //$display("@%0t LEE: Received final operation event for 17,9\n", $time);
            end
            begin
              @(final_operation[17][10]) ;
              //$display("@%0t LEE: Received final operation event for 17,10\n", $time);
            end
            begin
              @(final_operation[17][11]) ;
              //$display("@%0t LEE: Received final operation event for 17,11\n", $time);
            end
            begin
              @(final_operation[17][12]) ;
              //$display("@%0t LEE: Received final operation event for 17,12\n", $time);
            end
            begin
              @(final_operation[17][13]) ;
              //$display("@%0t LEE: Received final operation event for 17,13\n", $time);
            end
            begin
              @(final_operation[17][14]) ;
              //$display("@%0t LEE: Received final operation event for 17,14\n", $time);
            end
            begin
              @(final_operation[17][15]) ;
              //$display("@%0t LEE: Received final operation event for 17,15\n", $time);
            end
            begin
              @(final_operation[17][16]) ;
              //$display("@%0t LEE: Received final operation event for 17,16\n", $time);
            end
            begin
              @(final_operation[17][17]) ;
              //$display("@%0t LEE: Received final operation event for 17,17\n", $time);
            end
            begin
              @(final_operation[17][18]) ;
              //$display("@%0t LEE: Received final operation event for 17,18\n", $time);
            end
            begin
              @(final_operation[17][19]) ;
              //$display("@%0t LEE: Received final operation event for 17,19\n", $time);
            end
            begin
              @(final_operation[17][20]) ;
              //$display("@%0t LEE: Received final operation event for 17,20\n", $time);
            end
            begin
              @(final_operation[17][21]) ;
              //$display("@%0t LEE: Received final operation event for 17,21\n", $time);
            end
            begin
              @(final_operation[17][22]) ;
              //$display("@%0t LEE: Received final operation event for 17,22\n", $time);
            end
            begin
              @(final_operation[17][23]) ;
              //$display("@%0t LEE: Received final operation event for 17,23\n", $time);
            end
            begin
              @(final_operation[17][24]) ;
              //$display("@%0t LEE: Received final operation event for 17,24\n", $time);
            end
            begin
              @(final_operation[17][25]) ;
              //$display("@%0t LEE: Received final operation event for 17,25\n", $time);
            end
            begin
              @(final_operation[17][26]) ;
              //$display("@%0t LEE: Received final operation event for 17,26\n", $time);
            end
            begin
              @(final_operation[17][27]) ;
              //$display("@%0t LEE: Received final operation event for 17,27\n", $time);
            end
            begin
              @(final_operation[17][28]) ;
              //$display("@%0t LEE: Received final operation event for 17,28\n", $time);
            end
            begin
              @(final_operation[17][29]) ;
              //$display("@%0t LEE: Received final operation event for 17,29\n", $time);
            end
            begin
              @(final_operation[17][30]) ;
              //$display("@%0t LEE: Received final operation event for 17,30\n", $time);
            end
            begin
              @(final_operation[17][31]) ;
              //$display("@%0t LEE: Received final operation event for 17,31\n", $time);
            end

            begin
              @(final_operation[18][0]) ;
              //$display("@%0t LEE: Received final operation event for 18,0\n", $time);
            end
            begin
              @(final_operation[18][1]) ;
              //$display("@%0t LEE: Received final operation event for 18,1\n", $time);
            end
            begin
              @(final_operation[18][2]) ;
              //$display("@%0t LEE: Received final operation event for 18,2\n", $time);
            end
            begin
              @(final_operation[18][3]) ;
              //$display("@%0t LEE: Received final operation event for 18,3\n", $time);
            end
            begin
              @(final_operation[18][4]) ;
              //$display("@%0t LEE: Received final operation event for 18,4\n", $time);
            end
            begin
              @(final_operation[18][5]) ;
              //$display("@%0t LEE: Received final operation event for 18,5\n", $time);
            end
            begin
              @(final_operation[18][6]) ;
              //$display("@%0t LEE: Received final operation event for 18,6\n", $time);
            end
            begin
              @(final_operation[18][7]) ;
              //$display("@%0t LEE: Received final operation event for 18,7\n", $time);
            end
            begin
              @(final_operation[18][8]) ;
              //$display("@%0t LEE: Received final operation event for 18,8\n", $time);
            end
            begin
              @(final_operation[18][9]) ;
              //$display("@%0t LEE: Received final operation event for 18,9\n", $time);
            end
            begin
              @(final_operation[18][10]) ;
              //$display("@%0t LEE: Received final operation event for 18,10\n", $time);
            end
            begin
              @(final_operation[18][11]) ;
              //$display("@%0t LEE: Received final operation event for 18,11\n", $time);
            end
            begin
              @(final_operation[18][12]) ;
              //$display("@%0t LEE: Received final operation event for 18,12\n", $time);
            end
            begin
              @(final_operation[18][13]) ;
              //$display("@%0t LEE: Received final operation event for 18,13\n", $time);
            end
            begin
              @(final_operation[18][14]) ;
              //$display("@%0t LEE: Received final operation event for 18,14\n", $time);
            end
            begin
              @(final_operation[18][15]) ;
              //$display("@%0t LEE: Received final operation event for 18,15\n", $time);
            end
            begin
              @(final_operation[18][16]) ;
              //$display("@%0t LEE: Received final operation event for 18,16\n", $time);
            end
            begin
              @(final_operation[18][17]) ;
              //$display("@%0t LEE: Received final operation event for 18,17\n", $time);
            end
            begin
              @(final_operation[18][18]) ;
              //$display("@%0t LEE: Received final operation event for 18,18\n", $time);
            end
            begin
              @(final_operation[18][19]) ;
              //$display("@%0t LEE: Received final operation event for 18,19\n", $time);
            end
            begin
              @(final_operation[18][20]) ;
              //$display("@%0t LEE: Received final operation event for 18,20\n", $time);
            end
            begin
              @(final_operation[18][21]) ;
              //$display("@%0t LEE: Received final operation event for 18,21\n", $time);
            end
            begin
              @(final_operation[18][22]) ;
              //$display("@%0t LEE: Received final operation event for 18,22\n", $time);
            end
            begin
              @(final_operation[18][23]) ;
              //$display("@%0t LEE: Received final operation event for 18,23\n", $time);
            end
            begin
              @(final_operation[18][24]) ;
              //$display("@%0t LEE: Received final operation event for 18,24\n", $time);
            end
            begin
              @(final_operation[18][25]) ;
              //$display("@%0t LEE: Received final operation event for 18,25\n", $time);
            end
            begin
              @(final_operation[18][26]) ;
              //$display("@%0t LEE: Received final operation event for 18,26\n", $time);
            end
            begin
              @(final_operation[18][27]) ;
              //$display("@%0t LEE: Received final operation event for 18,27\n", $time);
            end
            begin
              @(final_operation[18][28]) ;
              //$display("@%0t LEE: Received final operation event for 18,28\n", $time);
            end
            begin
              @(final_operation[18][29]) ;
              //$display("@%0t LEE: Received final operation event for 18,29\n", $time);
            end
            begin
              @(final_operation[18][30]) ;
              //$display("@%0t LEE: Received final operation event for 18,30\n", $time);
            end
            begin
              @(final_operation[18][31]) ;
              //$display("@%0t LEE: Received final operation event for 18,31\n", $time);
            end

            begin
              @(final_operation[19][0]) ;
              //$display("@%0t LEE: Received final operation event for 19,0\n", $time);
            end
            begin
              @(final_operation[19][1]) ;
              //$display("@%0t LEE: Received final operation event for 19,1\n", $time);
            end
            begin
              @(final_operation[19][2]) ;
              //$display("@%0t LEE: Received final operation event for 19,2\n", $time);
            end
            begin
              @(final_operation[19][3]) ;
              //$display("@%0t LEE: Received final operation event for 19,3\n", $time);
            end
            begin
              @(final_operation[19][4]) ;
              //$display("@%0t LEE: Received final operation event for 19,4\n", $time);
            end
            begin
              @(final_operation[19][5]) ;
              //$display("@%0t LEE: Received final operation event for 19,5\n", $time);
            end
            begin
              @(final_operation[19][6]) ;
              //$display("@%0t LEE: Received final operation event for 19,6\n", $time);
            end
            begin
              @(final_operation[19][7]) ;
              //$display("@%0t LEE: Received final operation event for 19,7\n", $time);
            end
            begin
              @(final_operation[19][8]) ;
              //$display("@%0t LEE: Received final operation event for 19,8\n", $time);
            end
            begin
              @(final_operation[19][9]) ;
              //$display("@%0t LEE: Received final operation event for 19,9\n", $time);
            end
            begin
              @(final_operation[19][10]) ;
              //$display("@%0t LEE: Received final operation event for 19,10\n", $time);
            end
            begin
              @(final_operation[19][11]) ;
              //$display("@%0t LEE: Received final operation event for 19,11\n", $time);
            end
            begin
              @(final_operation[19][12]) ;
              //$display("@%0t LEE: Received final operation event for 19,12\n", $time);
            end
            begin
              @(final_operation[19][13]) ;
              //$display("@%0t LEE: Received final operation event for 19,13\n", $time);
            end
            begin
              @(final_operation[19][14]) ;
              //$display("@%0t LEE: Received final operation event for 19,14\n", $time);
            end
            begin
              @(final_operation[19][15]) ;
              //$display("@%0t LEE: Received final operation event for 19,15\n", $time);
            end
            begin
              @(final_operation[19][16]) ;
              //$display("@%0t LEE: Received final operation event for 19,16\n", $time);
            end
            begin
              @(final_operation[19][17]) ;
              //$display("@%0t LEE: Received final operation event for 19,17\n", $time);
            end
            begin
              @(final_operation[19][18]) ;
              //$display("@%0t LEE: Received final operation event for 19,18\n", $time);
            end
            begin
              @(final_operation[19][19]) ;
              //$display("@%0t LEE: Received final operation event for 19,19\n", $time);
            end
            begin
              @(final_operation[19][20]) ;
              //$display("@%0t LEE: Received final operation event for 19,20\n", $time);
            end
            begin
              @(final_operation[19][21]) ;
              //$display("@%0t LEE: Received final operation event for 19,21\n", $time);
            end
            begin
              @(final_operation[19][22]) ;
              //$display("@%0t LEE: Received final operation event for 19,22\n", $time);
            end
            begin
              @(final_operation[19][23]) ;
              //$display("@%0t LEE: Received final operation event for 19,23\n", $time);
            end
            begin
              @(final_operation[19][24]) ;
              //$display("@%0t LEE: Received final operation event for 19,24\n", $time);
            end
            begin
              @(final_operation[19][25]) ;
              //$display("@%0t LEE: Received final operation event for 19,25\n", $time);
            end
            begin
              @(final_operation[19][26]) ;
              //$display("@%0t LEE: Received final operation event for 19,26\n", $time);
            end
            begin
              @(final_operation[19][27]) ;
              //$display("@%0t LEE: Received final operation event for 19,27\n", $time);
            end
            begin
              @(final_operation[19][28]) ;
              //$display("@%0t LEE: Received final operation event for 19,28\n", $time);
            end
            begin
              @(final_operation[19][29]) ;
              //$display("@%0t LEE: Received final operation event for 19,29\n", $time);
            end
            begin
              @(final_operation[19][30]) ;
              //$display("@%0t LEE: Received final operation event for 19,30\n", $time);
            end
            begin
              @(final_operation[19][31]) ;
              //$display("@%0t LEE: Received final operation event for 19,31\n", $time);
            end

            begin
              @(final_operation[20][0]) ;
              //$display("@%0t LEE: Received final operation event for 20,0\n", $time);
            end
            begin
              @(final_operation[20][1]) ;
              //$display("@%0t LEE: Received final operation event for 20,1\n", $time);
            end
            begin
              @(final_operation[20][2]) ;
              //$display("@%0t LEE: Received final operation event for 20,2\n", $time);
            end
            begin
              @(final_operation[20][3]) ;
              //$display("@%0t LEE: Received final operation event for 20,3\n", $time);
            end
            begin
              @(final_operation[20][4]) ;
              //$display("@%0t LEE: Received final operation event for 20,4\n", $time);
            end
            begin
              @(final_operation[20][5]) ;
              //$display("@%0t LEE: Received final operation event for 20,5\n", $time);
            end
            begin
              @(final_operation[20][6]) ;
              //$display("@%0t LEE: Received final operation event for 20,6\n", $time);
            end
            begin
              @(final_operation[20][7]) ;
              //$display("@%0t LEE: Received final operation event for 20,7\n", $time);
            end
            begin
              @(final_operation[20][8]) ;
              //$display("@%0t LEE: Received final operation event for 20,8\n", $time);
            end
            begin
              @(final_operation[20][9]) ;
              //$display("@%0t LEE: Received final operation event for 20,9\n", $time);
            end
            begin
              @(final_operation[20][10]) ;
              //$display("@%0t LEE: Received final operation event for 20,10\n", $time);
            end
            begin
              @(final_operation[20][11]) ;
              //$display("@%0t LEE: Received final operation event for 20,11\n", $time);
            end
            begin
              @(final_operation[20][12]) ;
              //$display("@%0t LEE: Received final operation event for 20,12\n", $time);
            end
            begin
              @(final_operation[20][13]) ;
              //$display("@%0t LEE: Received final operation event for 20,13\n", $time);
            end
            begin
              @(final_operation[20][14]) ;
              //$display("@%0t LEE: Received final operation event for 20,14\n", $time);
            end
            begin
              @(final_operation[20][15]) ;
              //$display("@%0t LEE: Received final operation event for 20,15\n", $time);
            end
            begin
              @(final_operation[20][16]) ;
              //$display("@%0t LEE: Received final operation event for 20,16\n", $time);
            end
            begin
              @(final_operation[20][17]) ;
              //$display("@%0t LEE: Received final operation event for 20,17\n", $time);
            end
            begin
              @(final_operation[20][18]) ;
              //$display("@%0t LEE: Received final operation event for 20,18\n", $time);
            end
            begin
              @(final_operation[20][19]) ;
              //$display("@%0t LEE: Received final operation event for 20,19\n", $time);
            end
            begin
              @(final_operation[20][20]) ;
              //$display("@%0t LEE: Received final operation event for 20,20\n", $time);
            end
            begin
              @(final_operation[20][21]) ;
              //$display("@%0t LEE: Received final operation event for 20,21\n", $time);
            end
            begin
              @(final_operation[20][22]) ;
              //$display("@%0t LEE: Received final operation event for 20,22\n", $time);
            end
            begin
              @(final_operation[20][23]) ;
              //$display("@%0t LEE: Received final operation event for 20,23\n", $time);
            end
            begin
              @(final_operation[20][24]) ;
              //$display("@%0t LEE: Received final operation event for 20,24\n", $time);
            end
            begin
              @(final_operation[20][25]) ;
              //$display("@%0t LEE: Received final operation event for 20,25\n", $time);
            end
            begin
              @(final_operation[20][26]) ;
              //$display("@%0t LEE: Received final operation event for 20,26\n", $time);
            end
            begin
              @(final_operation[20][27]) ;
              //$display("@%0t LEE: Received final operation event for 20,27\n", $time);
            end
            begin
              @(final_operation[20][28]) ;
              //$display("@%0t LEE: Received final operation event for 20,28\n", $time);
            end
            begin
              @(final_operation[20][29]) ;
              //$display("@%0t LEE: Received final operation event for 20,29\n", $time);
            end
            begin
              @(final_operation[20][30]) ;
              //$display("@%0t LEE: Received final operation event for 20,30\n", $time);
            end
            begin
              @(final_operation[20][31]) ;
              //$display("@%0t LEE: Received final operation event for 20,31\n", $time);
            end

            begin
              @(final_operation[21][0]) ;
              //$display("@%0t LEE: Received final operation event for 21,0\n", $time);
            end
            begin
              @(final_operation[21][1]) ;
              //$display("@%0t LEE: Received final operation event for 21,1\n", $time);
            end
            begin
              @(final_operation[21][2]) ;
              //$display("@%0t LEE: Received final operation event for 21,2\n", $time);
            end
            begin
              @(final_operation[21][3]) ;
              //$display("@%0t LEE: Received final operation event for 21,3\n", $time);
            end
            begin
              @(final_operation[21][4]) ;
              //$display("@%0t LEE: Received final operation event for 21,4\n", $time);
            end
            begin
              @(final_operation[21][5]) ;
              //$display("@%0t LEE: Received final operation event for 21,5\n", $time);
            end
            begin
              @(final_operation[21][6]) ;
              //$display("@%0t LEE: Received final operation event for 21,6\n", $time);
            end
            begin
              @(final_operation[21][7]) ;
              //$display("@%0t LEE: Received final operation event for 21,7\n", $time);
            end
            begin
              @(final_operation[21][8]) ;
              //$display("@%0t LEE: Received final operation event for 21,8\n", $time);
            end
            begin
              @(final_operation[21][9]) ;
              //$display("@%0t LEE: Received final operation event for 21,9\n", $time);
            end
            begin
              @(final_operation[21][10]) ;
              //$display("@%0t LEE: Received final operation event for 21,10\n", $time);
            end
            begin
              @(final_operation[21][11]) ;
              //$display("@%0t LEE: Received final operation event for 21,11\n", $time);
            end
            begin
              @(final_operation[21][12]) ;
              //$display("@%0t LEE: Received final operation event for 21,12\n", $time);
            end
            begin
              @(final_operation[21][13]) ;
              //$display("@%0t LEE: Received final operation event for 21,13\n", $time);
            end
            begin
              @(final_operation[21][14]) ;
              //$display("@%0t LEE: Received final operation event for 21,14\n", $time);
            end
            begin
              @(final_operation[21][15]) ;
              //$display("@%0t LEE: Received final operation event for 21,15\n", $time);
            end
            begin
              @(final_operation[21][16]) ;
              //$display("@%0t LEE: Received final operation event for 21,16\n", $time);
            end
            begin
              @(final_operation[21][17]) ;
              //$display("@%0t LEE: Received final operation event for 21,17\n", $time);
            end
            begin
              @(final_operation[21][18]) ;
              //$display("@%0t LEE: Received final operation event for 21,18\n", $time);
            end
            begin
              @(final_operation[21][19]) ;
              //$display("@%0t LEE: Received final operation event for 21,19\n", $time);
            end
            begin
              @(final_operation[21][20]) ;
              //$display("@%0t LEE: Received final operation event for 21,20\n", $time);
            end
            begin
              @(final_operation[21][21]) ;
              //$display("@%0t LEE: Received final operation event for 21,21\n", $time);
            end
            begin
              @(final_operation[21][22]) ;
              //$display("@%0t LEE: Received final operation event for 21,22\n", $time);
            end
            begin
              @(final_operation[21][23]) ;
              //$display("@%0t LEE: Received final operation event for 21,23\n", $time);
            end
            begin
              @(final_operation[21][24]) ;
              //$display("@%0t LEE: Received final operation event for 21,24\n", $time);
            end
            begin
              @(final_operation[21][25]) ;
              //$display("@%0t LEE: Received final operation event for 21,25\n", $time);
            end
            begin
              @(final_operation[21][26]) ;
              //$display("@%0t LEE: Received final operation event for 21,26\n", $time);
            end
            begin
              @(final_operation[21][27]) ;
              //$display("@%0t LEE: Received final operation event for 21,27\n", $time);
            end
            begin
              @(final_operation[21][28]) ;
              //$display("@%0t LEE: Received final operation event for 21,28\n", $time);
            end
            begin
              @(final_operation[21][29]) ;
              //$display("@%0t LEE: Received final operation event for 21,29\n", $time);
            end
            begin
              @(final_operation[21][30]) ;
              //$display("@%0t LEE: Received final operation event for 21,30\n", $time);
            end
            begin
              @(final_operation[21][31]) ;
              //$display("@%0t LEE: Received final operation event for 21,31\n", $time);
            end

            begin
              @(final_operation[22][0]) ;
              //$display("@%0t LEE: Received final operation event for 22,0\n", $time);
            end
            begin
              @(final_operation[22][1]) ;
              //$display("@%0t LEE: Received final operation event for 22,1\n", $time);
            end
            begin
              @(final_operation[22][2]) ;
              //$display("@%0t LEE: Received final operation event for 22,2\n", $time);
            end
            begin
              @(final_operation[22][3]) ;
              //$display("@%0t LEE: Received final operation event for 22,3\n", $time);
            end
            begin
              @(final_operation[22][4]) ;
              //$display("@%0t LEE: Received final operation event for 22,4\n", $time);
            end
            begin
              @(final_operation[22][5]) ;
              //$display("@%0t LEE: Received final operation event for 22,5\n", $time);
            end
            begin
              @(final_operation[22][6]) ;
              //$display("@%0t LEE: Received final operation event for 22,6\n", $time);
            end
            begin
              @(final_operation[22][7]) ;
              //$display("@%0t LEE: Received final operation event for 22,7\n", $time);
            end
            begin
              @(final_operation[22][8]) ;
              //$display("@%0t LEE: Received final operation event for 22,8\n", $time);
            end
            begin
              @(final_operation[22][9]) ;
              //$display("@%0t LEE: Received final operation event for 22,9\n", $time);
            end
            begin
              @(final_operation[22][10]) ;
              //$display("@%0t LEE: Received final operation event for 22,10\n", $time);
            end
            begin
              @(final_operation[22][11]) ;
              //$display("@%0t LEE: Received final operation event for 22,11\n", $time);
            end
            begin
              @(final_operation[22][12]) ;
              //$display("@%0t LEE: Received final operation event for 22,12\n", $time);
            end
            begin
              @(final_operation[22][13]) ;
              //$display("@%0t LEE: Received final operation event for 22,13\n", $time);
            end
            begin
              @(final_operation[22][14]) ;
              //$display("@%0t LEE: Received final operation event for 22,14\n", $time);
            end
            begin
              @(final_operation[22][15]) ;
              //$display("@%0t LEE: Received final operation event for 22,15\n", $time);
            end
            begin
              @(final_operation[22][16]) ;
              //$display("@%0t LEE: Received final operation event for 22,16\n", $time);
            end
            begin
              @(final_operation[22][17]) ;
              //$display("@%0t LEE: Received final operation event for 22,17\n", $time);
            end
            begin
              @(final_operation[22][18]) ;
              //$display("@%0t LEE: Received final operation event for 22,18\n", $time);
            end
            begin
              @(final_operation[22][19]) ;
              //$display("@%0t LEE: Received final operation event for 22,19\n", $time);
            end
            begin
              @(final_operation[22][20]) ;
              //$display("@%0t LEE: Received final operation event for 22,20\n", $time);
            end
            begin
              @(final_operation[22][21]) ;
              //$display("@%0t LEE: Received final operation event for 22,21\n", $time);
            end
            begin
              @(final_operation[22][22]) ;
              //$display("@%0t LEE: Received final operation event for 22,22\n", $time);
            end
            begin
              @(final_operation[22][23]) ;
              //$display("@%0t LEE: Received final operation event for 22,23\n", $time);
            end
            begin
              @(final_operation[22][24]) ;
              //$display("@%0t LEE: Received final operation event for 22,24\n", $time);
            end
            begin
              @(final_operation[22][25]) ;
              //$display("@%0t LEE: Received final operation event for 22,25\n", $time);
            end
            begin
              @(final_operation[22][26]) ;
              //$display("@%0t LEE: Received final operation event for 22,26\n", $time);
            end
            begin
              @(final_operation[22][27]) ;
              //$display("@%0t LEE: Received final operation event for 22,27\n", $time);
            end
            begin
              @(final_operation[22][28]) ;
              //$display("@%0t LEE: Received final operation event for 22,28\n", $time);
            end
            begin
              @(final_operation[22][29]) ;
              //$display("@%0t LEE: Received final operation event for 22,29\n", $time);
            end
            begin
              @(final_operation[22][30]) ;
              //$display("@%0t LEE: Received final operation event for 22,30\n", $time);
            end
            begin
              @(final_operation[22][31]) ;
              //$display("@%0t LEE: Received final operation event for 22,31\n", $time);
            end

            begin
              @(final_operation[23][0]) ;
              //$display("@%0t LEE: Received final operation event for 23,0\n", $time);
            end
            begin
              @(final_operation[23][1]) ;
              //$display("@%0t LEE: Received final operation event for 23,1\n", $time);
            end
            begin
              @(final_operation[23][2]) ;
              //$display("@%0t LEE: Received final operation event for 23,2\n", $time);
            end
            begin
              @(final_operation[23][3]) ;
              //$display("@%0t LEE: Received final operation event for 23,3\n", $time);
            end
            begin
              @(final_operation[23][4]) ;
              //$display("@%0t LEE: Received final operation event for 23,4\n", $time);
            end
            begin
              @(final_operation[23][5]) ;
              //$display("@%0t LEE: Received final operation event for 23,5\n", $time);
            end
            begin
              @(final_operation[23][6]) ;
              //$display("@%0t LEE: Received final operation event for 23,6\n", $time);
            end
            begin
              @(final_operation[23][7]) ;
              //$display("@%0t LEE: Received final operation event for 23,7\n", $time);
            end
            begin
              @(final_operation[23][8]) ;
              //$display("@%0t LEE: Received final operation event for 23,8\n", $time);
            end
            begin
              @(final_operation[23][9]) ;
              //$display("@%0t LEE: Received final operation event for 23,9\n", $time);
            end
            begin
              @(final_operation[23][10]) ;
              //$display("@%0t LEE: Received final operation event for 23,10\n", $time);
            end
            begin
              @(final_operation[23][11]) ;
              //$display("@%0t LEE: Received final operation event for 23,11\n", $time);
            end
            begin
              @(final_operation[23][12]) ;
              //$display("@%0t LEE: Received final operation event for 23,12\n", $time);
            end
            begin
              @(final_operation[23][13]) ;
              //$display("@%0t LEE: Received final operation event for 23,13\n", $time);
            end
            begin
              @(final_operation[23][14]) ;
              //$display("@%0t LEE: Received final operation event for 23,14\n", $time);
            end
            begin
              @(final_operation[23][15]) ;
              //$display("@%0t LEE: Received final operation event for 23,15\n", $time);
            end
            begin
              @(final_operation[23][16]) ;
              //$display("@%0t LEE: Received final operation event for 23,16\n", $time);
            end
            begin
              @(final_operation[23][17]) ;
              //$display("@%0t LEE: Received final operation event for 23,17\n", $time);
            end
            begin
              @(final_operation[23][18]) ;
              //$display("@%0t LEE: Received final operation event for 23,18\n", $time);
            end
            begin
              @(final_operation[23][19]) ;
              //$display("@%0t LEE: Received final operation event for 23,19\n", $time);
            end
            begin
              @(final_operation[23][20]) ;
              //$display("@%0t LEE: Received final operation event for 23,20\n", $time);
            end
            begin
              @(final_operation[23][21]) ;
              //$display("@%0t LEE: Received final operation event for 23,21\n", $time);
            end
            begin
              @(final_operation[23][22]) ;
              //$display("@%0t LEE: Received final operation event for 23,22\n", $time);
            end
            begin
              @(final_operation[23][23]) ;
              //$display("@%0t LEE: Received final operation event for 23,23\n", $time);
            end
            begin
              @(final_operation[23][24]) ;
              //$display("@%0t LEE: Received final operation event for 23,24\n", $time);
            end
            begin
              @(final_operation[23][25]) ;
              //$display("@%0t LEE: Received final operation event for 23,25\n", $time);
            end
            begin
              @(final_operation[23][26]) ;
              //$display("@%0t LEE: Received final operation event for 23,26\n", $time);
            end
            begin
              @(final_operation[23][27]) ;
              //$display("@%0t LEE: Received final operation event for 23,27\n", $time);
            end
            begin
              @(final_operation[23][28]) ;
              //$display("@%0t LEE: Received final operation event for 23,28\n", $time);
            end
            begin
              @(final_operation[23][29]) ;
              //$display("@%0t LEE: Received final operation event for 23,29\n", $time);
            end
            begin
              @(final_operation[23][30]) ;
              //$display("@%0t LEE: Received final operation event for 23,30\n", $time);
            end
            begin
              @(final_operation[23][31]) ;
              //$display("@%0t LEE: Received final operation event for 23,31\n", $time);
            end

            begin
              @(final_operation[24][0]) ;
              //$display("@%0t LEE: Received final operation event for 24,0\n", $time);
            end
            begin
              @(final_operation[24][1]) ;
              //$display("@%0t LEE: Received final operation event for 24,1\n", $time);
            end
            begin
              @(final_operation[24][2]) ;
              //$display("@%0t LEE: Received final operation event for 24,2\n", $time);
            end
            begin
              @(final_operation[24][3]) ;
              //$display("@%0t LEE: Received final operation event for 24,3\n", $time);
            end
            begin
              @(final_operation[24][4]) ;
              //$display("@%0t LEE: Received final operation event for 24,4\n", $time);
            end
            begin
              @(final_operation[24][5]) ;
              //$display("@%0t LEE: Received final operation event for 24,5\n", $time);
            end
            begin
              @(final_operation[24][6]) ;
              //$display("@%0t LEE: Received final operation event for 24,6\n", $time);
            end
            begin
              @(final_operation[24][7]) ;
              //$display("@%0t LEE: Received final operation event for 24,7\n", $time);
            end
            begin
              @(final_operation[24][8]) ;
              //$display("@%0t LEE: Received final operation event for 24,8\n", $time);
            end
            begin
              @(final_operation[24][9]) ;
              //$display("@%0t LEE: Received final operation event for 24,9\n", $time);
            end
            begin
              @(final_operation[24][10]) ;
              //$display("@%0t LEE: Received final operation event for 24,10\n", $time);
            end
            begin
              @(final_operation[24][11]) ;
              //$display("@%0t LEE: Received final operation event for 24,11\n", $time);
            end
            begin
              @(final_operation[24][12]) ;
              //$display("@%0t LEE: Received final operation event for 24,12\n", $time);
            end
            begin
              @(final_operation[24][13]) ;
              //$display("@%0t LEE: Received final operation event for 24,13\n", $time);
            end
            begin
              @(final_operation[24][14]) ;
              //$display("@%0t LEE: Received final operation event for 24,14\n", $time);
            end
            begin
              @(final_operation[24][15]) ;
              //$display("@%0t LEE: Received final operation event for 24,15\n", $time);
            end
            begin
              @(final_operation[24][16]) ;
              //$display("@%0t LEE: Received final operation event for 24,16\n", $time);
            end
            begin
              @(final_operation[24][17]) ;
              //$display("@%0t LEE: Received final operation event for 24,17\n", $time);
            end
            begin
              @(final_operation[24][18]) ;
              //$display("@%0t LEE: Received final operation event for 24,18\n", $time);
            end
            begin
              @(final_operation[24][19]) ;
              //$display("@%0t LEE: Received final operation event for 24,19\n", $time);
            end
            begin
              @(final_operation[24][20]) ;
              //$display("@%0t LEE: Received final operation event for 24,20\n", $time);
            end
            begin
              @(final_operation[24][21]) ;
              //$display("@%0t LEE: Received final operation event for 24,21\n", $time);
            end
            begin
              @(final_operation[24][22]) ;
              //$display("@%0t LEE: Received final operation event for 24,22\n", $time);
            end
            begin
              @(final_operation[24][23]) ;
              //$display("@%0t LEE: Received final operation event for 24,23\n", $time);
            end
            begin
              @(final_operation[24][24]) ;
              //$display("@%0t LEE: Received final operation event for 24,24\n", $time);
            end
            begin
              @(final_operation[24][25]) ;
              //$display("@%0t LEE: Received final operation event for 24,25\n", $time);
            end
            begin
              @(final_operation[24][26]) ;
              //$display("@%0t LEE: Received final operation event for 24,26\n", $time);
            end
            begin
              @(final_operation[24][27]) ;
              //$display("@%0t LEE: Received final operation event for 24,27\n", $time);
            end
            begin
              @(final_operation[24][28]) ;
              //$display("@%0t LEE: Received final operation event for 24,28\n", $time);
            end
            begin
              @(final_operation[24][29]) ;
              //$display("@%0t LEE: Received final operation event for 24,29\n", $time);
            end
            begin
              @(final_operation[24][30]) ;
              //$display("@%0t LEE: Received final operation event for 24,30\n", $time);
            end
            begin
              @(final_operation[24][31]) ;
              //$display("@%0t LEE: Received final operation event for 24,31\n", $time);
            end

            begin
              @(final_operation[25][0]) ;
              //$display("@%0t LEE: Received final operation event for 25,0\n", $time);
            end
            begin
              @(final_operation[25][1]) ;
              //$display("@%0t LEE: Received final operation event for 25,1\n", $time);
            end
            begin
              @(final_operation[25][2]) ;
              //$display("@%0t LEE: Received final operation event for 25,2\n", $time);
            end
            begin
              @(final_operation[25][3]) ;
              //$display("@%0t LEE: Received final operation event for 25,3\n", $time);
            end
            begin
              @(final_operation[25][4]) ;
              //$display("@%0t LEE: Received final operation event for 25,4\n", $time);
            end
            begin
              @(final_operation[25][5]) ;
              //$display("@%0t LEE: Received final operation event for 25,5\n", $time);
            end
            begin
              @(final_operation[25][6]) ;
              //$display("@%0t LEE: Received final operation event for 25,6\n", $time);
            end
            begin
              @(final_operation[25][7]) ;
              //$display("@%0t LEE: Received final operation event for 25,7\n", $time);
            end
            begin
              @(final_operation[25][8]) ;
              //$display("@%0t LEE: Received final operation event for 25,8\n", $time);
            end
            begin
              @(final_operation[25][9]) ;
              //$display("@%0t LEE: Received final operation event for 25,9\n", $time);
            end
            begin
              @(final_operation[25][10]) ;
              //$display("@%0t LEE: Received final operation event for 25,10\n", $time);
            end
            begin
              @(final_operation[25][11]) ;
              //$display("@%0t LEE: Received final operation event for 25,11\n", $time);
            end
            begin
              @(final_operation[25][12]) ;
              //$display("@%0t LEE: Received final operation event for 25,12\n", $time);
            end
            begin
              @(final_operation[25][13]) ;
              //$display("@%0t LEE: Received final operation event for 25,13\n", $time);
            end
            begin
              @(final_operation[25][14]) ;
              //$display("@%0t LEE: Received final operation event for 25,14\n", $time);
            end
            begin
              @(final_operation[25][15]) ;
              //$display("@%0t LEE: Received final operation event for 25,15\n", $time);
            end
            begin
              @(final_operation[25][16]) ;
              //$display("@%0t LEE: Received final operation event for 25,16\n", $time);
            end
            begin
              @(final_operation[25][17]) ;
              //$display("@%0t LEE: Received final operation event for 25,17\n", $time);
            end
            begin
              @(final_operation[25][18]) ;
              //$display("@%0t LEE: Received final operation event for 25,18\n", $time);
            end
            begin
              @(final_operation[25][19]) ;
              //$display("@%0t LEE: Received final operation event for 25,19\n", $time);
            end
            begin
              @(final_operation[25][20]) ;
              //$display("@%0t LEE: Received final operation event for 25,20\n", $time);
            end
            begin
              @(final_operation[25][21]) ;
              //$display("@%0t LEE: Received final operation event for 25,21\n", $time);
            end
            begin
              @(final_operation[25][22]) ;
              //$display("@%0t LEE: Received final operation event for 25,22\n", $time);
            end
            begin
              @(final_operation[25][23]) ;
              //$display("@%0t LEE: Received final operation event for 25,23\n", $time);
            end
            begin
              @(final_operation[25][24]) ;
              //$display("@%0t LEE: Received final operation event for 25,24\n", $time);
            end
            begin
              @(final_operation[25][25]) ;
              //$display("@%0t LEE: Received final operation event for 25,25\n", $time);
            end
            begin
              @(final_operation[25][26]) ;
              //$display("@%0t LEE: Received final operation event for 25,26\n", $time);
            end
            begin
              @(final_operation[25][27]) ;
              //$display("@%0t LEE: Received final operation event for 25,27\n", $time);
            end
            begin
              @(final_operation[25][28]) ;
              //$display("@%0t LEE: Received final operation event for 25,28\n", $time);
            end
            begin
              @(final_operation[25][29]) ;
              //$display("@%0t LEE: Received final operation event for 25,29\n", $time);
            end
            begin
              @(final_operation[25][30]) ;
              //$display("@%0t LEE: Received final operation event for 25,30\n", $time);
            end
            begin
              @(final_operation[25][31]) ;
              //$display("@%0t LEE: Received final operation event for 25,31\n", $time);
            end

            begin
              @(final_operation[26][0]) ;
              //$display("@%0t LEE: Received final operation event for 26,0\n", $time);
            end
            begin
              @(final_operation[26][1]) ;
              //$display("@%0t LEE: Received final operation event for 26,1\n", $time);
            end
            begin
              @(final_operation[26][2]) ;
              //$display("@%0t LEE: Received final operation event for 26,2\n", $time);
            end
            begin
              @(final_operation[26][3]) ;
              //$display("@%0t LEE: Received final operation event for 26,3\n", $time);
            end
            begin
              @(final_operation[26][4]) ;
              //$display("@%0t LEE: Received final operation event for 26,4\n", $time);
            end
            begin
              @(final_operation[26][5]) ;
              //$display("@%0t LEE: Received final operation event for 26,5\n", $time);
            end
            begin
              @(final_operation[26][6]) ;
              //$display("@%0t LEE: Received final operation event for 26,6\n", $time);
            end
            begin
              @(final_operation[26][7]) ;
              //$display("@%0t LEE: Received final operation event for 26,7\n", $time);
            end
            begin
              @(final_operation[26][8]) ;
              //$display("@%0t LEE: Received final operation event for 26,8\n", $time);
            end
            begin
              @(final_operation[26][9]) ;
              //$display("@%0t LEE: Received final operation event for 26,9\n", $time);
            end
            begin
              @(final_operation[26][10]) ;
              //$display("@%0t LEE: Received final operation event for 26,10\n", $time);
            end
            begin
              @(final_operation[26][11]) ;
              //$display("@%0t LEE: Received final operation event for 26,11\n", $time);
            end
            begin
              @(final_operation[26][12]) ;
              //$display("@%0t LEE: Received final operation event for 26,12\n", $time);
            end
            begin
              @(final_operation[26][13]) ;
              //$display("@%0t LEE: Received final operation event for 26,13\n", $time);
            end
            begin
              @(final_operation[26][14]) ;
              //$display("@%0t LEE: Received final operation event for 26,14\n", $time);
            end
            begin
              @(final_operation[26][15]) ;
              //$display("@%0t LEE: Received final operation event for 26,15\n", $time);
            end
            begin
              @(final_operation[26][16]) ;
              //$display("@%0t LEE: Received final operation event for 26,16\n", $time);
            end
            begin
              @(final_operation[26][17]) ;
              //$display("@%0t LEE: Received final operation event for 26,17\n", $time);
            end
            begin
              @(final_operation[26][18]) ;
              //$display("@%0t LEE: Received final operation event for 26,18\n", $time);
            end
            begin
              @(final_operation[26][19]) ;
              //$display("@%0t LEE: Received final operation event for 26,19\n", $time);
            end
            begin
              @(final_operation[26][20]) ;
              //$display("@%0t LEE: Received final operation event for 26,20\n", $time);
            end
            begin
              @(final_operation[26][21]) ;
              //$display("@%0t LEE: Received final operation event for 26,21\n", $time);
            end
            begin
              @(final_operation[26][22]) ;
              //$display("@%0t LEE: Received final operation event for 26,22\n", $time);
            end
            begin
              @(final_operation[26][23]) ;
              //$display("@%0t LEE: Received final operation event for 26,23\n", $time);
            end
            begin
              @(final_operation[26][24]) ;
              //$display("@%0t LEE: Received final operation event for 26,24\n", $time);
            end
            begin
              @(final_operation[26][25]) ;
              //$display("@%0t LEE: Received final operation event for 26,25\n", $time);
            end
            begin
              @(final_operation[26][26]) ;
              //$display("@%0t LEE: Received final operation event for 26,26\n", $time);
            end
            begin
              @(final_operation[26][27]) ;
              //$display("@%0t LEE: Received final operation event for 26,27\n", $time);
            end
            begin
              @(final_operation[26][28]) ;
              //$display("@%0t LEE: Received final operation event for 26,28\n", $time);
            end
            begin
              @(final_operation[26][29]) ;
              //$display("@%0t LEE: Received final operation event for 26,29\n", $time);
            end
            begin
              @(final_operation[26][30]) ;
              //$display("@%0t LEE: Received final operation event for 26,30\n", $time);
            end
            begin
              @(final_operation[26][31]) ;
              //$display("@%0t LEE: Received final operation event for 26,31\n", $time);
            end

            begin
              @(final_operation[27][0]) ;
              //$display("@%0t LEE: Received final operation event for 27,0\n", $time);
            end
            begin
              @(final_operation[27][1]) ;
              //$display("@%0t LEE: Received final operation event for 27,1\n", $time);
            end
            begin
              @(final_operation[27][2]) ;
              //$display("@%0t LEE: Received final operation event for 27,2\n", $time);
            end
            begin
              @(final_operation[27][3]) ;
              //$display("@%0t LEE: Received final operation event for 27,3\n", $time);
            end
            begin
              @(final_operation[27][4]) ;
              //$display("@%0t LEE: Received final operation event for 27,4\n", $time);
            end
            begin
              @(final_operation[27][5]) ;
              //$display("@%0t LEE: Received final operation event for 27,5\n", $time);
            end
            begin
              @(final_operation[27][6]) ;
              //$display("@%0t LEE: Received final operation event for 27,6\n", $time);
            end
            begin
              @(final_operation[27][7]) ;
              //$display("@%0t LEE: Received final operation event for 27,7\n", $time);
            end
            begin
              @(final_operation[27][8]) ;
              //$display("@%0t LEE: Received final operation event for 27,8\n", $time);
            end
            begin
              @(final_operation[27][9]) ;
              //$display("@%0t LEE: Received final operation event for 27,9\n", $time);
            end
            begin
              @(final_operation[27][10]) ;
              //$display("@%0t LEE: Received final operation event for 27,10\n", $time);
            end
            begin
              @(final_operation[27][11]) ;
              //$display("@%0t LEE: Received final operation event for 27,11\n", $time);
            end
            begin
              @(final_operation[27][12]) ;
              //$display("@%0t LEE: Received final operation event for 27,12\n", $time);
            end
            begin
              @(final_operation[27][13]) ;
              //$display("@%0t LEE: Received final operation event for 27,13\n", $time);
            end
            begin
              @(final_operation[27][14]) ;
              //$display("@%0t LEE: Received final operation event for 27,14\n", $time);
            end
            begin
              @(final_operation[27][15]) ;
              //$display("@%0t LEE: Received final operation event for 27,15\n", $time);
            end
            begin
              @(final_operation[27][16]) ;
              //$display("@%0t LEE: Received final operation event for 27,16\n", $time);
            end
            begin
              @(final_operation[27][17]) ;
              //$display("@%0t LEE: Received final operation event for 27,17\n", $time);
            end
            begin
              @(final_operation[27][18]) ;
              //$display("@%0t LEE: Received final operation event for 27,18\n", $time);
            end
            begin
              @(final_operation[27][19]) ;
              //$display("@%0t LEE: Received final operation event for 27,19\n", $time);
            end
            begin
              @(final_operation[27][20]) ;
              //$display("@%0t LEE: Received final operation event for 27,20\n", $time);
            end
            begin
              @(final_operation[27][21]) ;
              //$display("@%0t LEE: Received final operation event for 27,21\n", $time);
            end
            begin
              @(final_operation[27][22]) ;
              //$display("@%0t LEE: Received final operation event for 27,22\n", $time);
            end
            begin
              @(final_operation[27][23]) ;
              //$display("@%0t LEE: Received final operation event for 27,23\n", $time);
            end
            begin
              @(final_operation[27][24]) ;
              //$display("@%0t LEE: Received final operation event for 27,24\n", $time);
            end
            begin
              @(final_operation[27][25]) ;
              //$display("@%0t LEE: Received final operation event for 27,25\n", $time);
            end
            begin
              @(final_operation[27][26]) ;
              //$display("@%0t LEE: Received final operation event for 27,26\n", $time);
            end
            begin
              @(final_operation[27][27]) ;
              //$display("@%0t LEE: Received final operation event for 27,27\n", $time);
            end
            begin
              @(final_operation[27][28]) ;
              //$display("@%0t LEE: Received final operation event for 27,28\n", $time);
            end
            begin
              @(final_operation[27][29]) ;
              //$display("@%0t LEE: Received final operation event for 27,29\n", $time);
            end
            begin
              @(final_operation[27][30]) ;
              //$display("@%0t LEE: Received final operation event for 27,30\n", $time);
            end
            begin
              @(final_operation[27][31]) ;
              //$display("@%0t LEE: Received final operation event for 27,31\n", $time);
            end

            begin
              @(final_operation[28][0]) ;
              //$display("@%0t LEE: Received final operation event for 28,0\n", $time);
            end
            begin
              @(final_operation[28][1]) ;
              //$display("@%0t LEE: Received final operation event for 28,1\n", $time);
            end
            begin
              @(final_operation[28][2]) ;
              //$display("@%0t LEE: Received final operation event for 28,2\n", $time);
            end
            begin
              @(final_operation[28][3]) ;
              //$display("@%0t LEE: Received final operation event for 28,3\n", $time);
            end
            begin
              @(final_operation[28][4]) ;
              //$display("@%0t LEE: Received final operation event for 28,4\n", $time);
            end
            begin
              @(final_operation[28][5]) ;
              //$display("@%0t LEE: Received final operation event for 28,5\n", $time);
            end
            begin
              @(final_operation[28][6]) ;
              //$display("@%0t LEE: Received final operation event for 28,6\n", $time);
            end
            begin
              @(final_operation[28][7]) ;
              //$display("@%0t LEE: Received final operation event for 28,7\n", $time);
            end
            begin
              @(final_operation[28][8]) ;
              //$display("@%0t LEE: Received final operation event for 28,8\n", $time);
            end
            begin
              @(final_operation[28][9]) ;
              //$display("@%0t LEE: Received final operation event for 28,9\n", $time);
            end
            begin
              @(final_operation[28][10]) ;
              //$display("@%0t LEE: Received final operation event for 28,10\n", $time);
            end
            begin
              @(final_operation[28][11]) ;
              //$display("@%0t LEE: Received final operation event for 28,11\n", $time);
            end
            begin
              @(final_operation[28][12]) ;
              //$display("@%0t LEE: Received final operation event for 28,12\n", $time);
            end
            begin
              @(final_operation[28][13]) ;
              //$display("@%0t LEE: Received final operation event for 28,13\n", $time);
            end
            begin
              @(final_operation[28][14]) ;
              //$display("@%0t LEE: Received final operation event for 28,14\n", $time);
            end
            begin
              @(final_operation[28][15]) ;
              //$display("@%0t LEE: Received final operation event for 28,15\n", $time);
            end
            begin
              @(final_operation[28][16]) ;
              //$display("@%0t LEE: Received final operation event for 28,16\n", $time);
            end
            begin
              @(final_operation[28][17]) ;
              //$display("@%0t LEE: Received final operation event for 28,17\n", $time);
            end
            begin
              @(final_operation[28][18]) ;
              //$display("@%0t LEE: Received final operation event for 28,18\n", $time);
            end
            begin
              @(final_operation[28][19]) ;
              //$display("@%0t LEE: Received final operation event for 28,19\n", $time);
            end
            begin
              @(final_operation[28][20]) ;
              //$display("@%0t LEE: Received final operation event for 28,20\n", $time);
            end
            begin
              @(final_operation[28][21]) ;
              //$display("@%0t LEE: Received final operation event for 28,21\n", $time);
            end
            begin
              @(final_operation[28][22]) ;
              //$display("@%0t LEE: Received final operation event for 28,22\n", $time);
            end
            begin
              @(final_operation[28][23]) ;
              //$display("@%0t LEE: Received final operation event for 28,23\n", $time);
            end
            begin
              @(final_operation[28][24]) ;
              //$display("@%0t LEE: Received final operation event for 28,24\n", $time);
            end
            begin
              @(final_operation[28][25]) ;
              //$display("@%0t LEE: Received final operation event for 28,25\n", $time);
            end
            begin
              @(final_operation[28][26]) ;
              //$display("@%0t LEE: Received final operation event for 28,26\n", $time);
            end
            begin
              @(final_operation[28][27]) ;
              //$display("@%0t LEE: Received final operation event for 28,27\n", $time);
            end
            begin
              @(final_operation[28][28]) ;
              //$display("@%0t LEE: Received final operation event for 28,28\n", $time);
            end
            begin
              @(final_operation[28][29]) ;
              //$display("@%0t LEE: Received final operation event for 28,29\n", $time);
            end
            begin
              @(final_operation[28][30]) ;
              //$display("@%0t LEE: Received final operation event for 28,30\n", $time);
            end
            begin
              @(final_operation[28][31]) ;
              //$display("@%0t LEE: Received final operation event for 28,31\n", $time);
            end

            begin
              @(final_operation[29][0]) ;
              //$display("@%0t LEE: Received final operation event for 29,0\n", $time);
            end
            begin
              @(final_operation[29][1]) ;
              //$display("@%0t LEE: Received final operation event for 29,1\n", $time);
            end
            begin
              @(final_operation[29][2]) ;
              //$display("@%0t LEE: Received final operation event for 29,2\n", $time);
            end
            begin
              @(final_operation[29][3]) ;
              //$display("@%0t LEE: Received final operation event for 29,3\n", $time);
            end
            begin
              @(final_operation[29][4]) ;
              //$display("@%0t LEE: Received final operation event for 29,4\n", $time);
            end
            begin
              @(final_operation[29][5]) ;
              //$display("@%0t LEE: Received final operation event for 29,5\n", $time);
            end
            begin
              @(final_operation[29][6]) ;
              //$display("@%0t LEE: Received final operation event for 29,6\n", $time);
            end
            begin
              @(final_operation[29][7]) ;
              //$display("@%0t LEE: Received final operation event for 29,7\n", $time);
            end
            begin
              @(final_operation[29][8]) ;
              //$display("@%0t LEE: Received final operation event for 29,8\n", $time);
            end
            begin
              @(final_operation[29][9]) ;
              //$display("@%0t LEE: Received final operation event for 29,9\n", $time);
            end
            begin
              @(final_operation[29][10]) ;
              //$display("@%0t LEE: Received final operation event for 29,10\n", $time);
            end
            begin
              @(final_operation[29][11]) ;
              //$display("@%0t LEE: Received final operation event for 29,11\n", $time);
            end
            begin
              @(final_operation[29][12]) ;
              //$display("@%0t LEE: Received final operation event for 29,12\n", $time);
            end
            begin
              @(final_operation[29][13]) ;
              //$display("@%0t LEE: Received final operation event for 29,13\n", $time);
            end
            begin
              @(final_operation[29][14]) ;
              //$display("@%0t LEE: Received final operation event for 29,14\n", $time);
            end
            begin
              @(final_operation[29][15]) ;
              //$display("@%0t LEE: Received final operation event for 29,15\n", $time);
            end
            begin
              @(final_operation[29][16]) ;
              //$display("@%0t LEE: Received final operation event for 29,16\n", $time);
            end
            begin
              @(final_operation[29][17]) ;
              //$display("@%0t LEE: Received final operation event for 29,17\n", $time);
            end
            begin
              @(final_operation[29][18]) ;
              //$display("@%0t LEE: Received final operation event for 29,18\n", $time);
            end
            begin
              @(final_operation[29][19]) ;
              //$display("@%0t LEE: Received final operation event for 29,19\n", $time);
            end
            begin
              @(final_operation[29][20]) ;
              //$display("@%0t LEE: Received final operation event for 29,20\n", $time);
            end
            begin
              @(final_operation[29][21]) ;
              //$display("@%0t LEE: Received final operation event for 29,21\n", $time);
            end
            begin
              @(final_operation[29][22]) ;
              //$display("@%0t LEE: Received final operation event for 29,22\n", $time);
            end
            begin
              @(final_operation[29][23]) ;
              //$display("@%0t LEE: Received final operation event for 29,23\n", $time);
            end
            begin
              @(final_operation[29][24]) ;
              //$display("@%0t LEE: Received final operation event for 29,24\n", $time);
            end
            begin
              @(final_operation[29][25]) ;
              //$display("@%0t LEE: Received final operation event for 29,25\n", $time);
            end
            begin
              @(final_operation[29][26]) ;
              //$display("@%0t LEE: Received final operation event for 29,26\n", $time);
            end
            begin
              @(final_operation[29][27]) ;
              //$display("@%0t LEE: Received final operation event for 29,27\n", $time);
            end
            begin
              @(final_operation[29][28]) ;
              //$display("@%0t LEE: Received final operation event for 29,28\n", $time);
            end
            begin
              @(final_operation[29][29]) ;
              //$display("@%0t LEE: Received final operation event for 29,29\n", $time);
            end
            begin
              @(final_operation[29][30]) ;
              //$display("@%0t LEE: Received final operation event for 29,30\n", $time);
            end
            begin
              @(final_operation[29][31]) ;
              //$display("@%0t LEE: Received final operation event for 29,31\n", $time);
            end

            begin
              @(final_operation[30][0]) ;
              //$display("@%0t LEE: Received final operation event for 30,0\n", $time);
            end
            begin
              @(final_operation[30][1]) ;
              //$display("@%0t LEE: Received final operation event for 30,1\n", $time);
            end
            begin
              @(final_operation[30][2]) ;
              //$display("@%0t LEE: Received final operation event for 30,2\n", $time);
            end
            begin
              @(final_operation[30][3]) ;
              //$display("@%0t LEE: Received final operation event for 30,3\n", $time);
            end
            begin
              @(final_operation[30][4]) ;
              //$display("@%0t LEE: Received final operation event for 30,4\n", $time);
            end
            begin
              @(final_operation[30][5]) ;
              //$display("@%0t LEE: Received final operation event for 30,5\n", $time);
            end
            begin
              @(final_operation[30][6]) ;
              //$display("@%0t LEE: Received final operation event for 30,6\n", $time);
            end
            begin
              @(final_operation[30][7]) ;
              //$display("@%0t LEE: Received final operation event for 30,7\n", $time);
            end
            begin
              @(final_operation[30][8]) ;
              //$display("@%0t LEE: Received final operation event for 30,8\n", $time);
            end
            begin
              @(final_operation[30][9]) ;
              //$display("@%0t LEE: Received final operation event for 30,9\n", $time);
            end
            begin
              @(final_operation[30][10]) ;
              //$display("@%0t LEE: Received final operation event for 30,10\n", $time);
            end
            begin
              @(final_operation[30][11]) ;
              //$display("@%0t LEE: Received final operation event for 30,11\n", $time);
            end
            begin
              @(final_operation[30][12]) ;
              //$display("@%0t LEE: Received final operation event for 30,12\n", $time);
            end
            begin
              @(final_operation[30][13]) ;
              //$display("@%0t LEE: Received final operation event for 30,13\n", $time);
            end
            begin
              @(final_operation[30][14]) ;
              //$display("@%0t LEE: Received final operation event for 30,14\n", $time);
            end
            begin
              @(final_operation[30][15]) ;
              //$display("@%0t LEE: Received final operation event for 30,15\n", $time);
            end
            begin
              @(final_operation[30][16]) ;
              //$display("@%0t LEE: Received final operation event for 30,16\n", $time);
            end
            begin
              @(final_operation[30][17]) ;
              //$display("@%0t LEE: Received final operation event for 30,17\n", $time);
            end
            begin
              @(final_operation[30][18]) ;
              //$display("@%0t LEE: Received final operation event for 30,18\n", $time);
            end
            begin
              @(final_operation[30][19]) ;
              //$display("@%0t LEE: Received final operation event for 30,19\n", $time);
            end
            begin
              @(final_operation[30][20]) ;
              //$display("@%0t LEE: Received final operation event for 30,20\n", $time);
            end
            begin
              @(final_operation[30][21]) ;
              //$display("@%0t LEE: Received final operation event for 30,21\n", $time);
            end
            begin
              @(final_operation[30][22]) ;
              //$display("@%0t LEE: Received final operation event for 30,22\n", $time);
            end
            begin
              @(final_operation[30][23]) ;
              //$display("@%0t LEE: Received final operation event for 30,23\n", $time);
            end
            begin
              @(final_operation[30][24]) ;
              //$display("@%0t LEE: Received final operation event for 30,24\n", $time);
            end
            begin
              @(final_operation[30][25]) ;
              //$display("@%0t LEE: Received final operation event for 30,25\n", $time);
            end
            begin
              @(final_operation[30][26]) ;
              //$display("@%0t LEE: Received final operation event for 30,26\n", $time);
            end
            begin
              @(final_operation[30][27]) ;
              //$display("@%0t LEE: Received final operation event for 30,27\n", $time);
            end
            begin
              @(final_operation[30][28]) ;
              //$display("@%0t LEE: Received final operation event for 30,28\n", $time);
            end
            begin
              @(final_operation[30][29]) ;
              //$display("@%0t LEE: Received final operation event for 30,29\n", $time);
            end
            begin
              @(final_operation[30][30]) ;
              //$display("@%0t LEE: Received final operation event for 30,30\n", $time);
            end
            begin
              @(final_operation[30][31]) ;
              //$display("@%0t LEE: Received final operation event for 30,31\n", $time);
            end

            begin
              @(final_operation[31][0]) ;
              //$display("@%0t LEE: Received final operation event for 31,0\n", $time);
            end
            begin
              @(final_operation[31][1]) ;
              //$display("@%0t LEE: Received final operation event for 31,1\n", $time);
            end
            begin
              @(final_operation[31][2]) ;
              //$display("@%0t LEE: Received final operation event for 31,2\n", $time);
            end
            begin
              @(final_operation[31][3]) ;
              //$display("@%0t LEE: Received final operation event for 31,3\n", $time);
            end
            begin
              @(final_operation[31][4]) ;
              //$display("@%0t LEE: Received final operation event for 31,4\n", $time);
            end
            begin
              @(final_operation[31][5]) ;
              //$display("@%0t LEE: Received final operation event for 31,5\n", $time);
            end
            begin
              @(final_operation[31][6]) ;
              //$display("@%0t LEE: Received final operation event for 31,6\n", $time);
            end
            begin
              @(final_operation[31][7]) ;
              //$display("@%0t LEE: Received final operation event for 31,7\n", $time);
            end
            begin
              @(final_operation[31][8]) ;
              //$display("@%0t LEE: Received final operation event for 31,8\n", $time);
            end
            begin
              @(final_operation[31][9]) ;
              //$display("@%0t LEE: Received final operation event for 31,9\n", $time);
            end
            begin
              @(final_operation[31][10]) ;
              //$display("@%0t LEE: Received final operation event for 31,10\n", $time);
            end
            begin
              @(final_operation[31][11]) ;
              //$display("@%0t LEE: Received final operation event for 31,11\n", $time);
            end
            begin
              @(final_operation[31][12]) ;
              //$display("@%0t LEE: Received final operation event for 31,12\n", $time);
            end
            begin
              @(final_operation[31][13]) ;
              //$display("@%0t LEE: Received final operation event for 31,13\n", $time);
            end
            begin
              @(final_operation[31][14]) ;
              //$display("@%0t LEE: Received final operation event for 31,14\n", $time);
            end
            begin
              @(final_operation[31][15]) ;
              //$display("@%0t LEE: Received final operation event for 31,15\n", $time);
            end
            begin
              @(final_operation[31][16]) ;
              //$display("@%0t LEE: Received final operation event for 31,16\n", $time);
            end
            begin
              @(final_operation[31][17]) ;
              //$display("@%0t LEE: Received final operation event for 31,17\n", $time);
            end
            begin
              @(final_operation[31][18]) ;
              //$display("@%0t LEE: Received final operation event for 31,18\n", $time);
            end
            begin
              @(final_operation[31][19]) ;
              //$display("@%0t LEE: Received final operation event for 31,19\n", $time);
            end
            begin
              @(final_operation[31][20]) ;
              //$display("@%0t LEE: Received final operation event for 31,20\n", $time);
            end
            begin
              @(final_operation[31][21]) ;
              //$display("@%0t LEE: Received final operation event for 31,21\n", $time);
            end
            begin
              @(final_operation[31][22]) ;
              //$display("@%0t LEE: Received final operation event for 31,22\n", $time);
            end
            begin
              @(final_operation[31][23]) ;
              //$display("@%0t LEE: Received final operation event for 31,23\n", $time);
            end
            begin
              @(final_operation[31][24]) ;
              //$display("@%0t LEE: Received final operation event for 31,24\n", $time);
            end
            begin
              @(final_operation[31][25]) ;
              //$display("@%0t LEE: Received final operation event for 31,25\n", $time);
            end
            begin
              @(final_operation[31][26]) ;
              //$display("@%0t LEE: Received final operation event for 31,26\n", $time);
            end
            begin
              @(final_operation[31][27]) ;
              //$display("@%0t LEE: Received final operation event for 31,27\n", $time);
            end
            begin
              @(final_operation[31][28]) ;
              //$display("@%0t LEE: Received final operation event for 31,28\n", $time);
            end
            begin
              @(final_operation[31][29]) ;
              //$display("@%0t LEE: Received final operation event for 31,29\n", $time);
            end
            begin
              @(final_operation[31][30]) ;
              //$display("@%0t LEE: Received final operation event for 31,30\n", $time);
            end
            begin
              @(final_operation[31][31]) ;
              //$display("@%0t LEE: Received final operation event for 31,31\n", $time);
            end

            begin
              @(final_operation[32][0]) ;
              //$display("@%0t LEE: Received final operation event for 32,0\n", $time);
            end
            begin
              @(final_operation[32][1]) ;
              //$display("@%0t LEE: Received final operation event for 32,1\n", $time);
            end
            begin
              @(final_operation[32][2]) ;
              //$display("@%0t LEE: Received final operation event for 32,2\n", $time);
            end
            begin
              @(final_operation[32][3]) ;
              //$display("@%0t LEE: Received final operation event for 32,3\n", $time);
            end
            begin
              @(final_operation[32][4]) ;
              //$display("@%0t LEE: Received final operation event for 32,4\n", $time);
            end
            begin
              @(final_operation[32][5]) ;
              //$display("@%0t LEE: Received final operation event for 32,5\n", $time);
            end
            begin
              @(final_operation[32][6]) ;
              //$display("@%0t LEE: Received final operation event for 32,6\n", $time);
            end
            begin
              @(final_operation[32][7]) ;
              //$display("@%0t LEE: Received final operation event for 32,7\n", $time);
            end
            begin
              @(final_operation[32][8]) ;
              //$display("@%0t LEE: Received final operation event for 32,8\n", $time);
            end
            begin
              @(final_operation[32][9]) ;
              //$display("@%0t LEE: Received final operation event for 32,9\n", $time);
            end
            begin
              @(final_operation[32][10]) ;
              //$display("@%0t LEE: Received final operation event for 32,10\n", $time);
            end
            begin
              @(final_operation[32][11]) ;
              //$display("@%0t LEE: Received final operation event for 32,11\n", $time);
            end
            begin
              @(final_operation[32][12]) ;
              //$display("@%0t LEE: Received final operation event for 32,12\n", $time);
            end
            begin
              @(final_operation[32][13]) ;
              //$display("@%0t LEE: Received final operation event for 32,13\n", $time);
            end
            begin
              @(final_operation[32][14]) ;
              //$display("@%0t LEE: Received final operation event for 32,14\n", $time);
            end
            begin
              @(final_operation[32][15]) ;
              //$display("@%0t LEE: Received final operation event for 32,15\n", $time);
            end
            begin
              @(final_operation[32][16]) ;
              //$display("@%0t LEE: Received final operation event for 32,16\n", $time);
            end
            begin
              @(final_operation[32][17]) ;
              //$display("@%0t LEE: Received final operation event for 32,17\n", $time);
            end
            begin
              @(final_operation[32][18]) ;
              //$display("@%0t LEE: Received final operation event for 32,18\n", $time);
            end
            begin
              @(final_operation[32][19]) ;
              //$display("@%0t LEE: Received final operation event for 32,19\n", $time);
            end
            begin
              @(final_operation[32][20]) ;
              //$display("@%0t LEE: Received final operation event for 32,20\n", $time);
            end
            begin
              @(final_operation[32][21]) ;
              //$display("@%0t LEE: Received final operation event for 32,21\n", $time);
            end
            begin
              @(final_operation[32][22]) ;
              //$display("@%0t LEE: Received final operation event for 32,22\n", $time);
            end
            begin
              @(final_operation[32][23]) ;
              //$display("@%0t LEE: Received final operation event for 32,23\n", $time);
            end
            begin
              @(final_operation[32][24]) ;
              //$display("@%0t LEE: Received final operation event for 32,24\n", $time);
            end
            begin
              @(final_operation[32][25]) ;
              //$display("@%0t LEE: Received final operation event for 32,25\n", $time);
            end
            begin
              @(final_operation[32][26]) ;
              //$display("@%0t LEE: Received final operation event for 32,26\n", $time);
            end
            begin
              @(final_operation[32][27]) ;
              //$display("@%0t LEE: Received final operation event for 32,27\n", $time);
            end
            begin
              @(final_operation[32][28]) ;
              //$display("@%0t LEE: Received final operation event for 32,28\n", $time);
            end
            begin
              @(final_operation[32][29]) ;
              //$display("@%0t LEE: Received final operation event for 32,29\n", $time);
            end
            begin
              @(final_operation[32][30]) ;
              //$display("@%0t LEE: Received final operation event for 32,30\n", $time);
            end
            begin
              @(final_operation[32][31]) ;
              //$display("@%0t LEE: Received final operation event for 32,31\n", $time);
            end

            begin
              @(final_operation[33][0]) ;
              //$display("@%0t LEE: Received final operation event for 33,0\n", $time);
            end
            begin
              @(final_operation[33][1]) ;
              //$display("@%0t LEE: Received final operation event for 33,1\n", $time);
            end
            begin
              @(final_operation[33][2]) ;
              //$display("@%0t LEE: Received final operation event for 33,2\n", $time);
            end
            begin
              @(final_operation[33][3]) ;
              //$display("@%0t LEE: Received final operation event for 33,3\n", $time);
            end
            begin
              @(final_operation[33][4]) ;
              //$display("@%0t LEE: Received final operation event for 33,4\n", $time);
            end
            begin
              @(final_operation[33][5]) ;
              //$display("@%0t LEE: Received final operation event for 33,5\n", $time);
            end
            begin
              @(final_operation[33][6]) ;
              //$display("@%0t LEE: Received final operation event for 33,6\n", $time);
            end
            begin
              @(final_operation[33][7]) ;
              //$display("@%0t LEE: Received final operation event for 33,7\n", $time);
            end
            begin
              @(final_operation[33][8]) ;
              //$display("@%0t LEE: Received final operation event for 33,8\n", $time);
            end
            begin
              @(final_operation[33][9]) ;
              //$display("@%0t LEE: Received final operation event for 33,9\n", $time);
            end
            begin
              @(final_operation[33][10]) ;
              //$display("@%0t LEE: Received final operation event for 33,10\n", $time);
            end
            begin
              @(final_operation[33][11]) ;
              //$display("@%0t LEE: Received final operation event for 33,11\n", $time);
            end
            begin
              @(final_operation[33][12]) ;
              //$display("@%0t LEE: Received final operation event for 33,12\n", $time);
            end
            begin
              @(final_operation[33][13]) ;
              //$display("@%0t LEE: Received final operation event for 33,13\n", $time);
            end
            begin
              @(final_operation[33][14]) ;
              //$display("@%0t LEE: Received final operation event for 33,14\n", $time);
            end
            begin
              @(final_operation[33][15]) ;
              //$display("@%0t LEE: Received final operation event for 33,15\n", $time);
            end
            begin
              @(final_operation[33][16]) ;
              //$display("@%0t LEE: Received final operation event for 33,16\n", $time);
            end
            begin
              @(final_operation[33][17]) ;
              //$display("@%0t LEE: Received final operation event for 33,17\n", $time);
            end
            begin
              @(final_operation[33][18]) ;
              //$display("@%0t LEE: Received final operation event for 33,18\n", $time);
            end
            begin
              @(final_operation[33][19]) ;
              //$display("@%0t LEE: Received final operation event for 33,19\n", $time);
            end
            begin
              @(final_operation[33][20]) ;
              //$display("@%0t LEE: Received final operation event for 33,20\n", $time);
            end
            begin
              @(final_operation[33][21]) ;
              //$display("@%0t LEE: Received final operation event for 33,21\n", $time);
            end
            begin
              @(final_operation[33][22]) ;
              //$display("@%0t LEE: Received final operation event for 33,22\n", $time);
            end
            begin
              @(final_operation[33][23]) ;
              //$display("@%0t LEE: Received final operation event for 33,23\n", $time);
            end
            begin
              @(final_operation[33][24]) ;
              //$display("@%0t LEE: Received final operation event for 33,24\n", $time);
            end
            begin
              @(final_operation[33][25]) ;
              //$display("@%0t LEE: Received final operation event for 33,25\n", $time);
            end
            begin
              @(final_operation[33][26]) ;
              //$display("@%0t LEE: Received final operation event for 33,26\n", $time);
            end
            begin
              @(final_operation[33][27]) ;
              //$display("@%0t LEE: Received final operation event for 33,27\n", $time);
            end
            begin
              @(final_operation[33][28]) ;
              //$display("@%0t LEE: Received final operation event for 33,28\n", $time);
            end
            begin
              @(final_operation[33][29]) ;
              //$display("@%0t LEE: Received final operation event for 33,29\n", $time);
            end
            begin
              @(final_operation[33][30]) ;
              //$display("@%0t LEE: Received final operation event for 33,30\n", $time);
            end
            begin
              @(final_operation[33][31]) ;
              //$display("@%0t LEE: Received final operation event for 33,31\n", $time);
            end

            begin
              @(final_operation[34][0]) ;
              //$display("@%0t LEE: Received final operation event for 34,0\n", $time);
            end
            begin
              @(final_operation[34][1]) ;
              //$display("@%0t LEE: Received final operation event for 34,1\n", $time);
            end
            begin
              @(final_operation[34][2]) ;
              //$display("@%0t LEE: Received final operation event for 34,2\n", $time);
            end
            begin
              @(final_operation[34][3]) ;
              //$display("@%0t LEE: Received final operation event for 34,3\n", $time);
            end
            begin
              @(final_operation[34][4]) ;
              //$display("@%0t LEE: Received final operation event for 34,4\n", $time);
            end
            begin
              @(final_operation[34][5]) ;
              //$display("@%0t LEE: Received final operation event for 34,5\n", $time);
            end
            begin
              @(final_operation[34][6]) ;
              //$display("@%0t LEE: Received final operation event for 34,6\n", $time);
            end
            begin
              @(final_operation[34][7]) ;
              //$display("@%0t LEE: Received final operation event for 34,7\n", $time);
            end
            begin
              @(final_operation[34][8]) ;
              //$display("@%0t LEE: Received final operation event for 34,8\n", $time);
            end
            begin
              @(final_operation[34][9]) ;
              //$display("@%0t LEE: Received final operation event for 34,9\n", $time);
            end
            begin
              @(final_operation[34][10]) ;
              //$display("@%0t LEE: Received final operation event for 34,10\n", $time);
            end
            begin
              @(final_operation[34][11]) ;
              //$display("@%0t LEE: Received final operation event for 34,11\n", $time);
            end
            begin
              @(final_operation[34][12]) ;
              //$display("@%0t LEE: Received final operation event for 34,12\n", $time);
            end
            begin
              @(final_operation[34][13]) ;
              //$display("@%0t LEE: Received final operation event for 34,13\n", $time);
            end
            begin
              @(final_operation[34][14]) ;
              //$display("@%0t LEE: Received final operation event for 34,14\n", $time);
            end
            begin
              @(final_operation[34][15]) ;
              //$display("@%0t LEE: Received final operation event for 34,15\n", $time);
            end
            begin
              @(final_operation[34][16]) ;
              //$display("@%0t LEE: Received final operation event for 34,16\n", $time);
            end
            begin
              @(final_operation[34][17]) ;
              //$display("@%0t LEE: Received final operation event for 34,17\n", $time);
            end
            begin
              @(final_operation[34][18]) ;
              //$display("@%0t LEE: Received final operation event for 34,18\n", $time);
            end
            begin
              @(final_operation[34][19]) ;
              //$display("@%0t LEE: Received final operation event for 34,19\n", $time);
            end
            begin
              @(final_operation[34][20]) ;
              //$display("@%0t LEE: Received final operation event for 34,20\n", $time);
            end
            begin
              @(final_operation[34][21]) ;
              //$display("@%0t LEE: Received final operation event for 34,21\n", $time);
            end
            begin
              @(final_operation[34][22]) ;
              //$display("@%0t LEE: Received final operation event for 34,22\n", $time);
            end
            begin
              @(final_operation[34][23]) ;
              //$display("@%0t LEE: Received final operation event for 34,23\n", $time);
            end
            begin
              @(final_operation[34][24]) ;
              //$display("@%0t LEE: Received final operation event for 34,24\n", $time);
            end
            begin
              @(final_operation[34][25]) ;
              //$display("@%0t LEE: Received final operation event for 34,25\n", $time);
            end
            begin
              @(final_operation[34][26]) ;
              //$display("@%0t LEE: Received final operation event for 34,26\n", $time);
            end
            begin
              @(final_operation[34][27]) ;
              //$display("@%0t LEE: Received final operation event for 34,27\n", $time);
            end
            begin
              @(final_operation[34][28]) ;
              //$display("@%0t LEE: Received final operation event for 34,28\n", $time);
            end
            begin
              @(final_operation[34][29]) ;
              //$display("@%0t LEE: Received final operation event for 34,29\n", $time);
            end
            begin
              @(final_operation[34][30]) ;
              //$display("@%0t LEE: Received final operation event for 34,30\n", $time);
            end
            begin
              @(final_operation[34][31]) ;
              //$display("@%0t LEE: Received final operation event for 34,31\n", $time);
            end

            begin
              @(final_operation[35][0]) ;
              //$display("@%0t LEE: Received final operation event for 35,0\n", $time);
            end
            begin
              @(final_operation[35][1]) ;
              //$display("@%0t LEE: Received final operation event for 35,1\n", $time);
            end
            begin
              @(final_operation[35][2]) ;
              //$display("@%0t LEE: Received final operation event for 35,2\n", $time);
            end
            begin
              @(final_operation[35][3]) ;
              //$display("@%0t LEE: Received final operation event for 35,3\n", $time);
            end
            begin
              @(final_operation[35][4]) ;
              //$display("@%0t LEE: Received final operation event for 35,4\n", $time);
            end
            begin
              @(final_operation[35][5]) ;
              //$display("@%0t LEE: Received final operation event for 35,5\n", $time);
            end
            begin
              @(final_operation[35][6]) ;
              //$display("@%0t LEE: Received final operation event for 35,6\n", $time);
            end
            begin
              @(final_operation[35][7]) ;
              //$display("@%0t LEE: Received final operation event for 35,7\n", $time);
            end
            begin
              @(final_operation[35][8]) ;
              //$display("@%0t LEE: Received final operation event for 35,8\n", $time);
            end
            begin
              @(final_operation[35][9]) ;
              //$display("@%0t LEE: Received final operation event for 35,9\n", $time);
            end
            begin
              @(final_operation[35][10]) ;
              //$display("@%0t LEE: Received final operation event for 35,10\n", $time);
            end
            begin
              @(final_operation[35][11]) ;
              //$display("@%0t LEE: Received final operation event for 35,11\n", $time);
            end
            begin
              @(final_operation[35][12]) ;
              //$display("@%0t LEE: Received final operation event for 35,12\n", $time);
            end
            begin
              @(final_operation[35][13]) ;
              //$display("@%0t LEE: Received final operation event for 35,13\n", $time);
            end
            begin
              @(final_operation[35][14]) ;
              //$display("@%0t LEE: Received final operation event for 35,14\n", $time);
            end
            begin
              @(final_operation[35][15]) ;
              //$display("@%0t LEE: Received final operation event for 35,15\n", $time);
            end
            begin
              @(final_operation[35][16]) ;
              //$display("@%0t LEE: Received final operation event for 35,16\n", $time);
            end
            begin
              @(final_operation[35][17]) ;
              //$display("@%0t LEE: Received final operation event for 35,17\n", $time);
            end
            begin
              @(final_operation[35][18]) ;
              //$display("@%0t LEE: Received final operation event for 35,18\n", $time);
            end
            begin
              @(final_operation[35][19]) ;
              //$display("@%0t LEE: Received final operation event for 35,19\n", $time);
            end
            begin
              @(final_operation[35][20]) ;
              //$display("@%0t LEE: Received final operation event for 35,20\n", $time);
            end
            begin
              @(final_operation[35][21]) ;
              //$display("@%0t LEE: Received final operation event for 35,21\n", $time);
            end
            begin
              @(final_operation[35][22]) ;
              //$display("@%0t LEE: Received final operation event for 35,22\n", $time);
            end
            begin
              @(final_operation[35][23]) ;
              //$display("@%0t LEE: Received final operation event for 35,23\n", $time);
            end
            begin
              @(final_operation[35][24]) ;
              //$display("@%0t LEE: Received final operation event for 35,24\n", $time);
            end
            begin
              @(final_operation[35][25]) ;
              //$display("@%0t LEE: Received final operation event for 35,25\n", $time);
            end
            begin
              @(final_operation[35][26]) ;
              //$display("@%0t LEE: Received final operation event for 35,26\n", $time);
            end
            begin
              @(final_operation[35][27]) ;
              //$display("@%0t LEE: Received final operation event for 35,27\n", $time);
            end
            begin
              @(final_operation[35][28]) ;
              //$display("@%0t LEE: Received final operation event for 35,28\n", $time);
            end
            begin
              @(final_operation[35][29]) ;
              //$display("@%0t LEE: Received final operation event for 35,29\n", $time);
            end
            begin
              @(final_operation[35][30]) ;
              //$display("@%0t LEE: Received final operation event for 35,30\n", $time);
            end
            begin
              @(final_operation[35][31]) ;
              //$display("@%0t LEE: Received final operation event for 35,31\n", $time);
            end

            begin
              @(final_operation[36][0]) ;
              //$display("@%0t LEE: Received final operation event for 36,0\n", $time);
            end
            begin
              @(final_operation[36][1]) ;
              //$display("@%0t LEE: Received final operation event for 36,1\n", $time);
            end
            begin
              @(final_operation[36][2]) ;
              //$display("@%0t LEE: Received final operation event for 36,2\n", $time);
            end
            begin
              @(final_operation[36][3]) ;
              //$display("@%0t LEE: Received final operation event for 36,3\n", $time);
            end
            begin
              @(final_operation[36][4]) ;
              //$display("@%0t LEE: Received final operation event for 36,4\n", $time);
            end
            begin
              @(final_operation[36][5]) ;
              //$display("@%0t LEE: Received final operation event for 36,5\n", $time);
            end
            begin
              @(final_operation[36][6]) ;
              //$display("@%0t LEE: Received final operation event for 36,6\n", $time);
            end
            begin
              @(final_operation[36][7]) ;
              //$display("@%0t LEE: Received final operation event for 36,7\n", $time);
            end
            begin
              @(final_operation[36][8]) ;
              //$display("@%0t LEE: Received final operation event for 36,8\n", $time);
            end
            begin
              @(final_operation[36][9]) ;
              //$display("@%0t LEE: Received final operation event for 36,9\n", $time);
            end
            begin
              @(final_operation[36][10]) ;
              //$display("@%0t LEE: Received final operation event for 36,10\n", $time);
            end
            begin
              @(final_operation[36][11]) ;
              //$display("@%0t LEE: Received final operation event for 36,11\n", $time);
            end
            begin
              @(final_operation[36][12]) ;
              //$display("@%0t LEE: Received final operation event for 36,12\n", $time);
            end
            begin
              @(final_operation[36][13]) ;
              //$display("@%0t LEE: Received final operation event for 36,13\n", $time);
            end
            begin
              @(final_operation[36][14]) ;
              //$display("@%0t LEE: Received final operation event for 36,14\n", $time);
            end
            begin
              @(final_operation[36][15]) ;
              //$display("@%0t LEE: Received final operation event for 36,15\n", $time);
            end
            begin
              @(final_operation[36][16]) ;
              //$display("@%0t LEE: Received final operation event for 36,16\n", $time);
            end
            begin
              @(final_operation[36][17]) ;
              //$display("@%0t LEE: Received final operation event for 36,17\n", $time);
            end
            begin
              @(final_operation[36][18]) ;
              //$display("@%0t LEE: Received final operation event for 36,18\n", $time);
            end
            begin
              @(final_operation[36][19]) ;
              //$display("@%0t LEE: Received final operation event for 36,19\n", $time);
            end
            begin
              @(final_operation[36][20]) ;
              //$display("@%0t LEE: Received final operation event for 36,20\n", $time);
            end
            begin
              @(final_operation[36][21]) ;
              //$display("@%0t LEE: Received final operation event for 36,21\n", $time);
            end
            begin
              @(final_operation[36][22]) ;
              //$display("@%0t LEE: Received final operation event for 36,22\n", $time);
            end
            begin
              @(final_operation[36][23]) ;
              //$display("@%0t LEE: Received final operation event for 36,23\n", $time);
            end
            begin
              @(final_operation[36][24]) ;
              //$display("@%0t LEE: Received final operation event for 36,24\n", $time);
            end
            begin
              @(final_operation[36][25]) ;
              //$display("@%0t LEE: Received final operation event for 36,25\n", $time);
            end
            begin
              @(final_operation[36][26]) ;
              //$display("@%0t LEE: Received final operation event for 36,26\n", $time);
            end
            begin
              @(final_operation[36][27]) ;
              //$display("@%0t LEE: Received final operation event for 36,27\n", $time);
            end
            begin
              @(final_operation[36][28]) ;
              //$display("@%0t LEE: Received final operation event for 36,28\n", $time);
            end
            begin
              @(final_operation[36][29]) ;
              //$display("@%0t LEE: Received final operation event for 36,29\n", $time);
            end
            begin
              @(final_operation[36][30]) ;
              //$display("@%0t LEE: Received final operation event for 36,30\n", $time);
            end
            begin
              @(final_operation[36][31]) ;
              //$display("@%0t LEE: Received final operation event for 36,31\n", $time);
            end

            begin
              @(final_operation[37][0]) ;
              //$display("@%0t LEE: Received final operation event for 37,0\n", $time);
            end
            begin
              @(final_operation[37][1]) ;
              //$display("@%0t LEE: Received final operation event for 37,1\n", $time);
            end
            begin
              @(final_operation[37][2]) ;
              //$display("@%0t LEE: Received final operation event for 37,2\n", $time);
            end
            begin
              @(final_operation[37][3]) ;
              //$display("@%0t LEE: Received final operation event for 37,3\n", $time);
            end
            begin
              @(final_operation[37][4]) ;
              //$display("@%0t LEE: Received final operation event for 37,4\n", $time);
            end
            begin
              @(final_operation[37][5]) ;
              //$display("@%0t LEE: Received final operation event for 37,5\n", $time);
            end
            begin
              @(final_operation[37][6]) ;
              //$display("@%0t LEE: Received final operation event for 37,6\n", $time);
            end
            begin
              @(final_operation[37][7]) ;
              //$display("@%0t LEE: Received final operation event for 37,7\n", $time);
            end
            begin
              @(final_operation[37][8]) ;
              //$display("@%0t LEE: Received final operation event for 37,8\n", $time);
            end
            begin
              @(final_operation[37][9]) ;
              //$display("@%0t LEE: Received final operation event for 37,9\n", $time);
            end
            begin
              @(final_operation[37][10]) ;
              //$display("@%0t LEE: Received final operation event for 37,10\n", $time);
            end
            begin
              @(final_operation[37][11]) ;
              //$display("@%0t LEE: Received final operation event for 37,11\n", $time);
            end
            begin
              @(final_operation[37][12]) ;
              //$display("@%0t LEE: Received final operation event for 37,12\n", $time);
            end
            begin
              @(final_operation[37][13]) ;
              //$display("@%0t LEE: Received final operation event for 37,13\n", $time);
            end
            begin
              @(final_operation[37][14]) ;
              //$display("@%0t LEE: Received final operation event for 37,14\n", $time);
            end
            begin
              @(final_operation[37][15]) ;
              //$display("@%0t LEE: Received final operation event for 37,15\n", $time);
            end
            begin
              @(final_operation[37][16]) ;
              //$display("@%0t LEE: Received final operation event for 37,16\n", $time);
            end
            begin
              @(final_operation[37][17]) ;
              //$display("@%0t LEE: Received final operation event for 37,17\n", $time);
            end
            begin
              @(final_operation[37][18]) ;
              //$display("@%0t LEE: Received final operation event for 37,18\n", $time);
            end
            begin
              @(final_operation[37][19]) ;
              //$display("@%0t LEE: Received final operation event for 37,19\n", $time);
            end
            begin
              @(final_operation[37][20]) ;
              //$display("@%0t LEE: Received final operation event for 37,20\n", $time);
            end
            begin
              @(final_operation[37][21]) ;
              //$display("@%0t LEE: Received final operation event for 37,21\n", $time);
            end
            begin
              @(final_operation[37][22]) ;
              //$display("@%0t LEE: Received final operation event for 37,22\n", $time);
            end
            begin
              @(final_operation[37][23]) ;
              //$display("@%0t LEE: Received final operation event for 37,23\n", $time);
            end
            begin
              @(final_operation[37][24]) ;
              //$display("@%0t LEE: Received final operation event for 37,24\n", $time);
            end
            begin
              @(final_operation[37][25]) ;
              //$display("@%0t LEE: Received final operation event for 37,25\n", $time);
            end
            begin
              @(final_operation[37][26]) ;
              //$display("@%0t LEE: Received final operation event for 37,26\n", $time);
            end
            begin
              @(final_operation[37][27]) ;
              //$display("@%0t LEE: Received final operation event for 37,27\n", $time);
            end
            begin
              @(final_operation[37][28]) ;
              //$display("@%0t LEE: Received final operation event for 37,28\n", $time);
            end
            begin
              @(final_operation[37][29]) ;
              //$display("@%0t LEE: Received final operation event for 37,29\n", $time);
            end
            begin
              @(final_operation[37][30]) ;
              //$display("@%0t LEE: Received final operation event for 37,30\n", $time);
            end
            begin
              @(final_operation[37][31]) ;
              //$display("@%0t LEE: Received final operation event for 37,31\n", $time);
            end

            begin
              @(final_operation[38][0]) ;
              //$display("@%0t LEE: Received final operation event for 38,0\n", $time);
            end
            begin
              @(final_operation[38][1]) ;
              //$display("@%0t LEE: Received final operation event for 38,1\n", $time);
            end
            begin
              @(final_operation[38][2]) ;
              //$display("@%0t LEE: Received final operation event for 38,2\n", $time);
            end
            begin
              @(final_operation[38][3]) ;
              //$display("@%0t LEE: Received final operation event for 38,3\n", $time);
            end
            begin
              @(final_operation[38][4]) ;
              //$display("@%0t LEE: Received final operation event for 38,4\n", $time);
            end
            begin
              @(final_operation[38][5]) ;
              //$display("@%0t LEE: Received final operation event for 38,5\n", $time);
            end
            begin
              @(final_operation[38][6]) ;
              //$display("@%0t LEE: Received final operation event for 38,6\n", $time);
            end
            begin
              @(final_operation[38][7]) ;
              //$display("@%0t LEE: Received final operation event for 38,7\n", $time);
            end
            begin
              @(final_operation[38][8]) ;
              //$display("@%0t LEE: Received final operation event for 38,8\n", $time);
            end
            begin
              @(final_operation[38][9]) ;
              //$display("@%0t LEE: Received final operation event for 38,9\n", $time);
            end
            begin
              @(final_operation[38][10]) ;
              //$display("@%0t LEE: Received final operation event for 38,10\n", $time);
            end
            begin
              @(final_operation[38][11]) ;
              //$display("@%0t LEE: Received final operation event for 38,11\n", $time);
            end
            begin
              @(final_operation[38][12]) ;
              //$display("@%0t LEE: Received final operation event for 38,12\n", $time);
            end
            begin
              @(final_operation[38][13]) ;
              //$display("@%0t LEE: Received final operation event for 38,13\n", $time);
            end
            begin
              @(final_operation[38][14]) ;
              //$display("@%0t LEE: Received final operation event for 38,14\n", $time);
            end
            begin
              @(final_operation[38][15]) ;
              //$display("@%0t LEE: Received final operation event for 38,15\n", $time);
            end
            begin
              @(final_operation[38][16]) ;
              //$display("@%0t LEE: Received final operation event for 38,16\n", $time);
            end
            begin
              @(final_operation[38][17]) ;
              //$display("@%0t LEE: Received final operation event for 38,17\n", $time);
            end
            begin
              @(final_operation[38][18]) ;
              //$display("@%0t LEE: Received final operation event for 38,18\n", $time);
            end
            begin
              @(final_operation[38][19]) ;
              //$display("@%0t LEE: Received final operation event for 38,19\n", $time);
            end
            begin
              @(final_operation[38][20]) ;
              //$display("@%0t LEE: Received final operation event for 38,20\n", $time);
            end
            begin
              @(final_operation[38][21]) ;
              //$display("@%0t LEE: Received final operation event for 38,21\n", $time);
            end
            begin
              @(final_operation[38][22]) ;
              //$display("@%0t LEE: Received final operation event for 38,22\n", $time);
            end
            begin
              @(final_operation[38][23]) ;
              //$display("@%0t LEE: Received final operation event for 38,23\n", $time);
            end
            begin
              @(final_operation[38][24]) ;
              //$display("@%0t LEE: Received final operation event for 38,24\n", $time);
            end
            begin
              @(final_operation[38][25]) ;
              //$display("@%0t LEE: Received final operation event for 38,25\n", $time);
            end
            begin
              @(final_operation[38][26]) ;
              //$display("@%0t LEE: Received final operation event for 38,26\n", $time);
            end
            begin
              @(final_operation[38][27]) ;
              //$display("@%0t LEE: Received final operation event for 38,27\n", $time);
            end
            begin
              @(final_operation[38][28]) ;
              //$display("@%0t LEE: Received final operation event for 38,28\n", $time);
            end
            begin
              @(final_operation[38][29]) ;
              //$display("@%0t LEE: Received final operation event for 38,29\n", $time);
            end
            begin
              @(final_operation[38][30]) ;
              //$display("@%0t LEE: Received final operation event for 38,30\n", $time);
            end
            begin
              @(final_operation[38][31]) ;
              //$display("@%0t LEE: Received final operation event for 38,31\n", $time);
            end

            begin
              @(final_operation[39][0]) ;
              //$display("@%0t LEE: Received final operation event for 39,0\n", $time);
            end
            begin
              @(final_operation[39][1]) ;
              //$display("@%0t LEE: Received final operation event for 39,1\n", $time);
            end
            begin
              @(final_operation[39][2]) ;
              //$display("@%0t LEE: Received final operation event for 39,2\n", $time);
            end
            begin
              @(final_operation[39][3]) ;
              //$display("@%0t LEE: Received final operation event for 39,3\n", $time);
            end
            begin
              @(final_operation[39][4]) ;
              //$display("@%0t LEE: Received final operation event for 39,4\n", $time);
            end
            begin
              @(final_operation[39][5]) ;
              //$display("@%0t LEE: Received final operation event for 39,5\n", $time);
            end
            begin
              @(final_operation[39][6]) ;
              //$display("@%0t LEE: Received final operation event for 39,6\n", $time);
            end
            begin
              @(final_operation[39][7]) ;
              //$display("@%0t LEE: Received final operation event for 39,7\n", $time);
            end
            begin
              @(final_operation[39][8]) ;
              //$display("@%0t LEE: Received final operation event for 39,8\n", $time);
            end
            begin
              @(final_operation[39][9]) ;
              //$display("@%0t LEE: Received final operation event for 39,9\n", $time);
            end
            begin
              @(final_operation[39][10]) ;
              //$display("@%0t LEE: Received final operation event for 39,10\n", $time);
            end
            begin
              @(final_operation[39][11]) ;
              //$display("@%0t LEE: Received final operation event for 39,11\n", $time);
            end
            begin
              @(final_operation[39][12]) ;
              //$display("@%0t LEE: Received final operation event for 39,12\n", $time);
            end
            begin
              @(final_operation[39][13]) ;
              //$display("@%0t LEE: Received final operation event for 39,13\n", $time);
            end
            begin
              @(final_operation[39][14]) ;
              //$display("@%0t LEE: Received final operation event for 39,14\n", $time);
            end
            begin
              @(final_operation[39][15]) ;
              //$display("@%0t LEE: Received final operation event for 39,15\n", $time);
            end
            begin
              @(final_operation[39][16]) ;
              //$display("@%0t LEE: Received final operation event for 39,16\n", $time);
            end
            begin
              @(final_operation[39][17]) ;
              //$display("@%0t LEE: Received final operation event for 39,17\n", $time);
            end
            begin
              @(final_operation[39][18]) ;
              //$display("@%0t LEE: Received final operation event for 39,18\n", $time);
            end
            begin
              @(final_operation[39][19]) ;
              //$display("@%0t LEE: Received final operation event for 39,19\n", $time);
            end
            begin
              @(final_operation[39][20]) ;
              //$display("@%0t LEE: Received final operation event for 39,20\n", $time);
            end
            begin
              @(final_operation[39][21]) ;
              //$display("@%0t LEE: Received final operation event for 39,21\n", $time);
            end
            begin
              @(final_operation[39][22]) ;
              //$display("@%0t LEE: Received final operation event for 39,22\n", $time);
            end
            begin
              @(final_operation[39][23]) ;
              //$display("@%0t LEE: Received final operation event for 39,23\n", $time);
            end
            begin
              @(final_operation[39][24]) ;
              //$display("@%0t LEE: Received final operation event for 39,24\n", $time);
            end
            begin
              @(final_operation[39][25]) ;
              //$display("@%0t LEE: Received final operation event for 39,25\n", $time);
            end
            begin
              @(final_operation[39][26]) ;
              //$display("@%0t LEE: Received final operation event for 39,26\n", $time);
            end
            begin
              @(final_operation[39][27]) ;
              //$display("@%0t LEE: Received final operation event for 39,27\n", $time);
            end
            begin
              @(final_operation[39][28]) ;
              //$display("@%0t LEE: Received final operation event for 39,28\n", $time);
            end
            begin
              @(final_operation[39][29]) ;
              //$display("@%0t LEE: Received final operation event for 39,29\n", $time);
            end
            begin
              @(final_operation[39][30]) ;
              //$display("@%0t LEE: Received final operation event for 39,30\n", $time);
            end
            begin
              @(final_operation[39][31]) ;
              //$display("@%0t LEE: Received final operation event for 39,31\n", $time);
            end

            begin
              @(final_operation[40][0]) ;
              //$display("@%0t LEE: Received final operation event for 40,0\n", $time);
            end
            begin
              @(final_operation[40][1]) ;
              //$display("@%0t LEE: Received final operation event for 40,1\n", $time);
            end
            begin
              @(final_operation[40][2]) ;
              //$display("@%0t LEE: Received final operation event for 40,2\n", $time);
            end
            begin
              @(final_operation[40][3]) ;
              //$display("@%0t LEE: Received final operation event for 40,3\n", $time);
            end
            begin
              @(final_operation[40][4]) ;
              //$display("@%0t LEE: Received final operation event for 40,4\n", $time);
            end
            begin
              @(final_operation[40][5]) ;
              //$display("@%0t LEE: Received final operation event for 40,5\n", $time);
            end
            begin
              @(final_operation[40][6]) ;
              //$display("@%0t LEE: Received final operation event for 40,6\n", $time);
            end
            begin
              @(final_operation[40][7]) ;
              //$display("@%0t LEE: Received final operation event for 40,7\n", $time);
            end
            begin
              @(final_operation[40][8]) ;
              //$display("@%0t LEE: Received final operation event for 40,8\n", $time);
            end
            begin
              @(final_operation[40][9]) ;
              //$display("@%0t LEE: Received final operation event for 40,9\n", $time);
            end
            begin
              @(final_operation[40][10]) ;
              //$display("@%0t LEE: Received final operation event for 40,10\n", $time);
            end
            begin
              @(final_operation[40][11]) ;
              //$display("@%0t LEE: Received final operation event for 40,11\n", $time);
            end
            begin
              @(final_operation[40][12]) ;
              //$display("@%0t LEE: Received final operation event for 40,12\n", $time);
            end
            begin
              @(final_operation[40][13]) ;
              //$display("@%0t LEE: Received final operation event for 40,13\n", $time);
            end
            begin
              @(final_operation[40][14]) ;
              //$display("@%0t LEE: Received final operation event for 40,14\n", $time);
            end
            begin
              @(final_operation[40][15]) ;
              //$display("@%0t LEE: Received final operation event for 40,15\n", $time);
            end
            begin
              @(final_operation[40][16]) ;
              //$display("@%0t LEE: Received final operation event for 40,16\n", $time);
            end
            begin
              @(final_operation[40][17]) ;
              //$display("@%0t LEE: Received final operation event for 40,17\n", $time);
            end
            begin
              @(final_operation[40][18]) ;
              //$display("@%0t LEE: Received final operation event for 40,18\n", $time);
            end
            begin
              @(final_operation[40][19]) ;
              //$display("@%0t LEE: Received final operation event for 40,19\n", $time);
            end
            begin
              @(final_operation[40][20]) ;
              //$display("@%0t LEE: Received final operation event for 40,20\n", $time);
            end
            begin
              @(final_operation[40][21]) ;
              //$display("@%0t LEE: Received final operation event for 40,21\n", $time);
            end
            begin
              @(final_operation[40][22]) ;
              //$display("@%0t LEE: Received final operation event for 40,22\n", $time);
            end
            begin
              @(final_operation[40][23]) ;
              //$display("@%0t LEE: Received final operation event for 40,23\n", $time);
            end
            begin
              @(final_operation[40][24]) ;
              //$display("@%0t LEE: Received final operation event for 40,24\n", $time);
            end
            begin
              @(final_operation[40][25]) ;
              //$display("@%0t LEE: Received final operation event for 40,25\n", $time);
            end
            begin
              @(final_operation[40][26]) ;
              //$display("@%0t LEE: Received final operation event for 40,26\n", $time);
            end
            begin
              @(final_operation[40][27]) ;
              //$display("@%0t LEE: Received final operation event for 40,27\n", $time);
            end
            begin
              @(final_operation[40][28]) ;
              //$display("@%0t LEE: Received final operation event for 40,28\n", $time);
            end
            begin
              @(final_operation[40][29]) ;
              //$display("@%0t LEE: Received final operation event for 40,29\n", $time);
            end
            begin
              @(final_operation[40][30]) ;
              //$display("@%0t LEE: Received final operation event for 40,30\n", $time);
            end
            begin
              @(final_operation[40][31]) ;
              //$display("@%0t LEE: Received final operation event for 40,31\n", $time);
            end

            begin
              @(final_operation[41][0]) ;
              //$display("@%0t LEE: Received final operation event for 41,0\n", $time);
            end
            begin
              @(final_operation[41][1]) ;
              //$display("@%0t LEE: Received final operation event for 41,1\n", $time);
            end
            begin
              @(final_operation[41][2]) ;
              //$display("@%0t LEE: Received final operation event for 41,2\n", $time);
            end
            begin
              @(final_operation[41][3]) ;
              //$display("@%0t LEE: Received final operation event for 41,3\n", $time);
            end
            begin
              @(final_operation[41][4]) ;
              //$display("@%0t LEE: Received final operation event for 41,4\n", $time);
            end
            begin
              @(final_operation[41][5]) ;
              //$display("@%0t LEE: Received final operation event for 41,5\n", $time);
            end
            begin
              @(final_operation[41][6]) ;
              //$display("@%0t LEE: Received final operation event for 41,6\n", $time);
            end
            begin
              @(final_operation[41][7]) ;
              //$display("@%0t LEE: Received final operation event for 41,7\n", $time);
            end
            begin
              @(final_operation[41][8]) ;
              //$display("@%0t LEE: Received final operation event for 41,8\n", $time);
            end
            begin
              @(final_operation[41][9]) ;
              //$display("@%0t LEE: Received final operation event for 41,9\n", $time);
            end
            begin
              @(final_operation[41][10]) ;
              //$display("@%0t LEE: Received final operation event for 41,10\n", $time);
            end
            begin
              @(final_operation[41][11]) ;
              //$display("@%0t LEE: Received final operation event for 41,11\n", $time);
            end
            begin
              @(final_operation[41][12]) ;
              //$display("@%0t LEE: Received final operation event for 41,12\n", $time);
            end
            begin
              @(final_operation[41][13]) ;
              //$display("@%0t LEE: Received final operation event for 41,13\n", $time);
            end
            begin
              @(final_operation[41][14]) ;
              //$display("@%0t LEE: Received final operation event for 41,14\n", $time);
            end
            begin
              @(final_operation[41][15]) ;
              //$display("@%0t LEE: Received final operation event for 41,15\n", $time);
            end
            begin
              @(final_operation[41][16]) ;
              //$display("@%0t LEE: Received final operation event for 41,16\n", $time);
            end
            begin
              @(final_operation[41][17]) ;
              //$display("@%0t LEE: Received final operation event for 41,17\n", $time);
            end
            begin
              @(final_operation[41][18]) ;
              //$display("@%0t LEE: Received final operation event for 41,18\n", $time);
            end
            begin
              @(final_operation[41][19]) ;
              //$display("@%0t LEE: Received final operation event for 41,19\n", $time);
            end
            begin
              @(final_operation[41][20]) ;
              //$display("@%0t LEE: Received final operation event for 41,20\n", $time);
            end
            begin
              @(final_operation[41][21]) ;
              //$display("@%0t LEE: Received final operation event for 41,21\n", $time);
            end
            begin
              @(final_operation[41][22]) ;
              //$display("@%0t LEE: Received final operation event for 41,22\n", $time);
            end
            begin
              @(final_operation[41][23]) ;
              //$display("@%0t LEE: Received final operation event for 41,23\n", $time);
            end
            begin
              @(final_operation[41][24]) ;
              //$display("@%0t LEE: Received final operation event for 41,24\n", $time);
            end
            begin
              @(final_operation[41][25]) ;
              //$display("@%0t LEE: Received final operation event for 41,25\n", $time);
            end
            begin
              @(final_operation[41][26]) ;
              //$display("@%0t LEE: Received final operation event for 41,26\n", $time);
            end
            begin
              @(final_operation[41][27]) ;
              //$display("@%0t LEE: Received final operation event for 41,27\n", $time);
            end
            begin
              @(final_operation[41][28]) ;
              //$display("@%0t LEE: Received final operation event for 41,28\n", $time);
            end
            begin
              @(final_operation[41][29]) ;
              //$display("@%0t LEE: Received final operation event for 41,29\n", $time);
            end
            begin
              @(final_operation[41][30]) ;
              //$display("@%0t LEE: Received final operation event for 41,30\n", $time);
            end
            begin
              @(final_operation[41][31]) ;
              //$display("@%0t LEE: Received final operation event for 41,31\n", $time);
            end

            begin
              @(final_operation[42][0]) ;
              //$display("@%0t LEE: Received final operation event for 42,0\n", $time);
            end
            begin
              @(final_operation[42][1]) ;
              //$display("@%0t LEE: Received final operation event for 42,1\n", $time);
            end
            begin
              @(final_operation[42][2]) ;
              //$display("@%0t LEE: Received final operation event for 42,2\n", $time);
            end
            begin
              @(final_operation[42][3]) ;
              //$display("@%0t LEE: Received final operation event for 42,3\n", $time);
            end
            begin
              @(final_operation[42][4]) ;
              //$display("@%0t LEE: Received final operation event for 42,4\n", $time);
            end
            begin
              @(final_operation[42][5]) ;
              //$display("@%0t LEE: Received final operation event for 42,5\n", $time);
            end
            begin
              @(final_operation[42][6]) ;
              //$display("@%0t LEE: Received final operation event for 42,6\n", $time);
            end
            begin
              @(final_operation[42][7]) ;
              //$display("@%0t LEE: Received final operation event for 42,7\n", $time);
            end
            begin
              @(final_operation[42][8]) ;
              //$display("@%0t LEE: Received final operation event for 42,8\n", $time);
            end
            begin
              @(final_operation[42][9]) ;
              //$display("@%0t LEE: Received final operation event for 42,9\n", $time);
            end
            begin
              @(final_operation[42][10]) ;
              //$display("@%0t LEE: Received final operation event for 42,10\n", $time);
            end
            begin
              @(final_operation[42][11]) ;
              //$display("@%0t LEE: Received final operation event for 42,11\n", $time);
            end
            begin
              @(final_operation[42][12]) ;
              //$display("@%0t LEE: Received final operation event for 42,12\n", $time);
            end
            begin
              @(final_operation[42][13]) ;
              //$display("@%0t LEE: Received final operation event for 42,13\n", $time);
            end
            begin
              @(final_operation[42][14]) ;
              //$display("@%0t LEE: Received final operation event for 42,14\n", $time);
            end
            begin
              @(final_operation[42][15]) ;
              //$display("@%0t LEE: Received final operation event for 42,15\n", $time);
            end
            begin
              @(final_operation[42][16]) ;
              //$display("@%0t LEE: Received final operation event for 42,16\n", $time);
            end
            begin
              @(final_operation[42][17]) ;
              //$display("@%0t LEE: Received final operation event for 42,17\n", $time);
            end
            begin
              @(final_operation[42][18]) ;
              //$display("@%0t LEE: Received final operation event for 42,18\n", $time);
            end
            begin
              @(final_operation[42][19]) ;
              //$display("@%0t LEE: Received final operation event for 42,19\n", $time);
            end
            begin
              @(final_operation[42][20]) ;
              //$display("@%0t LEE: Received final operation event for 42,20\n", $time);
            end
            begin
              @(final_operation[42][21]) ;
              //$display("@%0t LEE: Received final operation event for 42,21\n", $time);
            end
            begin
              @(final_operation[42][22]) ;
              //$display("@%0t LEE: Received final operation event for 42,22\n", $time);
            end
            begin
              @(final_operation[42][23]) ;
              //$display("@%0t LEE: Received final operation event for 42,23\n", $time);
            end
            begin
              @(final_operation[42][24]) ;
              //$display("@%0t LEE: Received final operation event for 42,24\n", $time);
            end
            begin
              @(final_operation[42][25]) ;
              //$display("@%0t LEE: Received final operation event for 42,25\n", $time);
            end
            begin
              @(final_operation[42][26]) ;
              //$display("@%0t LEE: Received final operation event for 42,26\n", $time);
            end
            begin
              @(final_operation[42][27]) ;
              //$display("@%0t LEE: Received final operation event for 42,27\n", $time);
            end
            begin
              @(final_operation[42][28]) ;
              //$display("@%0t LEE: Received final operation event for 42,28\n", $time);
            end
            begin
              @(final_operation[42][29]) ;
              //$display("@%0t LEE: Received final operation event for 42,29\n", $time);
            end
            begin
              @(final_operation[42][30]) ;
              //$display("@%0t LEE: Received final operation event for 42,30\n", $time);
            end
            begin
              @(final_operation[42][31]) ;
              //$display("@%0t LEE: Received final operation event for 42,31\n", $time);
            end

            begin
              @(final_operation[43][0]) ;
              //$display("@%0t LEE: Received final operation event for 43,0\n", $time);
            end
            begin
              @(final_operation[43][1]) ;
              //$display("@%0t LEE: Received final operation event for 43,1\n", $time);
            end
            begin
              @(final_operation[43][2]) ;
              //$display("@%0t LEE: Received final operation event for 43,2\n", $time);
            end
            begin
              @(final_operation[43][3]) ;
              //$display("@%0t LEE: Received final operation event for 43,3\n", $time);
            end
            begin
              @(final_operation[43][4]) ;
              //$display("@%0t LEE: Received final operation event for 43,4\n", $time);
            end
            begin
              @(final_operation[43][5]) ;
              //$display("@%0t LEE: Received final operation event for 43,5\n", $time);
            end
            begin
              @(final_operation[43][6]) ;
              //$display("@%0t LEE: Received final operation event for 43,6\n", $time);
            end
            begin
              @(final_operation[43][7]) ;
              //$display("@%0t LEE: Received final operation event for 43,7\n", $time);
            end
            begin
              @(final_operation[43][8]) ;
              //$display("@%0t LEE: Received final operation event for 43,8\n", $time);
            end
            begin
              @(final_operation[43][9]) ;
              //$display("@%0t LEE: Received final operation event for 43,9\n", $time);
            end
            begin
              @(final_operation[43][10]) ;
              //$display("@%0t LEE: Received final operation event for 43,10\n", $time);
            end
            begin
              @(final_operation[43][11]) ;
              //$display("@%0t LEE: Received final operation event for 43,11\n", $time);
            end
            begin
              @(final_operation[43][12]) ;
              //$display("@%0t LEE: Received final operation event for 43,12\n", $time);
            end
            begin
              @(final_operation[43][13]) ;
              //$display("@%0t LEE: Received final operation event for 43,13\n", $time);
            end
            begin
              @(final_operation[43][14]) ;
              //$display("@%0t LEE: Received final operation event for 43,14\n", $time);
            end
            begin
              @(final_operation[43][15]) ;
              //$display("@%0t LEE: Received final operation event for 43,15\n", $time);
            end
            begin
              @(final_operation[43][16]) ;
              //$display("@%0t LEE: Received final operation event for 43,16\n", $time);
            end
            begin
              @(final_operation[43][17]) ;
              //$display("@%0t LEE: Received final operation event for 43,17\n", $time);
            end
            begin
              @(final_operation[43][18]) ;
              //$display("@%0t LEE: Received final operation event for 43,18\n", $time);
            end
            begin
              @(final_operation[43][19]) ;
              //$display("@%0t LEE: Received final operation event for 43,19\n", $time);
            end
            begin
              @(final_operation[43][20]) ;
              //$display("@%0t LEE: Received final operation event for 43,20\n", $time);
            end
            begin
              @(final_operation[43][21]) ;
              //$display("@%0t LEE: Received final operation event for 43,21\n", $time);
            end
            begin
              @(final_operation[43][22]) ;
              //$display("@%0t LEE: Received final operation event for 43,22\n", $time);
            end
            begin
              @(final_operation[43][23]) ;
              //$display("@%0t LEE: Received final operation event for 43,23\n", $time);
            end
            begin
              @(final_operation[43][24]) ;
              //$display("@%0t LEE: Received final operation event for 43,24\n", $time);
            end
            begin
              @(final_operation[43][25]) ;
              //$display("@%0t LEE: Received final operation event for 43,25\n", $time);
            end
            begin
              @(final_operation[43][26]) ;
              //$display("@%0t LEE: Received final operation event for 43,26\n", $time);
            end
            begin
              @(final_operation[43][27]) ;
              //$display("@%0t LEE: Received final operation event for 43,27\n", $time);
            end
            begin
              @(final_operation[43][28]) ;
              //$display("@%0t LEE: Received final operation event for 43,28\n", $time);
            end
            begin
              @(final_operation[43][29]) ;
              //$display("@%0t LEE: Received final operation event for 43,29\n", $time);
            end
            begin
              @(final_operation[43][30]) ;
              //$display("@%0t LEE: Received final operation event for 43,30\n", $time);
            end
            begin
              @(final_operation[43][31]) ;
              //$display("@%0t LEE: Received final operation event for 43,31\n", $time);
            end

            begin
              @(final_operation[44][0]) ;
              //$display("@%0t LEE: Received final operation event for 44,0\n", $time);
            end
            begin
              @(final_operation[44][1]) ;
              //$display("@%0t LEE: Received final operation event for 44,1\n", $time);
            end
            begin
              @(final_operation[44][2]) ;
              //$display("@%0t LEE: Received final operation event for 44,2\n", $time);
            end
            begin
              @(final_operation[44][3]) ;
              //$display("@%0t LEE: Received final operation event for 44,3\n", $time);
            end
            begin
              @(final_operation[44][4]) ;
              //$display("@%0t LEE: Received final operation event for 44,4\n", $time);
            end
            begin
              @(final_operation[44][5]) ;
              //$display("@%0t LEE: Received final operation event for 44,5\n", $time);
            end
            begin
              @(final_operation[44][6]) ;
              //$display("@%0t LEE: Received final operation event for 44,6\n", $time);
            end
            begin
              @(final_operation[44][7]) ;
              //$display("@%0t LEE: Received final operation event for 44,7\n", $time);
            end
            begin
              @(final_operation[44][8]) ;
              //$display("@%0t LEE: Received final operation event for 44,8\n", $time);
            end
            begin
              @(final_operation[44][9]) ;
              //$display("@%0t LEE: Received final operation event for 44,9\n", $time);
            end
            begin
              @(final_operation[44][10]) ;
              //$display("@%0t LEE: Received final operation event for 44,10\n", $time);
            end
            begin
              @(final_operation[44][11]) ;
              //$display("@%0t LEE: Received final operation event for 44,11\n", $time);
            end
            begin
              @(final_operation[44][12]) ;
              //$display("@%0t LEE: Received final operation event for 44,12\n", $time);
            end
            begin
              @(final_operation[44][13]) ;
              //$display("@%0t LEE: Received final operation event for 44,13\n", $time);
            end
            begin
              @(final_operation[44][14]) ;
              //$display("@%0t LEE: Received final operation event for 44,14\n", $time);
            end
            begin
              @(final_operation[44][15]) ;
              //$display("@%0t LEE: Received final operation event for 44,15\n", $time);
            end
            begin
              @(final_operation[44][16]) ;
              //$display("@%0t LEE: Received final operation event for 44,16\n", $time);
            end
            begin
              @(final_operation[44][17]) ;
              //$display("@%0t LEE: Received final operation event for 44,17\n", $time);
            end
            begin
              @(final_operation[44][18]) ;
              //$display("@%0t LEE: Received final operation event for 44,18\n", $time);
            end
            begin
              @(final_operation[44][19]) ;
              //$display("@%0t LEE: Received final operation event for 44,19\n", $time);
            end
            begin
              @(final_operation[44][20]) ;
              //$display("@%0t LEE: Received final operation event for 44,20\n", $time);
            end
            begin
              @(final_operation[44][21]) ;
              //$display("@%0t LEE: Received final operation event for 44,21\n", $time);
            end
            begin
              @(final_operation[44][22]) ;
              //$display("@%0t LEE: Received final operation event for 44,22\n", $time);
            end
            begin
              @(final_operation[44][23]) ;
              //$display("@%0t LEE: Received final operation event for 44,23\n", $time);
            end
            begin
              @(final_operation[44][24]) ;
              //$display("@%0t LEE: Received final operation event for 44,24\n", $time);
            end
            begin
              @(final_operation[44][25]) ;
              //$display("@%0t LEE: Received final operation event for 44,25\n", $time);
            end
            begin
              @(final_operation[44][26]) ;
              //$display("@%0t LEE: Received final operation event for 44,26\n", $time);
            end
            begin
              @(final_operation[44][27]) ;
              //$display("@%0t LEE: Received final operation event for 44,27\n", $time);
            end
            begin
              @(final_operation[44][28]) ;
              //$display("@%0t LEE: Received final operation event for 44,28\n", $time);
            end
            begin
              @(final_operation[44][29]) ;
              //$display("@%0t LEE: Received final operation event for 44,29\n", $time);
            end
            begin
              @(final_operation[44][30]) ;
              //$display("@%0t LEE: Received final operation event for 44,30\n", $time);
            end
            begin
              @(final_operation[44][31]) ;
              //$display("@%0t LEE: Received final operation event for 44,31\n", $time);
            end

            begin
              @(final_operation[45][0]) ;
              //$display("@%0t LEE: Received final operation event for 45,0\n", $time);
            end
            begin
              @(final_operation[45][1]) ;
              //$display("@%0t LEE: Received final operation event for 45,1\n", $time);
            end
            begin
              @(final_operation[45][2]) ;
              //$display("@%0t LEE: Received final operation event for 45,2\n", $time);
            end
            begin
              @(final_operation[45][3]) ;
              //$display("@%0t LEE: Received final operation event for 45,3\n", $time);
            end
            begin
              @(final_operation[45][4]) ;
              //$display("@%0t LEE: Received final operation event for 45,4\n", $time);
            end
            begin
              @(final_operation[45][5]) ;
              //$display("@%0t LEE: Received final operation event for 45,5\n", $time);
            end
            begin
              @(final_operation[45][6]) ;
              //$display("@%0t LEE: Received final operation event for 45,6\n", $time);
            end
            begin
              @(final_operation[45][7]) ;
              //$display("@%0t LEE: Received final operation event for 45,7\n", $time);
            end
            begin
              @(final_operation[45][8]) ;
              //$display("@%0t LEE: Received final operation event for 45,8\n", $time);
            end
            begin
              @(final_operation[45][9]) ;
              //$display("@%0t LEE: Received final operation event for 45,9\n", $time);
            end
            begin
              @(final_operation[45][10]) ;
              //$display("@%0t LEE: Received final operation event for 45,10\n", $time);
            end
            begin
              @(final_operation[45][11]) ;
              //$display("@%0t LEE: Received final operation event for 45,11\n", $time);
            end
            begin
              @(final_operation[45][12]) ;
              //$display("@%0t LEE: Received final operation event for 45,12\n", $time);
            end
            begin
              @(final_operation[45][13]) ;
              //$display("@%0t LEE: Received final operation event for 45,13\n", $time);
            end
            begin
              @(final_operation[45][14]) ;
              //$display("@%0t LEE: Received final operation event for 45,14\n", $time);
            end
            begin
              @(final_operation[45][15]) ;
              //$display("@%0t LEE: Received final operation event for 45,15\n", $time);
            end
            begin
              @(final_operation[45][16]) ;
              //$display("@%0t LEE: Received final operation event for 45,16\n", $time);
            end
            begin
              @(final_operation[45][17]) ;
              //$display("@%0t LEE: Received final operation event for 45,17\n", $time);
            end
            begin
              @(final_operation[45][18]) ;
              //$display("@%0t LEE: Received final operation event for 45,18\n", $time);
            end
            begin
              @(final_operation[45][19]) ;
              //$display("@%0t LEE: Received final operation event for 45,19\n", $time);
            end
            begin
              @(final_operation[45][20]) ;
              //$display("@%0t LEE: Received final operation event for 45,20\n", $time);
            end
            begin
              @(final_operation[45][21]) ;
              //$display("@%0t LEE: Received final operation event for 45,21\n", $time);
            end
            begin
              @(final_operation[45][22]) ;
              //$display("@%0t LEE: Received final operation event for 45,22\n", $time);
            end
            begin
              @(final_operation[45][23]) ;
              //$display("@%0t LEE: Received final operation event for 45,23\n", $time);
            end
            begin
              @(final_operation[45][24]) ;
              //$display("@%0t LEE: Received final operation event for 45,24\n", $time);
            end
            begin
              @(final_operation[45][25]) ;
              //$display("@%0t LEE: Received final operation event for 45,25\n", $time);
            end
            begin
              @(final_operation[45][26]) ;
              //$display("@%0t LEE: Received final operation event for 45,26\n", $time);
            end
            begin
              @(final_operation[45][27]) ;
              //$display("@%0t LEE: Received final operation event for 45,27\n", $time);
            end
            begin
              @(final_operation[45][28]) ;
              //$display("@%0t LEE: Received final operation event for 45,28\n", $time);
            end
            begin
              @(final_operation[45][29]) ;
              //$display("@%0t LEE: Received final operation event for 45,29\n", $time);
            end
            begin
              @(final_operation[45][30]) ;
              //$display("@%0t LEE: Received final operation event for 45,30\n", $time);
            end
            begin
              @(final_operation[45][31]) ;
              //$display("@%0t LEE: Received final operation event for 45,31\n", $time);
            end

            begin
              @(final_operation[46][0]) ;
              //$display("@%0t LEE: Received final operation event for 46,0\n", $time);
            end
            begin
              @(final_operation[46][1]) ;
              //$display("@%0t LEE: Received final operation event for 46,1\n", $time);
            end
            begin
              @(final_operation[46][2]) ;
              //$display("@%0t LEE: Received final operation event for 46,2\n", $time);
            end
            begin
              @(final_operation[46][3]) ;
              //$display("@%0t LEE: Received final operation event for 46,3\n", $time);
            end
            begin
              @(final_operation[46][4]) ;
              //$display("@%0t LEE: Received final operation event for 46,4\n", $time);
            end
            begin
              @(final_operation[46][5]) ;
              //$display("@%0t LEE: Received final operation event for 46,5\n", $time);
            end
            begin
              @(final_operation[46][6]) ;
              //$display("@%0t LEE: Received final operation event for 46,6\n", $time);
            end
            begin
              @(final_operation[46][7]) ;
              //$display("@%0t LEE: Received final operation event for 46,7\n", $time);
            end
            begin
              @(final_operation[46][8]) ;
              //$display("@%0t LEE: Received final operation event for 46,8\n", $time);
            end
            begin
              @(final_operation[46][9]) ;
              //$display("@%0t LEE: Received final operation event for 46,9\n", $time);
            end
            begin
              @(final_operation[46][10]) ;
              //$display("@%0t LEE: Received final operation event for 46,10\n", $time);
            end
            begin
              @(final_operation[46][11]) ;
              //$display("@%0t LEE: Received final operation event for 46,11\n", $time);
            end
            begin
              @(final_operation[46][12]) ;
              //$display("@%0t LEE: Received final operation event for 46,12\n", $time);
            end
            begin
              @(final_operation[46][13]) ;
              //$display("@%0t LEE: Received final operation event for 46,13\n", $time);
            end
            begin
              @(final_operation[46][14]) ;
              //$display("@%0t LEE: Received final operation event for 46,14\n", $time);
            end
            begin
              @(final_operation[46][15]) ;
              //$display("@%0t LEE: Received final operation event for 46,15\n", $time);
            end
            begin
              @(final_operation[46][16]) ;
              //$display("@%0t LEE: Received final operation event for 46,16\n", $time);
            end
            begin
              @(final_operation[46][17]) ;
              //$display("@%0t LEE: Received final operation event for 46,17\n", $time);
            end
            begin
              @(final_operation[46][18]) ;
              //$display("@%0t LEE: Received final operation event for 46,18\n", $time);
            end
            begin
              @(final_operation[46][19]) ;
              //$display("@%0t LEE: Received final operation event for 46,19\n", $time);
            end
            begin
              @(final_operation[46][20]) ;
              //$display("@%0t LEE: Received final operation event for 46,20\n", $time);
            end
            begin
              @(final_operation[46][21]) ;
              //$display("@%0t LEE: Received final operation event for 46,21\n", $time);
            end
            begin
              @(final_operation[46][22]) ;
              //$display("@%0t LEE: Received final operation event for 46,22\n", $time);
            end
            begin
              @(final_operation[46][23]) ;
              //$display("@%0t LEE: Received final operation event for 46,23\n", $time);
            end
            begin
              @(final_operation[46][24]) ;
              //$display("@%0t LEE: Received final operation event for 46,24\n", $time);
            end
            begin
              @(final_operation[46][25]) ;
              //$display("@%0t LEE: Received final operation event for 46,25\n", $time);
            end
            begin
              @(final_operation[46][26]) ;
              //$display("@%0t LEE: Received final operation event for 46,26\n", $time);
            end
            begin
              @(final_operation[46][27]) ;
              //$display("@%0t LEE: Received final operation event for 46,27\n", $time);
            end
            begin
              @(final_operation[46][28]) ;
              //$display("@%0t LEE: Received final operation event for 46,28\n", $time);
            end
            begin
              @(final_operation[46][29]) ;
              //$display("@%0t LEE: Received final operation event for 46,29\n", $time);
            end
            begin
              @(final_operation[46][30]) ;
              //$display("@%0t LEE: Received final operation event for 46,30\n", $time);
            end
            begin
              @(final_operation[46][31]) ;
              //$display("@%0t LEE: Received final operation event for 46,31\n", $time);
            end

            begin
              @(final_operation[47][0]) ;
              //$display("@%0t LEE: Received final operation event for 47,0\n", $time);
            end
            begin
              @(final_operation[47][1]) ;
              //$display("@%0t LEE: Received final operation event for 47,1\n", $time);
            end
            begin
              @(final_operation[47][2]) ;
              //$display("@%0t LEE: Received final operation event for 47,2\n", $time);
            end
            begin
              @(final_operation[47][3]) ;
              //$display("@%0t LEE: Received final operation event for 47,3\n", $time);
            end
            begin
              @(final_operation[47][4]) ;
              //$display("@%0t LEE: Received final operation event for 47,4\n", $time);
            end
            begin
              @(final_operation[47][5]) ;
              //$display("@%0t LEE: Received final operation event for 47,5\n", $time);
            end
            begin
              @(final_operation[47][6]) ;
              //$display("@%0t LEE: Received final operation event for 47,6\n", $time);
            end
            begin
              @(final_operation[47][7]) ;
              //$display("@%0t LEE: Received final operation event for 47,7\n", $time);
            end
            begin
              @(final_operation[47][8]) ;
              //$display("@%0t LEE: Received final operation event for 47,8\n", $time);
            end
            begin
              @(final_operation[47][9]) ;
              //$display("@%0t LEE: Received final operation event for 47,9\n", $time);
            end
            begin
              @(final_operation[47][10]) ;
              //$display("@%0t LEE: Received final operation event for 47,10\n", $time);
            end
            begin
              @(final_operation[47][11]) ;
              //$display("@%0t LEE: Received final operation event for 47,11\n", $time);
            end
            begin
              @(final_operation[47][12]) ;
              //$display("@%0t LEE: Received final operation event for 47,12\n", $time);
            end
            begin
              @(final_operation[47][13]) ;
              //$display("@%0t LEE: Received final operation event for 47,13\n", $time);
            end
            begin
              @(final_operation[47][14]) ;
              //$display("@%0t LEE: Received final operation event for 47,14\n", $time);
            end
            begin
              @(final_operation[47][15]) ;
              //$display("@%0t LEE: Received final operation event for 47,15\n", $time);
            end
            begin
              @(final_operation[47][16]) ;
              //$display("@%0t LEE: Received final operation event for 47,16\n", $time);
            end
            begin
              @(final_operation[47][17]) ;
              //$display("@%0t LEE: Received final operation event for 47,17\n", $time);
            end
            begin
              @(final_operation[47][18]) ;
              //$display("@%0t LEE: Received final operation event for 47,18\n", $time);
            end
            begin
              @(final_operation[47][19]) ;
              //$display("@%0t LEE: Received final operation event for 47,19\n", $time);
            end
            begin
              @(final_operation[47][20]) ;
              //$display("@%0t LEE: Received final operation event for 47,20\n", $time);
            end
            begin
              @(final_operation[47][21]) ;
              //$display("@%0t LEE: Received final operation event for 47,21\n", $time);
            end
            begin
              @(final_operation[47][22]) ;
              //$display("@%0t LEE: Received final operation event for 47,22\n", $time);
            end
            begin
              @(final_operation[47][23]) ;
              //$display("@%0t LEE: Received final operation event for 47,23\n", $time);
            end
            begin
              @(final_operation[47][24]) ;
              //$display("@%0t LEE: Received final operation event for 47,24\n", $time);
            end
            begin
              @(final_operation[47][25]) ;
              //$display("@%0t LEE: Received final operation event for 47,25\n", $time);
            end
            begin
              @(final_operation[47][26]) ;
              //$display("@%0t LEE: Received final operation event for 47,26\n", $time);
            end
            begin
              @(final_operation[47][27]) ;
              //$display("@%0t LEE: Received final operation event for 47,27\n", $time);
            end
            begin
              @(final_operation[47][28]) ;
              //$display("@%0t LEE: Received final operation event for 47,28\n", $time);
            end
            begin
              @(final_operation[47][29]) ;
              //$display("@%0t LEE: Received final operation event for 47,29\n", $time);
            end
            begin
              @(final_operation[47][30]) ;
              //$display("@%0t LEE: Received final operation event for 47,30\n", $time);
            end
            begin
              @(final_operation[47][31]) ;
              //$display("@%0t LEE: Received final operation event for 47,31\n", $time);
            end

            begin
              @(final_operation[48][0]) ;
              //$display("@%0t LEE: Received final operation event for 48,0\n", $time);
            end
            begin
              @(final_operation[48][1]) ;
              //$display("@%0t LEE: Received final operation event for 48,1\n", $time);
            end
            begin
              @(final_operation[48][2]) ;
              //$display("@%0t LEE: Received final operation event for 48,2\n", $time);
            end
            begin
              @(final_operation[48][3]) ;
              //$display("@%0t LEE: Received final operation event for 48,3\n", $time);
            end
            begin
              @(final_operation[48][4]) ;
              //$display("@%0t LEE: Received final operation event for 48,4\n", $time);
            end
            begin
              @(final_operation[48][5]) ;
              //$display("@%0t LEE: Received final operation event for 48,5\n", $time);
            end
            begin
              @(final_operation[48][6]) ;
              //$display("@%0t LEE: Received final operation event for 48,6\n", $time);
            end
            begin
              @(final_operation[48][7]) ;
              //$display("@%0t LEE: Received final operation event for 48,7\n", $time);
            end
            begin
              @(final_operation[48][8]) ;
              //$display("@%0t LEE: Received final operation event for 48,8\n", $time);
            end
            begin
              @(final_operation[48][9]) ;
              //$display("@%0t LEE: Received final operation event for 48,9\n", $time);
            end
            begin
              @(final_operation[48][10]) ;
              //$display("@%0t LEE: Received final operation event for 48,10\n", $time);
            end
            begin
              @(final_operation[48][11]) ;
              //$display("@%0t LEE: Received final operation event for 48,11\n", $time);
            end
            begin
              @(final_operation[48][12]) ;
              //$display("@%0t LEE: Received final operation event for 48,12\n", $time);
            end
            begin
              @(final_operation[48][13]) ;
              //$display("@%0t LEE: Received final operation event for 48,13\n", $time);
            end
            begin
              @(final_operation[48][14]) ;
              //$display("@%0t LEE: Received final operation event for 48,14\n", $time);
            end
            begin
              @(final_operation[48][15]) ;
              //$display("@%0t LEE: Received final operation event for 48,15\n", $time);
            end
            begin
              @(final_operation[48][16]) ;
              //$display("@%0t LEE: Received final operation event for 48,16\n", $time);
            end
            begin
              @(final_operation[48][17]) ;
              //$display("@%0t LEE: Received final operation event for 48,17\n", $time);
            end
            begin
              @(final_operation[48][18]) ;
              //$display("@%0t LEE: Received final operation event for 48,18\n", $time);
            end
            begin
              @(final_operation[48][19]) ;
              //$display("@%0t LEE: Received final operation event for 48,19\n", $time);
            end
            begin
              @(final_operation[48][20]) ;
              //$display("@%0t LEE: Received final operation event for 48,20\n", $time);
            end
            begin
              @(final_operation[48][21]) ;
              //$display("@%0t LEE: Received final operation event for 48,21\n", $time);
            end
            begin
              @(final_operation[48][22]) ;
              //$display("@%0t LEE: Received final operation event for 48,22\n", $time);
            end
            begin
              @(final_operation[48][23]) ;
              //$display("@%0t LEE: Received final operation event for 48,23\n", $time);
            end
            begin
              @(final_operation[48][24]) ;
              //$display("@%0t LEE: Received final operation event for 48,24\n", $time);
            end
            begin
              @(final_operation[48][25]) ;
              //$display("@%0t LEE: Received final operation event for 48,25\n", $time);
            end
            begin
              @(final_operation[48][26]) ;
              //$display("@%0t LEE: Received final operation event for 48,26\n", $time);
            end
            begin
              @(final_operation[48][27]) ;
              //$display("@%0t LEE: Received final operation event for 48,27\n", $time);
            end
            begin
              @(final_operation[48][28]) ;
              //$display("@%0t LEE: Received final operation event for 48,28\n", $time);
            end
            begin
              @(final_operation[48][29]) ;
              //$display("@%0t LEE: Received final operation event for 48,29\n", $time);
            end
            begin
              @(final_operation[48][30]) ;
              //$display("@%0t LEE: Received final operation event for 48,30\n", $time);
            end
            begin
              @(final_operation[48][31]) ;
              //$display("@%0t LEE: Received final operation event for 48,31\n", $time);
            end

            begin
              @(final_operation[49][0]) ;
              //$display("@%0t LEE: Received final operation event for 49,0\n", $time);
            end
            begin
              @(final_operation[49][1]) ;
              //$display("@%0t LEE: Received final operation event for 49,1\n", $time);
            end
            begin
              @(final_operation[49][2]) ;
              //$display("@%0t LEE: Received final operation event for 49,2\n", $time);
            end
            begin
              @(final_operation[49][3]) ;
              //$display("@%0t LEE: Received final operation event for 49,3\n", $time);
            end
            begin
              @(final_operation[49][4]) ;
              //$display("@%0t LEE: Received final operation event for 49,4\n", $time);
            end
            begin
              @(final_operation[49][5]) ;
              //$display("@%0t LEE: Received final operation event for 49,5\n", $time);
            end
            begin
              @(final_operation[49][6]) ;
              //$display("@%0t LEE: Received final operation event for 49,6\n", $time);
            end
            begin
              @(final_operation[49][7]) ;
              //$display("@%0t LEE: Received final operation event for 49,7\n", $time);
            end
            begin
              @(final_operation[49][8]) ;
              //$display("@%0t LEE: Received final operation event for 49,8\n", $time);
            end
            begin
              @(final_operation[49][9]) ;
              //$display("@%0t LEE: Received final operation event for 49,9\n", $time);
            end
            begin
              @(final_operation[49][10]) ;
              //$display("@%0t LEE: Received final operation event for 49,10\n", $time);
            end
            begin
              @(final_operation[49][11]) ;
              //$display("@%0t LEE: Received final operation event for 49,11\n", $time);
            end
            begin
              @(final_operation[49][12]) ;
              //$display("@%0t LEE: Received final operation event for 49,12\n", $time);
            end
            begin
              @(final_operation[49][13]) ;
              //$display("@%0t LEE: Received final operation event for 49,13\n", $time);
            end
            begin
              @(final_operation[49][14]) ;
              //$display("@%0t LEE: Received final operation event for 49,14\n", $time);
            end
            begin
              @(final_operation[49][15]) ;
              //$display("@%0t LEE: Received final operation event for 49,15\n", $time);
            end
            begin
              @(final_operation[49][16]) ;
              //$display("@%0t LEE: Received final operation event for 49,16\n", $time);
            end
            begin
              @(final_operation[49][17]) ;
              //$display("@%0t LEE: Received final operation event for 49,17\n", $time);
            end
            begin
              @(final_operation[49][18]) ;
              //$display("@%0t LEE: Received final operation event for 49,18\n", $time);
            end
            begin
              @(final_operation[49][19]) ;
              //$display("@%0t LEE: Received final operation event for 49,19\n", $time);
            end
            begin
              @(final_operation[49][20]) ;
              //$display("@%0t LEE: Received final operation event for 49,20\n", $time);
            end
            begin
              @(final_operation[49][21]) ;
              //$display("@%0t LEE: Received final operation event for 49,21\n", $time);
            end
            begin
              @(final_operation[49][22]) ;
              //$display("@%0t LEE: Received final operation event for 49,22\n", $time);
            end
            begin
              @(final_operation[49][23]) ;
              //$display("@%0t LEE: Received final operation event for 49,23\n", $time);
            end
            begin
              @(final_operation[49][24]) ;
              //$display("@%0t LEE: Received final operation event for 49,24\n", $time);
            end
            begin
              @(final_operation[49][25]) ;
              //$display("@%0t LEE: Received final operation event for 49,25\n", $time);
            end
            begin
              @(final_operation[49][26]) ;
              //$display("@%0t LEE: Received final operation event for 49,26\n", $time);
            end
            begin
              @(final_operation[49][27]) ;
              //$display("@%0t LEE: Received final operation event for 49,27\n", $time);
            end
            begin
              @(final_operation[49][28]) ;
              //$display("@%0t LEE: Received final operation event for 49,28\n", $time);
            end
            begin
              @(final_operation[49][29]) ;
              //$display("@%0t LEE: Received final operation event for 49,29\n", $time);
            end
            begin
              @(final_operation[49][30]) ;
              //$display("@%0t LEE: Received final operation event for 49,30\n", $time);
            end
            begin
              @(final_operation[49][31]) ;
              //$display("@%0t LEE: Received final operation event for 49,31\n", $time);
            end

            begin
              @(final_operation[50][0]) ;
              //$display("@%0t LEE: Received final operation event for 50,0\n", $time);
            end
            begin
              @(final_operation[50][1]) ;
              //$display("@%0t LEE: Received final operation event for 50,1\n", $time);
            end
            begin
              @(final_operation[50][2]) ;
              //$display("@%0t LEE: Received final operation event for 50,2\n", $time);
            end
            begin
              @(final_operation[50][3]) ;
              //$display("@%0t LEE: Received final operation event for 50,3\n", $time);
            end
            begin
              @(final_operation[50][4]) ;
              //$display("@%0t LEE: Received final operation event for 50,4\n", $time);
            end
            begin
              @(final_operation[50][5]) ;
              //$display("@%0t LEE: Received final operation event for 50,5\n", $time);
            end
            begin
              @(final_operation[50][6]) ;
              //$display("@%0t LEE: Received final operation event for 50,6\n", $time);
            end
            begin
              @(final_operation[50][7]) ;
              //$display("@%0t LEE: Received final operation event for 50,7\n", $time);
            end
            begin
              @(final_operation[50][8]) ;
              //$display("@%0t LEE: Received final operation event for 50,8\n", $time);
            end
            begin
              @(final_operation[50][9]) ;
              //$display("@%0t LEE: Received final operation event for 50,9\n", $time);
            end
            begin
              @(final_operation[50][10]) ;
              //$display("@%0t LEE: Received final operation event for 50,10\n", $time);
            end
            begin
              @(final_operation[50][11]) ;
              //$display("@%0t LEE: Received final operation event for 50,11\n", $time);
            end
            begin
              @(final_operation[50][12]) ;
              //$display("@%0t LEE: Received final operation event for 50,12\n", $time);
            end
            begin
              @(final_operation[50][13]) ;
              //$display("@%0t LEE: Received final operation event for 50,13\n", $time);
            end
            begin
              @(final_operation[50][14]) ;
              //$display("@%0t LEE: Received final operation event for 50,14\n", $time);
            end
            begin
              @(final_operation[50][15]) ;
              //$display("@%0t LEE: Received final operation event for 50,15\n", $time);
            end
            begin
              @(final_operation[50][16]) ;
              //$display("@%0t LEE: Received final operation event for 50,16\n", $time);
            end
            begin
              @(final_operation[50][17]) ;
              //$display("@%0t LEE: Received final operation event for 50,17\n", $time);
            end
            begin
              @(final_operation[50][18]) ;
              //$display("@%0t LEE: Received final operation event for 50,18\n", $time);
            end
            begin
              @(final_operation[50][19]) ;
              //$display("@%0t LEE: Received final operation event for 50,19\n", $time);
            end
            begin
              @(final_operation[50][20]) ;
              //$display("@%0t LEE: Received final operation event for 50,20\n", $time);
            end
            begin
              @(final_operation[50][21]) ;
              //$display("@%0t LEE: Received final operation event for 50,21\n", $time);
            end
            begin
              @(final_operation[50][22]) ;
              //$display("@%0t LEE: Received final operation event for 50,22\n", $time);
            end
            begin
              @(final_operation[50][23]) ;
              //$display("@%0t LEE: Received final operation event for 50,23\n", $time);
            end
            begin
              @(final_operation[50][24]) ;
              //$display("@%0t LEE: Received final operation event for 50,24\n", $time);
            end
            begin
              @(final_operation[50][25]) ;
              //$display("@%0t LEE: Received final operation event for 50,25\n", $time);
            end
            begin
              @(final_operation[50][26]) ;
              //$display("@%0t LEE: Received final operation event for 50,26\n", $time);
            end
            begin
              @(final_operation[50][27]) ;
              //$display("@%0t LEE: Received final operation event for 50,27\n", $time);
            end
            begin
              @(final_operation[50][28]) ;
              //$display("@%0t LEE: Received final operation event for 50,28\n", $time);
            end
            begin
              @(final_operation[50][29]) ;
              //$display("@%0t LEE: Received final operation event for 50,29\n", $time);
            end
            begin
              @(final_operation[50][30]) ;
              //$display("@%0t LEE: Received final operation event for 50,30\n", $time);
            end
            begin
              @(final_operation[50][31]) ;
              //$display("@%0t LEE: Received final operation event for 50,31\n", $time);
            end

            begin
              @(final_operation[51][0]) ;
              //$display("@%0t LEE: Received final operation event for 51,0\n", $time);
            end
            begin
              @(final_operation[51][1]) ;
              //$display("@%0t LEE: Received final operation event for 51,1\n", $time);
            end
            begin
              @(final_operation[51][2]) ;
              //$display("@%0t LEE: Received final operation event for 51,2\n", $time);
            end
            begin
              @(final_operation[51][3]) ;
              //$display("@%0t LEE: Received final operation event for 51,3\n", $time);
            end
            begin
              @(final_operation[51][4]) ;
              //$display("@%0t LEE: Received final operation event for 51,4\n", $time);
            end
            begin
              @(final_operation[51][5]) ;
              //$display("@%0t LEE: Received final operation event for 51,5\n", $time);
            end
            begin
              @(final_operation[51][6]) ;
              //$display("@%0t LEE: Received final operation event for 51,6\n", $time);
            end
            begin
              @(final_operation[51][7]) ;
              //$display("@%0t LEE: Received final operation event for 51,7\n", $time);
            end
            begin
              @(final_operation[51][8]) ;
              //$display("@%0t LEE: Received final operation event for 51,8\n", $time);
            end
            begin
              @(final_operation[51][9]) ;
              //$display("@%0t LEE: Received final operation event for 51,9\n", $time);
            end
            begin
              @(final_operation[51][10]) ;
              //$display("@%0t LEE: Received final operation event for 51,10\n", $time);
            end
            begin
              @(final_operation[51][11]) ;
              //$display("@%0t LEE: Received final operation event for 51,11\n", $time);
            end
            begin
              @(final_operation[51][12]) ;
              //$display("@%0t LEE: Received final operation event for 51,12\n", $time);
            end
            begin
              @(final_operation[51][13]) ;
              //$display("@%0t LEE: Received final operation event for 51,13\n", $time);
            end
            begin
              @(final_operation[51][14]) ;
              //$display("@%0t LEE: Received final operation event for 51,14\n", $time);
            end
            begin
              @(final_operation[51][15]) ;
              //$display("@%0t LEE: Received final operation event for 51,15\n", $time);
            end
            begin
              @(final_operation[51][16]) ;
              //$display("@%0t LEE: Received final operation event for 51,16\n", $time);
            end
            begin
              @(final_operation[51][17]) ;
              //$display("@%0t LEE: Received final operation event for 51,17\n", $time);
            end
            begin
              @(final_operation[51][18]) ;
              //$display("@%0t LEE: Received final operation event for 51,18\n", $time);
            end
            begin
              @(final_operation[51][19]) ;
              //$display("@%0t LEE: Received final operation event for 51,19\n", $time);
            end
            begin
              @(final_operation[51][20]) ;
              //$display("@%0t LEE: Received final operation event for 51,20\n", $time);
            end
            begin
              @(final_operation[51][21]) ;
              //$display("@%0t LEE: Received final operation event for 51,21\n", $time);
            end
            begin
              @(final_operation[51][22]) ;
              //$display("@%0t LEE: Received final operation event for 51,22\n", $time);
            end
            begin
              @(final_operation[51][23]) ;
              //$display("@%0t LEE: Received final operation event for 51,23\n", $time);
            end
            begin
              @(final_operation[51][24]) ;
              //$display("@%0t LEE: Received final operation event for 51,24\n", $time);
            end
            begin
              @(final_operation[51][25]) ;
              //$display("@%0t LEE: Received final operation event for 51,25\n", $time);
            end
            begin
              @(final_operation[51][26]) ;
              //$display("@%0t LEE: Received final operation event for 51,26\n", $time);
            end
            begin
              @(final_operation[51][27]) ;
              //$display("@%0t LEE: Received final operation event for 51,27\n", $time);
            end
            begin
              @(final_operation[51][28]) ;
              //$display("@%0t LEE: Received final operation event for 51,28\n", $time);
            end
            begin
              @(final_operation[51][29]) ;
              //$display("@%0t LEE: Received final operation event for 51,29\n", $time);
            end
            begin
              @(final_operation[51][30]) ;
              //$display("@%0t LEE: Received final operation event for 51,30\n", $time);
            end
            begin
              @(final_operation[51][31]) ;
              //$display("@%0t LEE: Received final operation event for 51,31\n", $time);
            end

            begin
              @(final_operation[52][0]) ;
              //$display("@%0t LEE: Received final operation event for 52,0\n", $time);
            end
            begin
              @(final_operation[52][1]) ;
              //$display("@%0t LEE: Received final operation event for 52,1\n", $time);
            end
            begin
              @(final_operation[52][2]) ;
              //$display("@%0t LEE: Received final operation event for 52,2\n", $time);
            end
            begin
              @(final_operation[52][3]) ;
              //$display("@%0t LEE: Received final operation event for 52,3\n", $time);
            end
            begin
              @(final_operation[52][4]) ;
              //$display("@%0t LEE: Received final operation event for 52,4\n", $time);
            end
            begin
              @(final_operation[52][5]) ;
              //$display("@%0t LEE: Received final operation event for 52,5\n", $time);
            end
            begin
              @(final_operation[52][6]) ;
              //$display("@%0t LEE: Received final operation event for 52,6\n", $time);
            end
            begin
              @(final_operation[52][7]) ;
              //$display("@%0t LEE: Received final operation event for 52,7\n", $time);
            end
            begin
              @(final_operation[52][8]) ;
              //$display("@%0t LEE: Received final operation event for 52,8\n", $time);
            end
            begin
              @(final_operation[52][9]) ;
              //$display("@%0t LEE: Received final operation event for 52,9\n", $time);
            end
            begin
              @(final_operation[52][10]) ;
              //$display("@%0t LEE: Received final operation event for 52,10\n", $time);
            end
            begin
              @(final_operation[52][11]) ;
              //$display("@%0t LEE: Received final operation event for 52,11\n", $time);
            end
            begin
              @(final_operation[52][12]) ;
              //$display("@%0t LEE: Received final operation event for 52,12\n", $time);
            end
            begin
              @(final_operation[52][13]) ;
              //$display("@%0t LEE: Received final operation event for 52,13\n", $time);
            end
            begin
              @(final_operation[52][14]) ;
              //$display("@%0t LEE: Received final operation event for 52,14\n", $time);
            end
            begin
              @(final_operation[52][15]) ;
              //$display("@%0t LEE: Received final operation event for 52,15\n", $time);
            end
            begin
              @(final_operation[52][16]) ;
              //$display("@%0t LEE: Received final operation event for 52,16\n", $time);
            end
            begin
              @(final_operation[52][17]) ;
              //$display("@%0t LEE: Received final operation event for 52,17\n", $time);
            end
            begin
              @(final_operation[52][18]) ;
              //$display("@%0t LEE: Received final operation event for 52,18\n", $time);
            end
            begin
              @(final_operation[52][19]) ;
              //$display("@%0t LEE: Received final operation event for 52,19\n", $time);
            end
            begin
              @(final_operation[52][20]) ;
              //$display("@%0t LEE: Received final operation event for 52,20\n", $time);
            end
            begin
              @(final_operation[52][21]) ;
              //$display("@%0t LEE: Received final operation event for 52,21\n", $time);
            end
            begin
              @(final_operation[52][22]) ;
              //$display("@%0t LEE: Received final operation event for 52,22\n", $time);
            end
            begin
              @(final_operation[52][23]) ;
              //$display("@%0t LEE: Received final operation event for 52,23\n", $time);
            end
            begin
              @(final_operation[52][24]) ;
              //$display("@%0t LEE: Received final operation event for 52,24\n", $time);
            end
            begin
              @(final_operation[52][25]) ;
              //$display("@%0t LEE: Received final operation event for 52,25\n", $time);
            end
            begin
              @(final_operation[52][26]) ;
              //$display("@%0t LEE: Received final operation event for 52,26\n", $time);
            end
            begin
              @(final_operation[52][27]) ;
              //$display("@%0t LEE: Received final operation event for 52,27\n", $time);
            end
            begin
              @(final_operation[52][28]) ;
              //$display("@%0t LEE: Received final operation event for 52,28\n", $time);
            end
            begin
              @(final_operation[52][29]) ;
              //$display("@%0t LEE: Received final operation event for 52,29\n", $time);
            end
            begin
              @(final_operation[52][30]) ;
              //$display("@%0t LEE: Received final operation event for 52,30\n", $time);
            end
            begin
              @(final_operation[52][31]) ;
              //$display("@%0t LEE: Received final operation event for 52,31\n", $time);
            end

            begin
              @(final_operation[53][0]) ;
              //$display("@%0t LEE: Received final operation event for 53,0\n", $time);
            end
            begin
              @(final_operation[53][1]) ;
              //$display("@%0t LEE: Received final operation event for 53,1\n", $time);
            end
            begin
              @(final_operation[53][2]) ;
              //$display("@%0t LEE: Received final operation event for 53,2\n", $time);
            end
            begin
              @(final_operation[53][3]) ;
              //$display("@%0t LEE: Received final operation event for 53,3\n", $time);
            end
            begin
              @(final_operation[53][4]) ;
              //$display("@%0t LEE: Received final operation event for 53,4\n", $time);
            end
            begin
              @(final_operation[53][5]) ;
              //$display("@%0t LEE: Received final operation event for 53,5\n", $time);
            end
            begin
              @(final_operation[53][6]) ;
              //$display("@%0t LEE: Received final operation event for 53,6\n", $time);
            end
            begin
              @(final_operation[53][7]) ;
              //$display("@%0t LEE: Received final operation event for 53,7\n", $time);
            end
            begin
              @(final_operation[53][8]) ;
              //$display("@%0t LEE: Received final operation event for 53,8\n", $time);
            end
            begin
              @(final_operation[53][9]) ;
              //$display("@%0t LEE: Received final operation event for 53,9\n", $time);
            end
            begin
              @(final_operation[53][10]) ;
              //$display("@%0t LEE: Received final operation event for 53,10\n", $time);
            end
            begin
              @(final_operation[53][11]) ;
              //$display("@%0t LEE: Received final operation event for 53,11\n", $time);
            end
            begin
              @(final_operation[53][12]) ;
              //$display("@%0t LEE: Received final operation event for 53,12\n", $time);
            end
            begin
              @(final_operation[53][13]) ;
              //$display("@%0t LEE: Received final operation event for 53,13\n", $time);
            end
            begin
              @(final_operation[53][14]) ;
              //$display("@%0t LEE: Received final operation event for 53,14\n", $time);
            end
            begin
              @(final_operation[53][15]) ;
              //$display("@%0t LEE: Received final operation event for 53,15\n", $time);
            end
            begin
              @(final_operation[53][16]) ;
              //$display("@%0t LEE: Received final operation event for 53,16\n", $time);
            end
            begin
              @(final_operation[53][17]) ;
              //$display("@%0t LEE: Received final operation event for 53,17\n", $time);
            end
            begin
              @(final_operation[53][18]) ;
              //$display("@%0t LEE: Received final operation event for 53,18\n", $time);
            end
            begin
              @(final_operation[53][19]) ;
              //$display("@%0t LEE: Received final operation event for 53,19\n", $time);
            end
            begin
              @(final_operation[53][20]) ;
              //$display("@%0t LEE: Received final operation event for 53,20\n", $time);
            end
            begin
              @(final_operation[53][21]) ;
              //$display("@%0t LEE: Received final operation event for 53,21\n", $time);
            end
            begin
              @(final_operation[53][22]) ;
              //$display("@%0t LEE: Received final operation event for 53,22\n", $time);
            end
            begin
              @(final_operation[53][23]) ;
              //$display("@%0t LEE: Received final operation event for 53,23\n", $time);
            end
            begin
              @(final_operation[53][24]) ;
              //$display("@%0t LEE: Received final operation event for 53,24\n", $time);
            end
            begin
              @(final_operation[53][25]) ;
              //$display("@%0t LEE: Received final operation event for 53,25\n", $time);
            end
            begin
              @(final_operation[53][26]) ;
              //$display("@%0t LEE: Received final operation event for 53,26\n", $time);
            end
            begin
              @(final_operation[53][27]) ;
              //$display("@%0t LEE: Received final operation event for 53,27\n", $time);
            end
            begin
              @(final_operation[53][28]) ;
              //$display("@%0t LEE: Received final operation event for 53,28\n", $time);
            end
            begin
              @(final_operation[53][29]) ;
              //$display("@%0t LEE: Received final operation event for 53,29\n", $time);
            end
            begin
              @(final_operation[53][30]) ;
              //$display("@%0t LEE: Received final operation event for 53,30\n", $time);
            end
            begin
              @(final_operation[53][31]) ;
              //$display("@%0t LEE: Received final operation event for 53,31\n", $time);
            end

            begin
              @(final_operation[54][0]) ;
              //$display("@%0t LEE: Received final operation event for 54,0\n", $time);
            end
            begin
              @(final_operation[54][1]) ;
              //$display("@%0t LEE: Received final operation event for 54,1\n", $time);
            end
            begin
              @(final_operation[54][2]) ;
              //$display("@%0t LEE: Received final operation event for 54,2\n", $time);
            end
            begin
              @(final_operation[54][3]) ;
              //$display("@%0t LEE: Received final operation event for 54,3\n", $time);
            end
            begin
              @(final_operation[54][4]) ;
              //$display("@%0t LEE: Received final operation event for 54,4\n", $time);
            end
            begin
              @(final_operation[54][5]) ;
              //$display("@%0t LEE: Received final operation event for 54,5\n", $time);
            end
            begin
              @(final_operation[54][6]) ;
              //$display("@%0t LEE: Received final operation event for 54,6\n", $time);
            end
            begin
              @(final_operation[54][7]) ;
              //$display("@%0t LEE: Received final operation event for 54,7\n", $time);
            end
            begin
              @(final_operation[54][8]) ;
              //$display("@%0t LEE: Received final operation event for 54,8\n", $time);
            end
            begin
              @(final_operation[54][9]) ;
              //$display("@%0t LEE: Received final operation event for 54,9\n", $time);
            end
            begin
              @(final_operation[54][10]) ;
              //$display("@%0t LEE: Received final operation event for 54,10\n", $time);
            end
            begin
              @(final_operation[54][11]) ;
              //$display("@%0t LEE: Received final operation event for 54,11\n", $time);
            end
            begin
              @(final_operation[54][12]) ;
              //$display("@%0t LEE: Received final operation event for 54,12\n", $time);
            end
            begin
              @(final_operation[54][13]) ;
              //$display("@%0t LEE: Received final operation event for 54,13\n", $time);
            end
            begin
              @(final_operation[54][14]) ;
              //$display("@%0t LEE: Received final operation event for 54,14\n", $time);
            end
            begin
              @(final_operation[54][15]) ;
              //$display("@%0t LEE: Received final operation event for 54,15\n", $time);
            end
            begin
              @(final_operation[54][16]) ;
              //$display("@%0t LEE: Received final operation event for 54,16\n", $time);
            end
            begin
              @(final_operation[54][17]) ;
              //$display("@%0t LEE: Received final operation event for 54,17\n", $time);
            end
            begin
              @(final_operation[54][18]) ;
              //$display("@%0t LEE: Received final operation event for 54,18\n", $time);
            end
            begin
              @(final_operation[54][19]) ;
              //$display("@%0t LEE: Received final operation event for 54,19\n", $time);
            end
            begin
              @(final_operation[54][20]) ;
              //$display("@%0t LEE: Received final operation event for 54,20\n", $time);
            end
            begin
              @(final_operation[54][21]) ;
              //$display("@%0t LEE: Received final operation event for 54,21\n", $time);
            end
            begin
              @(final_operation[54][22]) ;
              //$display("@%0t LEE: Received final operation event for 54,22\n", $time);
            end
            begin
              @(final_operation[54][23]) ;
              //$display("@%0t LEE: Received final operation event for 54,23\n", $time);
            end
            begin
              @(final_operation[54][24]) ;
              //$display("@%0t LEE: Received final operation event for 54,24\n", $time);
            end
            begin
              @(final_operation[54][25]) ;
              //$display("@%0t LEE: Received final operation event for 54,25\n", $time);
            end
            begin
              @(final_operation[54][26]) ;
              //$display("@%0t LEE: Received final operation event for 54,26\n", $time);
            end
            begin
              @(final_operation[54][27]) ;
              //$display("@%0t LEE: Received final operation event for 54,27\n", $time);
            end
            begin
              @(final_operation[54][28]) ;
              //$display("@%0t LEE: Received final operation event for 54,28\n", $time);
            end
            begin
              @(final_operation[54][29]) ;
              //$display("@%0t LEE: Received final operation event for 54,29\n", $time);
            end
            begin
              @(final_operation[54][30]) ;
              //$display("@%0t LEE: Received final operation event for 54,30\n", $time);
            end
            begin
              @(final_operation[54][31]) ;
              //$display("@%0t LEE: Received final operation event for 54,31\n", $time);
            end

            begin
              @(final_operation[55][0]) ;
              //$display("@%0t LEE: Received final operation event for 55,0\n", $time);
            end
            begin
              @(final_operation[55][1]) ;
              //$display("@%0t LEE: Received final operation event for 55,1\n", $time);
            end
            begin
              @(final_operation[55][2]) ;
              //$display("@%0t LEE: Received final operation event for 55,2\n", $time);
            end
            begin
              @(final_operation[55][3]) ;
              //$display("@%0t LEE: Received final operation event for 55,3\n", $time);
            end
            begin
              @(final_operation[55][4]) ;
              //$display("@%0t LEE: Received final operation event for 55,4\n", $time);
            end
            begin
              @(final_operation[55][5]) ;
              //$display("@%0t LEE: Received final operation event for 55,5\n", $time);
            end
            begin
              @(final_operation[55][6]) ;
              //$display("@%0t LEE: Received final operation event for 55,6\n", $time);
            end
            begin
              @(final_operation[55][7]) ;
              //$display("@%0t LEE: Received final operation event for 55,7\n", $time);
            end
            begin
              @(final_operation[55][8]) ;
              //$display("@%0t LEE: Received final operation event for 55,8\n", $time);
            end
            begin
              @(final_operation[55][9]) ;
              //$display("@%0t LEE: Received final operation event for 55,9\n", $time);
            end
            begin
              @(final_operation[55][10]) ;
              //$display("@%0t LEE: Received final operation event for 55,10\n", $time);
            end
            begin
              @(final_operation[55][11]) ;
              //$display("@%0t LEE: Received final operation event for 55,11\n", $time);
            end
            begin
              @(final_operation[55][12]) ;
              //$display("@%0t LEE: Received final operation event for 55,12\n", $time);
            end
            begin
              @(final_operation[55][13]) ;
              //$display("@%0t LEE: Received final operation event for 55,13\n", $time);
            end
            begin
              @(final_operation[55][14]) ;
              //$display("@%0t LEE: Received final operation event for 55,14\n", $time);
            end
            begin
              @(final_operation[55][15]) ;
              //$display("@%0t LEE: Received final operation event for 55,15\n", $time);
            end
            begin
              @(final_operation[55][16]) ;
              //$display("@%0t LEE: Received final operation event for 55,16\n", $time);
            end
            begin
              @(final_operation[55][17]) ;
              //$display("@%0t LEE: Received final operation event for 55,17\n", $time);
            end
            begin
              @(final_operation[55][18]) ;
              //$display("@%0t LEE: Received final operation event for 55,18\n", $time);
            end
            begin
              @(final_operation[55][19]) ;
              //$display("@%0t LEE: Received final operation event for 55,19\n", $time);
            end
            begin
              @(final_operation[55][20]) ;
              //$display("@%0t LEE: Received final operation event for 55,20\n", $time);
            end
            begin
              @(final_operation[55][21]) ;
              //$display("@%0t LEE: Received final operation event for 55,21\n", $time);
            end
            begin
              @(final_operation[55][22]) ;
              //$display("@%0t LEE: Received final operation event for 55,22\n", $time);
            end
            begin
              @(final_operation[55][23]) ;
              //$display("@%0t LEE: Received final operation event for 55,23\n", $time);
            end
            begin
              @(final_operation[55][24]) ;
              //$display("@%0t LEE: Received final operation event for 55,24\n", $time);
            end
            begin
              @(final_operation[55][25]) ;
              //$display("@%0t LEE: Received final operation event for 55,25\n", $time);
            end
            begin
              @(final_operation[55][26]) ;
              //$display("@%0t LEE: Received final operation event for 55,26\n", $time);
            end
            begin
              @(final_operation[55][27]) ;
              //$display("@%0t LEE: Received final operation event for 55,27\n", $time);
            end
            begin
              @(final_operation[55][28]) ;
              //$display("@%0t LEE: Received final operation event for 55,28\n", $time);
            end
            begin
              @(final_operation[55][29]) ;
              //$display("@%0t LEE: Received final operation event for 55,29\n", $time);
            end
            begin
              @(final_operation[55][30]) ;
              //$display("@%0t LEE: Received final operation event for 55,30\n", $time);
            end
            begin
              @(final_operation[55][31]) ;
              //$display("@%0t LEE: Received final operation event for 55,31\n", $time);
            end

            begin
              @(final_operation[56][0]) ;
              //$display("@%0t LEE: Received final operation event for 56,0\n", $time);
            end
            begin
              @(final_operation[56][1]) ;
              //$display("@%0t LEE: Received final operation event for 56,1\n", $time);
            end
            begin
              @(final_operation[56][2]) ;
              //$display("@%0t LEE: Received final operation event for 56,2\n", $time);
            end
            begin
              @(final_operation[56][3]) ;
              //$display("@%0t LEE: Received final operation event for 56,3\n", $time);
            end
            begin
              @(final_operation[56][4]) ;
              //$display("@%0t LEE: Received final operation event for 56,4\n", $time);
            end
            begin
              @(final_operation[56][5]) ;
              //$display("@%0t LEE: Received final operation event for 56,5\n", $time);
            end
            begin
              @(final_operation[56][6]) ;
              //$display("@%0t LEE: Received final operation event for 56,6\n", $time);
            end
            begin
              @(final_operation[56][7]) ;
              //$display("@%0t LEE: Received final operation event for 56,7\n", $time);
            end
            begin
              @(final_operation[56][8]) ;
              //$display("@%0t LEE: Received final operation event for 56,8\n", $time);
            end
            begin
              @(final_operation[56][9]) ;
              //$display("@%0t LEE: Received final operation event for 56,9\n", $time);
            end
            begin
              @(final_operation[56][10]) ;
              //$display("@%0t LEE: Received final operation event for 56,10\n", $time);
            end
            begin
              @(final_operation[56][11]) ;
              //$display("@%0t LEE: Received final operation event for 56,11\n", $time);
            end
            begin
              @(final_operation[56][12]) ;
              //$display("@%0t LEE: Received final operation event for 56,12\n", $time);
            end
            begin
              @(final_operation[56][13]) ;
              //$display("@%0t LEE: Received final operation event for 56,13\n", $time);
            end
            begin
              @(final_operation[56][14]) ;
              //$display("@%0t LEE: Received final operation event for 56,14\n", $time);
            end
            begin
              @(final_operation[56][15]) ;
              //$display("@%0t LEE: Received final operation event for 56,15\n", $time);
            end
            begin
              @(final_operation[56][16]) ;
              //$display("@%0t LEE: Received final operation event for 56,16\n", $time);
            end
            begin
              @(final_operation[56][17]) ;
              //$display("@%0t LEE: Received final operation event for 56,17\n", $time);
            end
            begin
              @(final_operation[56][18]) ;
              //$display("@%0t LEE: Received final operation event for 56,18\n", $time);
            end
            begin
              @(final_operation[56][19]) ;
              //$display("@%0t LEE: Received final operation event for 56,19\n", $time);
            end
            begin
              @(final_operation[56][20]) ;
              //$display("@%0t LEE: Received final operation event for 56,20\n", $time);
            end
            begin
              @(final_operation[56][21]) ;
              //$display("@%0t LEE: Received final operation event for 56,21\n", $time);
            end
            begin
              @(final_operation[56][22]) ;
              //$display("@%0t LEE: Received final operation event for 56,22\n", $time);
            end
            begin
              @(final_operation[56][23]) ;
              //$display("@%0t LEE: Received final operation event for 56,23\n", $time);
            end
            begin
              @(final_operation[56][24]) ;
              //$display("@%0t LEE: Received final operation event for 56,24\n", $time);
            end
            begin
              @(final_operation[56][25]) ;
              //$display("@%0t LEE: Received final operation event for 56,25\n", $time);
            end
            begin
              @(final_operation[56][26]) ;
              //$display("@%0t LEE: Received final operation event for 56,26\n", $time);
            end
            begin
              @(final_operation[56][27]) ;
              //$display("@%0t LEE: Received final operation event for 56,27\n", $time);
            end
            begin
              @(final_operation[56][28]) ;
              //$display("@%0t LEE: Received final operation event for 56,28\n", $time);
            end
            begin
              @(final_operation[56][29]) ;
              //$display("@%0t LEE: Received final operation event for 56,29\n", $time);
            end
            begin
              @(final_operation[56][30]) ;
              //$display("@%0t LEE: Received final operation event for 56,30\n", $time);
            end
            begin
              @(final_operation[56][31]) ;
              //$display("@%0t LEE: Received final operation event for 56,31\n", $time);
            end

            begin
              @(final_operation[57][0]) ;
              //$display("@%0t LEE: Received final operation event for 57,0\n", $time);
            end
            begin
              @(final_operation[57][1]) ;
              //$display("@%0t LEE: Received final operation event for 57,1\n", $time);
            end
            begin
              @(final_operation[57][2]) ;
              //$display("@%0t LEE: Received final operation event for 57,2\n", $time);
            end
            begin
              @(final_operation[57][3]) ;
              //$display("@%0t LEE: Received final operation event for 57,3\n", $time);
            end
            begin
              @(final_operation[57][4]) ;
              //$display("@%0t LEE: Received final operation event for 57,4\n", $time);
            end
            begin
              @(final_operation[57][5]) ;
              //$display("@%0t LEE: Received final operation event for 57,5\n", $time);
            end
            begin
              @(final_operation[57][6]) ;
              //$display("@%0t LEE: Received final operation event for 57,6\n", $time);
            end
            begin
              @(final_operation[57][7]) ;
              //$display("@%0t LEE: Received final operation event for 57,7\n", $time);
            end
            begin
              @(final_operation[57][8]) ;
              //$display("@%0t LEE: Received final operation event for 57,8\n", $time);
            end
            begin
              @(final_operation[57][9]) ;
              //$display("@%0t LEE: Received final operation event for 57,9\n", $time);
            end
            begin
              @(final_operation[57][10]) ;
              //$display("@%0t LEE: Received final operation event for 57,10\n", $time);
            end
            begin
              @(final_operation[57][11]) ;
              //$display("@%0t LEE: Received final operation event for 57,11\n", $time);
            end
            begin
              @(final_operation[57][12]) ;
              //$display("@%0t LEE: Received final operation event for 57,12\n", $time);
            end
            begin
              @(final_operation[57][13]) ;
              //$display("@%0t LEE: Received final operation event for 57,13\n", $time);
            end
            begin
              @(final_operation[57][14]) ;
              //$display("@%0t LEE: Received final operation event for 57,14\n", $time);
            end
            begin
              @(final_operation[57][15]) ;
              //$display("@%0t LEE: Received final operation event for 57,15\n", $time);
            end
            begin
              @(final_operation[57][16]) ;
              //$display("@%0t LEE: Received final operation event for 57,16\n", $time);
            end
            begin
              @(final_operation[57][17]) ;
              //$display("@%0t LEE: Received final operation event for 57,17\n", $time);
            end
            begin
              @(final_operation[57][18]) ;
              //$display("@%0t LEE: Received final operation event for 57,18\n", $time);
            end
            begin
              @(final_operation[57][19]) ;
              //$display("@%0t LEE: Received final operation event for 57,19\n", $time);
            end
            begin
              @(final_operation[57][20]) ;
              //$display("@%0t LEE: Received final operation event for 57,20\n", $time);
            end
            begin
              @(final_operation[57][21]) ;
              //$display("@%0t LEE: Received final operation event for 57,21\n", $time);
            end
            begin
              @(final_operation[57][22]) ;
              //$display("@%0t LEE: Received final operation event for 57,22\n", $time);
            end
            begin
              @(final_operation[57][23]) ;
              //$display("@%0t LEE: Received final operation event for 57,23\n", $time);
            end
            begin
              @(final_operation[57][24]) ;
              //$display("@%0t LEE: Received final operation event for 57,24\n", $time);
            end
            begin
              @(final_operation[57][25]) ;
              //$display("@%0t LEE: Received final operation event for 57,25\n", $time);
            end
            begin
              @(final_operation[57][26]) ;
              //$display("@%0t LEE: Received final operation event for 57,26\n", $time);
            end
            begin
              @(final_operation[57][27]) ;
              //$display("@%0t LEE: Received final operation event for 57,27\n", $time);
            end
            begin
              @(final_operation[57][28]) ;
              //$display("@%0t LEE: Received final operation event for 57,28\n", $time);
            end
            begin
              @(final_operation[57][29]) ;
              //$display("@%0t LEE: Received final operation event for 57,29\n", $time);
            end
            begin
              @(final_operation[57][30]) ;
              //$display("@%0t LEE: Received final operation event for 57,30\n", $time);
            end
            begin
              @(final_operation[57][31]) ;
              //$display("@%0t LEE: Received final operation event for 57,31\n", $time);
            end

            begin
              @(final_operation[58][0]) ;
              //$display("@%0t LEE: Received final operation event for 58,0\n", $time);
            end
            begin
              @(final_operation[58][1]) ;
              //$display("@%0t LEE: Received final operation event for 58,1\n", $time);
            end
            begin
              @(final_operation[58][2]) ;
              //$display("@%0t LEE: Received final operation event for 58,2\n", $time);
            end
            begin
              @(final_operation[58][3]) ;
              //$display("@%0t LEE: Received final operation event for 58,3\n", $time);
            end
            begin
              @(final_operation[58][4]) ;
              //$display("@%0t LEE: Received final operation event for 58,4\n", $time);
            end
            begin
              @(final_operation[58][5]) ;
              //$display("@%0t LEE: Received final operation event for 58,5\n", $time);
            end
            begin
              @(final_operation[58][6]) ;
              //$display("@%0t LEE: Received final operation event for 58,6\n", $time);
            end
            begin
              @(final_operation[58][7]) ;
              //$display("@%0t LEE: Received final operation event for 58,7\n", $time);
            end
            begin
              @(final_operation[58][8]) ;
              //$display("@%0t LEE: Received final operation event for 58,8\n", $time);
            end
            begin
              @(final_operation[58][9]) ;
              //$display("@%0t LEE: Received final operation event for 58,9\n", $time);
            end
            begin
              @(final_operation[58][10]) ;
              //$display("@%0t LEE: Received final operation event for 58,10\n", $time);
            end
            begin
              @(final_operation[58][11]) ;
              //$display("@%0t LEE: Received final operation event for 58,11\n", $time);
            end
            begin
              @(final_operation[58][12]) ;
              //$display("@%0t LEE: Received final operation event for 58,12\n", $time);
            end
            begin
              @(final_operation[58][13]) ;
              //$display("@%0t LEE: Received final operation event for 58,13\n", $time);
            end
            begin
              @(final_operation[58][14]) ;
              //$display("@%0t LEE: Received final operation event for 58,14\n", $time);
            end
            begin
              @(final_operation[58][15]) ;
              //$display("@%0t LEE: Received final operation event for 58,15\n", $time);
            end
            begin
              @(final_operation[58][16]) ;
              //$display("@%0t LEE: Received final operation event for 58,16\n", $time);
            end
            begin
              @(final_operation[58][17]) ;
              //$display("@%0t LEE: Received final operation event for 58,17\n", $time);
            end
            begin
              @(final_operation[58][18]) ;
              //$display("@%0t LEE: Received final operation event for 58,18\n", $time);
            end
            begin
              @(final_operation[58][19]) ;
              //$display("@%0t LEE: Received final operation event for 58,19\n", $time);
            end
            begin
              @(final_operation[58][20]) ;
              //$display("@%0t LEE: Received final operation event for 58,20\n", $time);
            end
            begin
              @(final_operation[58][21]) ;
              //$display("@%0t LEE: Received final operation event for 58,21\n", $time);
            end
            begin
              @(final_operation[58][22]) ;
              //$display("@%0t LEE: Received final operation event for 58,22\n", $time);
            end
            begin
              @(final_operation[58][23]) ;
              //$display("@%0t LEE: Received final operation event for 58,23\n", $time);
            end
            begin
              @(final_operation[58][24]) ;
              //$display("@%0t LEE: Received final operation event for 58,24\n", $time);
            end
            begin
              @(final_operation[58][25]) ;
              //$display("@%0t LEE: Received final operation event for 58,25\n", $time);
            end
            begin
              @(final_operation[58][26]) ;
              //$display("@%0t LEE: Received final operation event for 58,26\n", $time);
            end
            begin
              @(final_operation[58][27]) ;
              //$display("@%0t LEE: Received final operation event for 58,27\n", $time);
            end
            begin
              @(final_operation[58][28]) ;
              //$display("@%0t LEE: Received final operation event for 58,28\n", $time);
            end
            begin
              @(final_operation[58][29]) ;
              //$display("@%0t LEE: Received final operation event for 58,29\n", $time);
            end
            begin
              @(final_operation[58][30]) ;
              //$display("@%0t LEE: Received final operation event for 58,30\n", $time);
            end
            begin
              @(final_operation[58][31]) ;
              //$display("@%0t LEE: Received final operation event for 58,31\n", $time);
            end

            begin
              @(final_operation[59][0]) ;
              //$display("@%0t LEE: Received final operation event for 59,0\n", $time);
            end
            begin
              @(final_operation[59][1]) ;
              //$display("@%0t LEE: Received final operation event for 59,1\n", $time);
            end
            begin
              @(final_operation[59][2]) ;
              //$display("@%0t LEE: Received final operation event for 59,2\n", $time);
            end
            begin
              @(final_operation[59][3]) ;
              //$display("@%0t LEE: Received final operation event for 59,3\n", $time);
            end
            begin
              @(final_operation[59][4]) ;
              //$display("@%0t LEE: Received final operation event for 59,4\n", $time);
            end
            begin
              @(final_operation[59][5]) ;
              //$display("@%0t LEE: Received final operation event for 59,5\n", $time);
            end
            begin
              @(final_operation[59][6]) ;
              //$display("@%0t LEE: Received final operation event for 59,6\n", $time);
            end
            begin
              @(final_operation[59][7]) ;
              //$display("@%0t LEE: Received final operation event for 59,7\n", $time);
            end
            begin
              @(final_operation[59][8]) ;
              //$display("@%0t LEE: Received final operation event for 59,8\n", $time);
            end
            begin
              @(final_operation[59][9]) ;
              //$display("@%0t LEE: Received final operation event for 59,9\n", $time);
            end
            begin
              @(final_operation[59][10]) ;
              //$display("@%0t LEE: Received final operation event for 59,10\n", $time);
            end
            begin
              @(final_operation[59][11]) ;
              //$display("@%0t LEE: Received final operation event for 59,11\n", $time);
            end
            begin
              @(final_operation[59][12]) ;
              //$display("@%0t LEE: Received final operation event for 59,12\n", $time);
            end
            begin
              @(final_operation[59][13]) ;
              //$display("@%0t LEE: Received final operation event for 59,13\n", $time);
            end
            begin
              @(final_operation[59][14]) ;
              //$display("@%0t LEE: Received final operation event for 59,14\n", $time);
            end
            begin
              @(final_operation[59][15]) ;
              //$display("@%0t LEE: Received final operation event for 59,15\n", $time);
            end
            begin
              @(final_operation[59][16]) ;
              //$display("@%0t LEE: Received final operation event for 59,16\n", $time);
            end
            begin
              @(final_operation[59][17]) ;
              //$display("@%0t LEE: Received final operation event for 59,17\n", $time);
            end
            begin
              @(final_operation[59][18]) ;
              //$display("@%0t LEE: Received final operation event for 59,18\n", $time);
            end
            begin
              @(final_operation[59][19]) ;
              //$display("@%0t LEE: Received final operation event for 59,19\n", $time);
            end
            begin
              @(final_operation[59][20]) ;
              //$display("@%0t LEE: Received final operation event for 59,20\n", $time);
            end
            begin
              @(final_operation[59][21]) ;
              //$display("@%0t LEE: Received final operation event for 59,21\n", $time);
            end
            begin
              @(final_operation[59][22]) ;
              //$display("@%0t LEE: Received final operation event for 59,22\n", $time);
            end
            begin
              @(final_operation[59][23]) ;
              //$display("@%0t LEE: Received final operation event for 59,23\n", $time);
            end
            begin
              @(final_operation[59][24]) ;
              //$display("@%0t LEE: Received final operation event for 59,24\n", $time);
            end
            begin
              @(final_operation[59][25]) ;
              //$display("@%0t LEE: Received final operation event for 59,25\n", $time);
            end
            begin
              @(final_operation[59][26]) ;
              //$display("@%0t LEE: Received final operation event for 59,26\n", $time);
            end
            begin
              @(final_operation[59][27]) ;
              //$display("@%0t LEE: Received final operation event for 59,27\n", $time);
            end
            begin
              @(final_operation[59][28]) ;
              //$display("@%0t LEE: Received final operation event for 59,28\n", $time);
            end
            begin
              @(final_operation[59][29]) ;
              //$display("@%0t LEE: Received final operation event for 59,29\n", $time);
            end
            begin
              @(final_operation[59][30]) ;
              //$display("@%0t LEE: Received final operation event for 59,30\n", $time);
            end
            begin
              @(final_operation[59][31]) ;
              //$display("@%0t LEE: Received final operation event for 59,31\n", $time);
            end

            begin
              @(final_operation[60][0]) ;
              //$display("@%0t LEE: Received final operation event for 60,0\n", $time);
            end
            begin
              @(final_operation[60][1]) ;
              //$display("@%0t LEE: Received final operation event for 60,1\n", $time);
            end
            begin
              @(final_operation[60][2]) ;
              //$display("@%0t LEE: Received final operation event for 60,2\n", $time);
            end
            begin
              @(final_operation[60][3]) ;
              //$display("@%0t LEE: Received final operation event for 60,3\n", $time);
            end
            begin
              @(final_operation[60][4]) ;
              //$display("@%0t LEE: Received final operation event for 60,4\n", $time);
            end
            begin
              @(final_operation[60][5]) ;
              //$display("@%0t LEE: Received final operation event for 60,5\n", $time);
            end
            begin
              @(final_operation[60][6]) ;
              //$display("@%0t LEE: Received final operation event for 60,6\n", $time);
            end
            begin
              @(final_operation[60][7]) ;
              //$display("@%0t LEE: Received final operation event for 60,7\n", $time);
            end
            begin
              @(final_operation[60][8]) ;
              //$display("@%0t LEE: Received final operation event for 60,8\n", $time);
            end
            begin
              @(final_operation[60][9]) ;
              //$display("@%0t LEE: Received final operation event for 60,9\n", $time);
            end
            begin
              @(final_operation[60][10]) ;
              //$display("@%0t LEE: Received final operation event for 60,10\n", $time);
            end
            begin
              @(final_operation[60][11]) ;
              //$display("@%0t LEE: Received final operation event for 60,11\n", $time);
            end
            begin
              @(final_operation[60][12]) ;
              //$display("@%0t LEE: Received final operation event for 60,12\n", $time);
            end
            begin
              @(final_operation[60][13]) ;
              //$display("@%0t LEE: Received final operation event for 60,13\n", $time);
            end
            begin
              @(final_operation[60][14]) ;
              //$display("@%0t LEE: Received final operation event for 60,14\n", $time);
            end
            begin
              @(final_operation[60][15]) ;
              //$display("@%0t LEE: Received final operation event for 60,15\n", $time);
            end
            begin
              @(final_operation[60][16]) ;
              //$display("@%0t LEE: Received final operation event for 60,16\n", $time);
            end
            begin
              @(final_operation[60][17]) ;
              //$display("@%0t LEE: Received final operation event for 60,17\n", $time);
            end
            begin
              @(final_operation[60][18]) ;
              //$display("@%0t LEE: Received final operation event for 60,18\n", $time);
            end
            begin
              @(final_operation[60][19]) ;
              //$display("@%0t LEE: Received final operation event for 60,19\n", $time);
            end
            begin
              @(final_operation[60][20]) ;
              //$display("@%0t LEE: Received final operation event for 60,20\n", $time);
            end
            begin
              @(final_operation[60][21]) ;
              //$display("@%0t LEE: Received final operation event for 60,21\n", $time);
            end
            begin
              @(final_operation[60][22]) ;
              //$display("@%0t LEE: Received final operation event for 60,22\n", $time);
            end
            begin
              @(final_operation[60][23]) ;
              //$display("@%0t LEE: Received final operation event for 60,23\n", $time);
            end
            begin
              @(final_operation[60][24]) ;
              //$display("@%0t LEE: Received final operation event for 60,24\n", $time);
            end
            begin
              @(final_operation[60][25]) ;
              //$display("@%0t LEE: Received final operation event for 60,25\n", $time);
            end
            begin
              @(final_operation[60][26]) ;
              //$display("@%0t LEE: Received final operation event for 60,26\n", $time);
            end
            begin
              @(final_operation[60][27]) ;
              //$display("@%0t LEE: Received final operation event for 60,27\n", $time);
            end
            begin
              @(final_operation[60][28]) ;
              //$display("@%0t LEE: Received final operation event for 60,28\n", $time);
            end
            begin
              @(final_operation[60][29]) ;
              //$display("@%0t LEE: Received final operation event for 60,29\n", $time);
            end
            begin
              @(final_operation[60][30]) ;
              //$display("@%0t LEE: Received final operation event for 60,30\n", $time);
            end
            begin
              @(final_operation[60][31]) ;
              //$display("@%0t LEE: Received final operation event for 60,31\n", $time);
            end

            begin
              @(final_operation[61][0]) ;
              //$display("@%0t LEE: Received final operation event for 61,0\n", $time);
            end
            begin
              @(final_operation[61][1]) ;
              //$display("@%0t LEE: Received final operation event for 61,1\n", $time);
            end
            begin
              @(final_operation[61][2]) ;
              //$display("@%0t LEE: Received final operation event for 61,2\n", $time);
            end
            begin
              @(final_operation[61][3]) ;
              //$display("@%0t LEE: Received final operation event for 61,3\n", $time);
            end
            begin
              @(final_operation[61][4]) ;
              //$display("@%0t LEE: Received final operation event for 61,4\n", $time);
            end
            begin
              @(final_operation[61][5]) ;
              //$display("@%0t LEE: Received final operation event for 61,5\n", $time);
            end
            begin
              @(final_operation[61][6]) ;
              //$display("@%0t LEE: Received final operation event for 61,6\n", $time);
            end
            begin
              @(final_operation[61][7]) ;
              //$display("@%0t LEE: Received final operation event for 61,7\n", $time);
            end
            begin
              @(final_operation[61][8]) ;
              //$display("@%0t LEE: Received final operation event for 61,8\n", $time);
            end
            begin
              @(final_operation[61][9]) ;
              //$display("@%0t LEE: Received final operation event for 61,9\n", $time);
            end
            begin
              @(final_operation[61][10]) ;
              //$display("@%0t LEE: Received final operation event for 61,10\n", $time);
            end
            begin
              @(final_operation[61][11]) ;
              //$display("@%0t LEE: Received final operation event for 61,11\n", $time);
            end
            begin
              @(final_operation[61][12]) ;
              //$display("@%0t LEE: Received final operation event for 61,12\n", $time);
            end
            begin
              @(final_operation[61][13]) ;
              //$display("@%0t LEE: Received final operation event for 61,13\n", $time);
            end
            begin
              @(final_operation[61][14]) ;
              //$display("@%0t LEE: Received final operation event for 61,14\n", $time);
            end
            begin
              @(final_operation[61][15]) ;
              //$display("@%0t LEE: Received final operation event for 61,15\n", $time);
            end
            begin
              @(final_operation[61][16]) ;
              //$display("@%0t LEE: Received final operation event for 61,16\n", $time);
            end
            begin
              @(final_operation[61][17]) ;
              //$display("@%0t LEE: Received final operation event for 61,17\n", $time);
            end
            begin
              @(final_operation[61][18]) ;
              //$display("@%0t LEE: Received final operation event for 61,18\n", $time);
            end
            begin
              @(final_operation[61][19]) ;
              //$display("@%0t LEE: Received final operation event for 61,19\n", $time);
            end
            begin
              @(final_operation[61][20]) ;
              //$display("@%0t LEE: Received final operation event for 61,20\n", $time);
            end
            begin
              @(final_operation[61][21]) ;
              //$display("@%0t LEE: Received final operation event for 61,21\n", $time);
            end
            begin
              @(final_operation[61][22]) ;
              //$display("@%0t LEE: Received final operation event for 61,22\n", $time);
            end
            begin
              @(final_operation[61][23]) ;
              //$display("@%0t LEE: Received final operation event for 61,23\n", $time);
            end
            begin
              @(final_operation[61][24]) ;
              //$display("@%0t LEE: Received final operation event for 61,24\n", $time);
            end
            begin
              @(final_operation[61][25]) ;
              //$display("@%0t LEE: Received final operation event for 61,25\n", $time);
            end
            begin
              @(final_operation[61][26]) ;
              //$display("@%0t LEE: Received final operation event for 61,26\n", $time);
            end
            begin
              @(final_operation[61][27]) ;
              //$display("@%0t LEE: Received final operation event for 61,27\n", $time);
            end
            begin
              @(final_operation[61][28]) ;
              //$display("@%0t LEE: Received final operation event for 61,28\n", $time);
            end
            begin
              @(final_operation[61][29]) ;
              //$display("@%0t LEE: Received final operation event for 61,29\n", $time);
            end
            begin
              @(final_operation[61][30]) ;
              //$display("@%0t LEE: Received final operation event for 61,30\n", $time);
            end
            begin
              @(final_operation[61][31]) ;
              //$display("@%0t LEE: Received final operation event for 61,31\n", $time);
            end

            begin
              @(final_operation[62][0]) ;
              //$display("@%0t LEE: Received final operation event for 62,0\n", $time);
            end
            begin
              @(final_operation[62][1]) ;
              //$display("@%0t LEE: Received final operation event for 62,1\n", $time);
            end
            begin
              @(final_operation[62][2]) ;
              //$display("@%0t LEE: Received final operation event for 62,2\n", $time);
            end
            begin
              @(final_operation[62][3]) ;
              //$display("@%0t LEE: Received final operation event for 62,3\n", $time);
            end
            begin
              @(final_operation[62][4]) ;
              //$display("@%0t LEE: Received final operation event for 62,4\n", $time);
            end
            begin
              @(final_operation[62][5]) ;
              //$display("@%0t LEE: Received final operation event for 62,5\n", $time);
            end
            begin
              @(final_operation[62][6]) ;
              //$display("@%0t LEE: Received final operation event for 62,6\n", $time);
            end
            begin
              @(final_operation[62][7]) ;
              //$display("@%0t LEE: Received final operation event for 62,7\n", $time);
            end
            begin
              @(final_operation[62][8]) ;
              //$display("@%0t LEE: Received final operation event for 62,8\n", $time);
            end
            begin
              @(final_operation[62][9]) ;
              //$display("@%0t LEE: Received final operation event for 62,9\n", $time);
            end
            begin
              @(final_operation[62][10]) ;
              //$display("@%0t LEE: Received final operation event for 62,10\n", $time);
            end
            begin
              @(final_operation[62][11]) ;
              //$display("@%0t LEE: Received final operation event for 62,11\n", $time);
            end
            begin
              @(final_operation[62][12]) ;
              //$display("@%0t LEE: Received final operation event for 62,12\n", $time);
            end
            begin
              @(final_operation[62][13]) ;
              //$display("@%0t LEE: Received final operation event for 62,13\n", $time);
            end
            begin
              @(final_operation[62][14]) ;
              //$display("@%0t LEE: Received final operation event for 62,14\n", $time);
            end
            begin
              @(final_operation[62][15]) ;
              //$display("@%0t LEE: Received final operation event for 62,15\n", $time);
            end
            begin
              @(final_operation[62][16]) ;
              //$display("@%0t LEE: Received final operation event for 62,16\n", $time);
            end
            begin
              @(final_operation[62][17]) ;
              //$display("@%0t LEE: Received final operation event for 62,17\n", $time);
            end
            begin
              @(final_operation[62][18]) ;
              //$display("@%0t LEE: Received final operation event for 62,18\n", $time);
            end
            begin
              @(final_operation[62][19]) ;
              //$display("@%0t LEE: Received final operation event for 62,19\n", $time);
            end
            begin
              @(final_operation[62][20]) ;
              //$display("@%0t LEE: Received final operation event for 62,20\n", $time);
            end
            begin
              @(final_operation[62][21]) ;
              //$display("@%0t LEE: Received final operation event for 62,21\n", $time);
            end
            begin
              @(final_operation[62][22]) ;
              //$display("@%0t LEE: Received final operation event for 62,22\n", $time);
            end
            begin
              @(final_operation[62][23]) ;
              //$display("@%0t LEE: Received final operation event for 62,23\n", $time);
            end
            begin
              @(final_operation[62][24]) ;
              //$display("@%0t LEE: Received final operation event for 62,24\n", $time);
            end
            begin
              @(final_operation[62][25]) ;
              //$display("@%0t LEE: Received final operation event for 62,25\n", $time);
            end
            begin
              @(final_operation[62][26]) ;
              //$display("@%0t LEE: Received final operation event for 62,26\n", $time);
            end
            begin
              @(final_operation[62][27]) ;
              //$display("@%0t LEE: Received final operation event for 62,27\n", $time);
            end
            begin
              @(final_operation[62][28]) ;
              //$display("@%0t LEE: Received final operation event for 62,28\n", $time);
            end
            begin
              @(final_operation[62][29]) ;
              //$display("@%0t LEE: Received final operation event for 62,29\n", $time);
            end
            begin
              @(final_operation[62][30]) ;
              //$display("@%0t LEE: Received final operation event for 62,30\n", $time);
            end
            begin
              @(final_operation[62][31]) ;
              //$display("@%0t LEE: Received final operation event for 62,31\n", $time);
            end

            begin
              @(final_operation[63][0]) ;
              //$display("@%0t LEE: Received final operation event for 63,0\n", $time);
            end
            begin
              @(final_operation[63][1]) ;
              //$display("@%0t LEE: Received final operation event for 63,1\n", $time);
            end
            begin
              @(final_operation[63][2]) ;
              //$display("@%0t LEE: Received final operation event for 63,2\n", $time);
            end
            begin
              @(final_operation[63][3]) ;
              //$display("@%0t LEE: Received final operation event for 63,3\n", $time);
            end
            begin
              @(final_operation[63][4]) ;
              //$display("@%0t LEE: Received final operation event for 63,4\n", $time);
            end
            begin
              @(final_operation[63][5]) ;
              //$display("@%0t LEE: Received final operation event for 63,5\n", $time);
            end
            begin
              @(final_operation[63][6]) ;
              //$display("@%0t LEE: Received final operation event for 63,6\n", $time);
            end
            begin
              @(final_operation[63][7]) ;
              //$display("@%0t LEE: Received final operation event for 63,7\n", $time);
            end
            begin
              @(final_operation[63][8]) ;
              //$display("@%0t LEE: Received final operation event for 63,8\n", $time);
            end
            begin
              @(final_operation[63][9]) ;
              //$display("@%0t LEE: Received final operation event for 63,9\n", $time);
            end
            begin
              @(final_operation[63][10]) ;
              //$display("@%0t LEE: Received final operation event for 63,10\n", $time);
            end
            begin
              @(final_operation[63][11]) ;
              //$display("@%0t LEE: Received final operation event for 63,11\n", $time);
            end
            begin
              @(final_operation[63][12]) ;
              //$display("@%0t LEE: Received final operation event for 63,12\n", $time);
            end
            begin
              @(final_operation[63][13]) ;
              //$display("@%0t LEE: Received final operation event for 63,13\n", $time);
            end
            begin
              @(final_operation[63][14]) ;
              //$display("@%0t LEE: Received final operation event for 63,14\n", $time);
            end
            begin
              @(final_operation[63][15]) ;
              //$display("@%0t LEE: Received final operation event for 63,15\n", $time);
            end
            begin
              @(final_operation[63][16]) ;
              //$display("@%0t LEE: Received final operation event for 63,16\n", $time);
            end
            begin
              @(final_operation[63][17]) ;
              //$display("@%0t LEE: Received final operation event for 63,17\n", $time);
            end
            begin
              @(final_operation[63][18]) ;
              //$display("@%0t LEE: Received final operation event for 63,18\n", $time);
            end
            begin
              @(final_operation[63][19]) ;
              //$display("@%0t LEE: Received final operation event for 63,19\n", $time);
            end
            begin
              @(final_operation[63][20]) ;
              //$display("@%0t LEE: Received final operation event for 63,20\n", $time);
            end
            begin
              @(final_operation[63][21]) ;
              //$display("@%0t LEE: Received final operation event for 63,21\n", $time);
            end
            begin
              @(final_operation[63][22]) ;
              //$display("@%0t LEE: Received final operation event for 63,22\n", $time);
            end
            begin
              @(final_operation[63][23]) ;
              //$display("@%0t LEE: Received final operation event for 63,23\n", $time);
            end
            begin
              @(final_operation[63][24]) ;
              //$display("@%0t LEE: Received final operation event for 63,24\n", $time);
            end
            begin
              @(final_operation[63][25]) ;
              //$display("@%0t LEE: Received final operation event for 63,25\n", $time);
            end
            begin
              @(final_operation[63][26]) ;
              //$display("@%0t LEE: Received final operation event for 63,26\n", $time);
            end
            begin
              @(final_operation[63][27]) ;
              //$display("@%0t LEE: Received final operation event for 63,27\n", $time);
            end
            begin
              @(final_operation[63][28]) ;
              //$display("@%0t LEE: Received final operation event for 63,28\n", $time);
            end
            begin
              @(final_operation[63][29]) ;
              //$display("@%0t LEE: Received final operation event for 63,29\n", $time);
            end
            begin
              @(final_operation[63][30]) ;
              //$display("@%0t LEE: Received final operation event for 63,30\n", $time);
            end
            begin
              @(final_operation[63][31]) ;
              //$display("@%0t LEE: Received final operation event for 63,31\n", $time);
            end
