package virtual_interface;
`timescale 1ns/10ps
    typedef virtual std_pe_lane_ifc.vSys2PeArray_T  vSys2PeArray_T ;
    typedef virtual pe_dma2mem_ifc.vDma2Mem_T       vDma2Mem_T     ;
    // FIXME : add more see MC 
endpackage:virtual_interface
    
