
            begin
                @vSys2PeArray[0][0].cb_test                                      ;
                vSys2PeArray [0][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][1].cb_test                                      ;
                vSys2PeArray [0][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][2].cb_test                                      ;
                vSys2PeArray [0][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][3].cb_test                                      ;
                vSys2PeArray [0][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][4].cb_test                                      ;
                vSys2PeArray [0][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][5].cb_test                                      ;
                vSys2PeArray [0][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][6].cb_test                                      ;
                vSys2PeArray [0][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][7].cb_test                                      ;
                vSys2PeArray [0][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][8].cb_test                                      ;
                vSys2PeArray [0][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][9].cb_test                                      ;
                vSys2PeArray [0][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][10].cb_test                                      ;
                vSys2PeArray [0][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][11].cb_test                                      ;
                vSys2PeArray [0][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][12].cb_test                                      ;
                vSys2PeArray [0][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][13].cb_test                                      ;
                vSys2PeArray [0][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][14].cb_test                                      ;
                vSys2PeArray [0][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][15].cb_test                                      ;
                vSys2PeArray [0][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][16].cb_test                                      ;
                vSys2PeArray [0][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][17].cb_test                                      ;
                vSys2PeArray [0][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][18].cb_test                                      ;
                vSys2PeArray [0][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][19].cb_test                                      ;
                vSys2PeArray [0][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][20].cb_test                                      ;
                vSys2PeArray [0][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][21].cb_test                                      ;
                vSys2PeArray [0][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][22].cb_test                                      ;
                vSys2PeArray [0][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][23].cb_test                                      ;
                vSys2PeArray [0][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][24].cb_test                                      ;
                vSys2PeArray [0][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][25].cb_test                                      ;
                vSys2PeArray [0][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][26].cb_test                                      ;
                vSys2PeArray [0][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][27].cb_test                                      ;
                vSys2PeArray [0][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][28].cb_test                                      ;
                vSys2PeArray [0][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][29].cb_test                                      ;
                vSys2PeArray [0][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][30].cb_test                                      ;
                vSys2PeArray [0][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[0][31].cb_test                                      ;
                vSys2PeArray [0][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [0][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[1][0].cb_test                                      ;
                vSys2PeArray [1][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][1].cb_test                                      ;
                vSys2PeArray [1][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][2].cb_test                                      ;
                vSys2PeArray [1][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][3].cb_test                                      ;
                vSys2PeArray [1][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][4].cb_test                                      ;
                vSys2PeArray [1][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][5].cb_test                                      ;
                vSys2PeArray [1][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][6].cb_test                                      ;
                vSys2PeArray [1][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][7].cb_test                                      ;
                vSys2PeArray [1][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][8].cb_test                                      ;
                vSys2PeArray [1][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][9].cb_test                                      ;
                vSys2PeArray [1][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][10].cb_test                                      ;
                vSys2PeArray [1][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][11].cb_test                                      ;
                vSys2PeArray [1][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][12].cb_test                                      ;
                vSys2PeArray [1][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][13].cb_test                                      ;
                vSys2PeArray [1][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][14].cb_test                                      ;
                vSys2PeArray [1][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][15].cb_test                                      ;
                vSys2PeArray [1][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][16].cb_test                                      ;
                vSys2PeArray [1][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][17].cb_test                                      ;
                vSys2PeArray [1][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][18].cb_test                                      ;
                vSys2PeArray [1][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][19].cb_test                                      ;
                vSys2PeArray [1][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][20].cb_test                                      ;
                vSys2PeArray [1][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][21].cb_test                                      ;
                vSys2PeArray [1][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][22].cb_test                                      ;
                vSys2PeArray [1][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][23].cb_test                                      ;
                vSys2PeArray [1][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][24].cb_test                                      ;
                vSys2PeArray [1][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][25].cb_test                                      ;
                vSys2PeArray [1][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][26].cb_test                                      ;
                vSys2PeArray [1][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][27].cb_test                                      ;
                vSys2PeArray [1][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][28].cb_test                                      ;
                vSys2PeArray [1][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][29].cb_test                                      ;
                vSys2PeArray [1][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][30].cb_test                                      ;
                vSys2PeArray [1][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[1][31].cb_test                                      ;
                vSys2PeArray [1][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [1][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[2][0].cb_test                                      ;
                vSys2PeArray [2][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][1].cb_test                                      ;
                vSys2PeArray [2][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][2].cb_test                                      ;
                vSys2PeArray [2][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][3].cb_test                                      ;
                vSys2PeArray [2][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][4].cb_test                                      ;
                vSys2PeArray [2][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][5].cb_test                                      ;
                vSys2PeArray [2][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][6].cb_test                                      ;
                vSys2PeArray [2][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][7].cb_test                                      ;
                vSys2PeArray [2][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][8].cb_test                                      ;
                vSys2PeArray [2][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][9].cb_test                                      ;
                vSys2PeArray [2][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][10].cb_test                                      ;
                vSys2PeArray [2][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][11].cb_test                                      ;
                vSys2PeArray [2][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][12].cb_test                                      ;
                vSys2PeArray [2][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][13].cb_test                                      ;
                vSys2PeArray [2][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][14].cb_test                                      ;
                vSys2PeArray [2][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][15].cb_test                                      ;
                vSys2PeArray [2][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][16].cb_test                                      ;
                vSys2PeArray [2][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][17].cb_test                                      ;
                vSys2PeArray [2][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][18].cb_test                                      ;
                vSys2PeArray [2][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][19].cb_test                                      ;
                vSys2PeArray [2][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][20].cb_test                                      ;
                vSys2PeArray [2][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][21].cb_test                                      ;
                vSys2PeArray [2][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][22].cb_test                                      ;
                vSys2PeArray [2][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][23].cb_test                                      ;
                vSys2PeArray [2][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][24].cb_test                                      ;
                vSys2PeArray [2][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][25].cb_test                                      ;
                vSys2PeArray [2][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][26].cb_test                                      ;
                vSys2PeArray [2][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][27].cb_test                                      ;
                vSys2PeArray [2][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][28].cb_test                                      ;
                vSys2PeArray [2][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][29].cb_test                                      ;
                vSys2PeArray [2][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][30].cb_test                                      ;
                vSys2PeArray [2][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[2][31].cb_test                                      ;
                vSys2PeArray [2][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [2][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[3][0].cb_test                                      ;
                vSys2PeArray [3][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][1].cb_test                                      ;
                vSys2PeArray [3][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][2].cb_test                                      ;
                vSys2PeArray [3][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][3].cb_test                                      ;
                vSys2PeArray [3][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][4].cb_test                                      ;
                vSys2PeArray [3][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][5].cb_test                                      ;
                vSys2PeArray [3][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][6].cb_test                                      ;
                vSys2PeArray [3][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][7].cb_test                                      ;
                vSys2PeArray [3][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][8].cb_test                                      ;
                vSys2PeArray [3][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][9].cb_test                                      ;
                vSys2PeArray [3][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][10].cb_test                                      ;
                vSys2PeArray [3][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][11].cb_test                                      ;
                vSys2PeArray [3][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][12].cb_test                                      ;
                vSys2PeArray [3][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][13].cb_test                                      ;
                vSys2PeArray [3][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][14].cb_test                                      ;
                vSys2PeArray [3][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][15].cb_test                                      ;
                vSys2PeArray [3][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][16].cb_test                                      ;
                vSys2PeArray [3][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][17].cb_test                                      ;
                vSys2PeArray [3][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][18].cb_test                                      ;
                vSys2PeArray [3][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][19].cb_test                                      ;
                vSys2PeArray [3][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][20].cb_test                                      ;
                vSys2PeArray [3][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][21].cb_test                                      ;
                vSys2PeArray [3][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][22].cb_test                                      ;
                vSys2PeArray [3][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][23].cb_test                                      ;
                vSys2PeArray [3][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][24].cb_test                                      ;
                vSys2PeArray [3][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][25].cb_test                                      ;
                vSys2PeArray [3][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][26].cb_test                                      ;
                vSys2PeArray [3][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][27].cb_test                                      ;
                vSys2PeArray [3][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][28].cb_test                                      ;
                vSys2PeArray [3][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][29].cb_test                                      ;
                vSys2PeArray [3][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][30].cb_test                                      ;
                vSys2PeArray [3][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[3][31].cb_test                                      ;
                vSys2PeArray [3][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [3][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[4][0].cb_test                                      ;
                vSys2PeArray [4][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][1].cb_test                                      ;
                vSys2PeArray [4][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][2].cb_test                                      ;
                vSys2PeArray [4][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][3].cb_test                                      ;
                vSys2PeArray [4][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][4].cb_test                                      ;
                vSys2PeArray [4][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][5].cb_test                                      ;
                vSys2PeArray [4][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][6].cb_test                                      ;
                vSys2PeArray [4][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][7].cb_test                                      ;
                vSys2PeArray [4][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][8].cb_test                                      ;
                vSys2PeArray [4][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][9].cb_test                                      ;
                vSys2PeArray [4][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][10].cb_test                                      ;
                vSys2PeArray [4][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][11].cb_test                                      ;
                vSys2PeArray [4][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][12].cb_test                                      ;
                vSys2PeArray [4][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][13].cb_test                                      ;
                vSys2PeArray [4][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][14].cb_test                                      ;
                vSys2PeArray [4][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][15].cb_test                                      ;
                vSys2PeArray [4][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][16].cb_test                                      ;
                vSys2PeArray [4][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][17].cb_test                                      ;
                vSys2PeArray [4][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][18].cb_test                                      ;
                vSys2PeArray [4][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][19].cb_test                                      ;
                vSys2PeArray [4][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][20].cb_test                                      ;
                vSys2PeArray [4][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][21].cb_test                                      ;
                vSys2PeArray [4][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][22].cb_test                                      ;
                vSys2PeArray [4][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][23].cb_test                                      ;
                vSys2PeArray [4][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][24].cb_test                                      ;
                vSys2PeArray [4][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][25].cb_test                                      ;
                vSys2PeArray [4][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][26].cb_test                                      ;
                vSys2PeArray [4][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][27].cb_test                                      ;
                vSys2PeArray [4][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][28].cb_test                                      ;
                vSys2PeArray [4][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][29].cb_test                                      ;
                vSys2PeArray [4][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][30].cb_test                                      ;
                vSys2PeArray [4][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[4][31].cb_test                                      ;
                vSys2PeArray [4][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [4][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[5][0].cb_test                                      ;
                vSys2PeArray [5][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][1].cb_test                                      ;
                vSys2PeArray [5][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][2].cb_test                                      ;
                vSys2PeArray [5][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][3].cb_test                                      ;
                vSys2PeArray [5][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][4].cb_test                                      ;
                vSys2PeArray [5][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][5].cb_test                                      ;
                vSys2PeArray [5][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][6].cb_test                                      ;
                vSys2PeArray [5][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][7].cb_test                                      ;
                vSys2PeArray [5][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][8].cb_test                                      ;
                vSys2PeArray [5][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][9].cb_test                                      ;
                vSys2PeArray [5][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][10].cb_test                                      ;
                vSys2PeArray [5][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][11].cb_test                                      ;
                vSys2PeArray [5][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][12].cb_test                                      ;
                vSys2PeArray [5][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][13].cb_test                                      ;
                vSys2PeArray [5][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][14].cb_test                                      ;
                vSys2PeArray [5][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][15].cb_test                                      ;
                vSys2PeArray [5][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][16].cb_test                                      ;
                vSys2PeArray [5][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][17].cb_test                                      ;
                vSys2PeArray [5][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][18].cb_test                                      ;
                vSys2PeArray [5][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][19].cb_test                                      ;
                vSys2PeArray [5][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][20].cb_test                                      ;
                vSys2PeArray [5][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][21].cb_test                                      ;
                vSys2PeArray [5][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][22].cb_test                                      ;
                vSys2PeArray [5][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][23].cb_test                                      ;
                vSys2PeArray [5][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][24].cb_test                                      ;
                vSys2PeArray [5][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][25].cb_test                                      ;
                vSys2PeArray [5][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][26].cb_test                                      ;
                vSys2PeArray [5][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][27].cb_test                                      ;
                vSys2PeArray [5][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][28].cb_test                                      ;
                vSys2PeArray [5][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][29].cb_test                                      ;
                vSys2PeArray [5][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][30].cb_test                                      ;
                vSys2PeArray [5][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[5][31].cb_test                                      ;
                vSys2PeArray [5][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [5][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[6][0].cb_test                                      ;
                vSys2PeArray [6][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][1].cb_test                                      ;
                vSys2PeArray [6][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][2].cb_test                                      ;
                vSys2PeArray [6][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][3].cb_test                                      ;
                vSys2PeArray [6][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][4].cb_test                                      ;
                vSys2PeArray [6][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][5].cb_test                                      ;
                vSys2PeArray [6][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][6].cb_test                                      ;
                vSys2PeArray [6][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][7].cb_test                                      ;
                vSys2PeArray [6][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][8].cb_test                                      ;
                vSys2PeArray [6][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][9].cb_test                                      ;
                vSys2PeArray [6][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][10].cb_test                                      ;
                vSys2PeArray [6][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][11].cb_test                                      ;
                vSys2PeArray [6][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][12].cb_test                                      ;
                vSys2PeArray [6][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][13].cb_test                                      ;
                vSys2PeArray [6][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][14].cb_test                                      ;
                vSys2PeArray [6][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][15].cb_test                                      ;
                vSys2PeArray [6][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][16].cb_test                                      ;
                vSys2PeArray [6][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][17].cb_test                                      ;
                vSys2PeArray [6][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][18].cb_test                                      ;
                vSys2PeArray [6][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][19].cb_test                                      ;
                vSys2PeArray [6][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][20].cb_test                                      ;
                vSys2PeArray [6][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][21].cb_test                                      ;
                vSys2PeArray [6][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][22].cb_test                                      ;
                vSys2PeArray [6][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][23].cb_test                                      ;
                vSys2PeArray [6][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][24].cb_test                                      ;
                vSys2PeArray [6][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][25].cb_test                                      ;
                vSys2PeArray [6][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][26].cb_test                                      ;
                vSys2PeArray [6][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][27].cb_test                                      ;
                vSys2PeArray [6][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][28].cb_test                                      ;
                vSys2PeArray [6][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][29].cb_test                                      ;
                vSys2PeArray [6][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][30].cb_test                                      ;
                vSys2PeArray [6][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[6][31].cb_test                                      ;
                vSys2PeArray [6][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [6][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[7][0].cb_test                                      ;
                vSys2PeArray [7][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][1].cb_test                                      ;
                vSys2PeArray [7][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][2].cb_test                                      ;
                vSys2PeArray [7][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][3].cb_test                                      ;
                vSys2PeArray [7][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][4].cb_test                                      ;
                vSys2PeArray [7][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][5].cb_test                                      ;
                vSys2PeArray [7][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][6].cb_test                                      ;
                vSys2PeArray [7][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][7].cb_test                                      ;
                vSys2PeArray [7][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][8].cb_test                                      ;
                vSys2PeArray [7][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][9].cb_test                                      ;
                vSys2PeArray [7][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][10].cb_test                                      ;
                vSys2PeArray [7][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][11].cb_test                                      ;
                vSys2PeArray [7][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][12].cb_test                                      ;
                vSys2PeArray [7][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][13].cb_test                                      ;
                vSys2PeArray [7][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][14].cb_test                                      ;
                vSys2PeArray [7][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][15].cb_test                                      ;
                vSys2PeArray [7][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][16].cb_test                                      ;
                vSys2PeArray [7][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][17].cb_test                                      ;
                vSys2PeArray [7][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][18].cb_test                                      ;
                vSys2PeArray [7][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][19].cb_test                                      ;
                vSys2PeArray [7][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][20].cb_test                                      ;
                vSys2PeArray [7][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][21].cb_test                                      ;
                vSys2PeArray [7][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][22].cb_test                                      ;
                vSys2PeArray [7][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][23].cb_test                                      ;
                vSys2PeArray [7][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][24].cb_test                                      ;
                vSys2PeArray [7][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][25].cb_test                                      ;
                vSys2PeArray [7][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][26].cb_test                                      ;
                vSys2PeArray [7][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][27].cb_test                                      ;
                vSys2PeArray [7][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][28].cb_test                                      ;
                vSys2PeArray [7][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][29].cb_test                                      ;
                vSys2PeArray [7][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][30].cb_test                                      ;
                vSys2PeArray [7][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[7][31].cb_test                                      ;
                vSys2PeArray [7][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [7][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[8][0].cb_test                                      ;
                vSys2PeArray [8][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][1].cb_test                                      ;
                vSys2PeArray [8][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][2].cb_test                                      ;
                vSys2PeArray [8][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][3].cb_test                                      ;
                vSys2PeArray [8][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][4].cb_test                                      ;
                vSys2PeArray [8][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][5].cb_test                                      ;
                vSys2PeArray [8][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][6].cb_test                                      ;
                vSys2PeArray [8][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][7].cb_test                                      ;
                vSys2PeArray [8][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][8].cb_test                                      ;
                vSys2PeArray [8][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][9].cb_test                                      ;
                vSys2PeArray [8][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][10].cb_test                                      ;
                vSys2PeArray [8][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][11].cb_test                                      ;
                vSys2PeArray [8][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][12].cb_test                                      ;
                vSys2PeArray [8][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][13].cb_test                                      ;
                vSys2PeArray [8][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][14].cb_test                                      ;
                vSys2PeArray [8][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][15].cb_test                                      ;
                vSys2PeArray [8][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][16].cb_test                                      ;
                vSys2PeArray [8][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][17].cb_test                                      ;
                vSys2PeArray [8][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][18].cb_test                                      ;
                vSys2PeArray [8][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][19].cb_test                                      ;
                vSys2PeArray [8][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][20].cb_test                                      ;
                vSys2PeArray [8][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][21].cb_test                                      ;
                vSys2PeArray [8][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][22].cb_test                                      ;
                vSys2PeArray [8][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][23].cb_test                                      ;
                vSys2PeArray [8][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][24].cb_test                                      ;
                vSys2PeArray [8][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][25].cb_test                                      ;
                vSys2PeArray [8][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][26].cb_test                                      ;
                vSys2PeArray [8][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][27].cb_test                                      ;
                vSys2PeArray [8][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][28].cb_test                                      ;
                vSys2PeArray [8][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][29].cb_test                                      ;
                vSys2PeArray [8][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][30].cb_test                                      ;
                vSys2PeArray [8][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[8][31].cb_test                                      ;
                vSys2PeArray [8][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [8][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[9][0].cb_test                                      ;
                vSys2PeArray [9][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][1].cb_test                                      ;
                vSys2PeArray [9][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][2].cb_test                                      ;
                vSys2PeArray [9][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][3].cb_test                                      ;
                vSys2PeArray [9][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][4].cb_test                                      ;
                vSys2PeArray [9][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][5].cb_test                                      ;
                vSys2PeArray [9][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][6].cb_test                                      ;
                vSys2PeArray [9][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][7].cb_test                                      ;
                vSys2PeArray [9][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][8].cb_test                                      ;
                vSys2PeArray [9][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][9].cb_test                                      ;
                vSys2PeArray [9][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][10].cb_test                                      ;
                vSys2PeArray [9][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][11].cb_test                                      ;
                vSys2PeArray [9][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][12].cb_test                                      ;
                vSys2PeArray [9][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][13].cb_test                                      ;
                vSys2PeArray [9][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][14].cb_test                                      ;
                vSys2PeArray [9][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][15].cb_test                                      ;
                vSys2PeArray [9][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][16].cb_test                                      ;
                vSys2PeArray [9][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][17].cb_test                                      ;
                vSys2PeArray [9][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][18].cb_test                                      ;
                vSys2PeArray [9][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][19].cb_test                                      ;
                vSys2PeArray [9][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][20].cb_test                                      ;
                vSys2PeArray [9][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][21].cb_test                                      ;
                vSys2PeArray [9][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][22].cb_test                                      ;
                vSys2PeArray [9][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][23].cb_test                                      ;
                vSys2PeArray [9][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][24].cb_test                                      ;
                vSys2PeArray [9][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][25].cb_test                                      ;
                vSys2PeArray [9][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][26].cb_test                                      ;
                vSys2PeArray [9][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][27].cb_test                                      ;
                vSys2PeArray [9][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][28].cb_test                                      ;
                vSys2PeArray [9][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][29].cb_test                                      ;
                vSys2PeArray [9][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][30].cb_test                                      ;
                vSys2PeArray [9][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[9][31].cb_test                                      ;
                vSys2PeArray [9][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [9][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[10][0].cb_test                                      ;
                vSys2PeArray [10][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][1].cb_test                                      ;
                vSys2PeArray [10][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][2].cb_test                                      ;
                vSys2PeArray [10][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][3].cb_test                                      ;
                vSys2PeArray [10][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][4].cb_test                                      ;
                vSys2PeArray [10][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][5].cb_test                                      ;
                vSys2PeArray [10][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][6].cb_test                                      ;
                vSys2PeArray [10][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][7].cb_test                                      ;
                vSys2PeArray [10][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][8].cb_test                                      ;
                vSys2PeArray [10][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][9].cb_test                                      ;
                vSys2PeArray [10][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][10].cb_test                                      ;
                vSys2PeArray [10][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][11].cb_test                                      ;
                vSys2PeArray [10][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][12].cb_test                                      ;
                vSys2PeArray [10][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][13].cb_test                                      ;
                vSys2PeArray [10][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][14].cb_test                                      ;
                vSys2PeArray [10][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][15].cb_test                                      ;
                vSys2PeArray [10][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][16].cb_test                                      ;
                vSys2PeArray [10][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][17].cb_test                                      ;
                vSys2PeArray [10][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][18].cb_test                                      ;
                vSys2PeArray [10][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][19].cb_test                                      ;
                vSys2PeArray [10][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][20].cb_test                                      ;
                vSys2PeArray [10][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][21].cb_test                                      ;
                vSys2PeArray [10][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][22].cb_test                                      ;
                vSys2PeArray [10][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][23].cb_test                                      ;
                vSys2PeArray [10][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][24].cb_test                                      ;
                vSys2PeArray [10][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][25].cb_test                                      ;
                vSys2PeArray [10][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][26].cb_test                                      ;
                vSys2PeArray [10][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][27].cb_test                                      ;
                vSys2PeArray [10][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][28].cb_test                                      ;
                vSys2PeArray [10][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][29].cb_test                                      ;
                vSys2PeArray [10][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][30].cb_test                                      ;
                vSys2PeArray [10][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[10][31].cb_test                                      ;
                vSys2PeArray [10][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [10][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[11][0].cb_test                                      ;
                vSys2PeArray [11][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][1].cb_test                                      ;
                vSys2PeArray [11][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][2].cb_test                                      ;
                vSys2PeArray [11][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][3].cb_test                                      ;
                vSys2PeArray [11][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][4].cb_test                                      ;
                vSys2PeArray [11][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][5].cb_test                                      ;
                vSys2PeArray [11][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][6].cb_test                                      ;
                vSys2PeArray [11][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][7].cb_test                                      ;
                vSys2PeArray [11][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][8].cb_test                                      ;
                vSys2PeArray [11][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][9].cb_test                                      ;
                vSys2PeArray [11][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][10].cb_test                                      ;
                vSys2PeArray [11][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][11].cb_test                                      ;
                vSys2PeArray [11][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][12].cb_test                                      ;
                vSys2PeArray [11][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][13].cb_test                                      ;
                vSys2PeArray [11][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][14].cb_test                                      ;
                vSys2PeArray [11][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][15].cb_test                                      ;
                vSys2PeArray [11][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][16].cb_test                                      ;
                vSys2PeArray [11][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][17].cb_test                                      ;
                vSys2PeArray [11][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][18].cb_test                                      ;
                vSys2PeArray [11][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][19].cb_test                                      ;
                vSys2PeArray [11][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][20].cb_test                                      ;
                vSys2PeArray [11][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][21].cb_test                                      ;
                vSys2PeArray [11][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][22].cb_test                                      ;
                vSys2PeArray [11][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][23].cb_test                                      ;
                vSys2PeArray [11][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][24].cb_test                                      ;
                vSys2PeArray [11][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][25].cb_test                                      ;
                vSys2PeArray [11][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][26].cb_test                                      ;
                vSys2PeArray [11][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][27].cb_test                                      ;
                vSys2PeArray [11][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][28].cb_test                                      ;
                vSys2PeArray [11][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][29].cb_test                                      ;
                vSys2PeArray [11][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][30].cb_test                                      ;
                vSys2PeArray [11][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[11][31].cb_test                                      ;
                vSys2PeArray [11][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [11][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[12][0].cb_test                                      ;
                vSys2PeArray [12][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][1].cb_test                                      ;
                vSys2PeArray [12][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][2].cb_test                                      ;
                vSys2PeArray [12][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][3].cb_test                                      ;
                vSys2PeArray [12][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][4].cb_test                                      ;
                vSys2PeArray [12][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][5].cb_test                                      ;
                vSys2PeArray [12][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][6].cb_test                                      ;
                vSys2PeArray [12][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][7].cb_test                                      ;
                vSys2PeArray [12][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][8].cb_test                                      ;
                vSys2PeArray [12][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][9].cb_test                                      ;
                vSys2PeArray [12][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][10].cb_test                                      ;
                vSys2PeArray [12][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][11].cb_test                                      ;
                vSys2PeArray [12][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][12].cb_test                                      ;
                vSys2PeArray [12][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][13].cb_test                                      ;
                vSys2PeArray [12][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][14].cb_test                                      ;
                vSys2PeArray [12][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][15].cb_test                                      ;
                vSys2PeArray [12][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][16].cb_test                                      ;
                vSys2PeArray [12][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][17].cb_test                                      ;
                vSys2PeArray [12][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][18].cb_test                                      ;
                vSys2PeArray [12][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][19].cb_test                                      ;
                vSys2PeArray [12][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][20].cb_test                                      ;
                vSys2PeArray [12][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][21].cb_test                                      ;
                vSys2PeArray [12][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][22].cb_test                                      ;
                vSys2PeArray [12][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][23].cb_test                                      ;
                vSys2PeArray [12][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][24].cb_test                                      ;
                vSys2PeArray [12][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][25].cb_test                                      ;
                vSys2PeArray [12][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][26].cb_test                                      ;
                vSys2PeArray [12][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][27].cb_test                                      ;
                vSys2PeArray [12][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][28].cb_test                                      ;
                vSys2PeArray [12][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][29].cb_test                                      ;
                vSys2PeArray [12][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][30].cb_test                                      ;
                vSys2PeArray [12][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[12][31].cb_test                                      ;
                vSys2PeArray [12][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [12][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[13][0].cb_test                                      ;
                vSys2PeArray [13][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][1].cb_test                                      ;
                vSys2PeArray [13][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][2].cb_test                                      ;
                vSys2PeArray [13][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][3].cb_test                                      ;
                vSys2PeArray [13][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][4].cb_test                                      ;
                vSys2PeArray [13][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][5].cb_test                                      ;
                vSys2PeArray [13][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][6].cb_test                                      ;
                vSys2PeArray [13][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][7].cb_test                                      ;
                vSys2PeArray [13][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][8].cb_test                                      ;
                vSys2PeArray [13][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][9].cb_test                                      ;
                vSys2PeArray [13][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][10].cb_test                                      ;
                vSys2PeArray [13][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][11].cb_test                                      ;
                vSys2PeArray [13][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][12].cb_test                                      ;
                vSys2PeArray [13][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][13].cb_test                                      ;
                vSys2PeArray [13][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][14].cb_test                                      ;
                vSys2PeArray [13][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][15].cb_test                                      ;
                vSys2PeArray [13][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][16].cb_test                                      ;
                vSys2PeArray [13][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][17].cb_test                                      ;
                vSys2PeArray [13][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][18].cb_test                                      ;
                vSys2PeArray [13][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][19].cb_test                                      ;
                vSys2PeArray [13][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][20].cb_test                                      ;
                vSys2PeArray [13][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][21].cb_test                                      ;
                vSys2PeArray [13][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][22].cb_test                                      ;
                vSys2PeArray [13][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][23].cb_test                                      ;
                vSys2PeArray [13][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][24].cb_test                                      ;
                vSys2PeArray [13][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][25].cb_test                                      ;
                vSys2PeArray [13][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][26].cb_test                                      ;
                vSys2PeArray [13][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][27].cb_test                                      ;
                vSys2PeArray [13][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][28].cb_test                                      ;
                vSys2PeArray [13][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][29].cb_test                                      ;
                vSys2PeArray [13][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][30].cb_test                                      ;
                vSys2PeArray [13][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[13][31].cb_test                                      ;
                vSys2PeArray [13][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [13][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[14][0].cb_test                                      ;
                vSys2PeArray [14][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][1].cb_test                                      ;
                vSys2PeArray [14][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][2].cb_test                                      ;
                vSys2PeArray [14][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][3].cb_test                                      ;
                vSys2PeArray [14][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][4].cb_test                                      ;
                vSys2PeArray [14][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][5].cb_test                                      ;
                vSys2PeArray [14][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][6].cb_test                                      ;
                vSys2PeArray [14][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][7].cb_test                                      ;
                vSys2PeArray [14][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][8].cb_test                                      ;
                vSys2PeArray [14][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][9].cb_test                                      ;
                vSys2PeArray [14][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][10].cb_test                                      ;
                vSys2PeArray [14][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][11].cb_test                                      ;
                vSys2PeArray [14][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][12].cb_test                                      ;
                vSys2PeArray [14][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][13].cb_test                                      ;
                vSys2PeArray [14][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][14].cb_test                                      ;
                vSys2PeArray [14][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][15].cb_test                                      ;
                vSys2PeArray [14][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][16].cb_test                                      ;
                vSys2PeArray [14][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][17].cb_test                                      ;
                vSys2PeArray [14][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][18].cb_test                                      ;
                vSys2PeArray [14][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][19].cb_test                                      ;
                vSys2PeArray [14][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][20].cb_test                                      ;
                vSys2PeArray [14][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][21].cb_test                                      ;
                vSys2PeArray [14][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][22].cb_test                                      ;
                vSys2PeArray [14][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][23].cb_test                                      ;
                vSys2PeArray [14][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][24].cb_test                                      ;
                vSys2PeArray [14][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][25].cb_test                                      ;
                vSys2PeArray [14][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][26].cb_test                                      ;
                vSys2PeArray [14][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][27].cb_test                                      ;
                vSys2PeArray [14][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][28].cb_test                                      ;
                vSys2PeArray [14][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][29].cb_test                                      ;
                vSys2PeArray [14][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][30].cb_test                                      ;
                vSys2PeArray [14][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[14][31].cb_test                                      ;
                vSys2PeArray [14][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [14][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[15][0].cb_test                                      ;
                vSys2PeArray [15][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][1].cb_test                                      ;
                vSys2PeArray [15][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][2].cb_test                                      ;
                vSys2PeArray [15][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][3].cb_test                                      ;
                vSys2PeArray [15][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][4].cb_test                                      ;
                vSys2PeArray [15][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][5].cb_test                                      ;
                vSys2PeArray [15][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][6].cb_test                                      ;
                vSys2PeArray [15][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][7].cb_test                                      ;
                vSys2PeArray [15][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][8].cb_test                                      ;
                vSys2PeArray [15][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][9].cb_test                                      ;
                vSys2PeArray [15][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][10].cb_test                                      ;
                vSys2PeArray [15][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][11].cb_test                                      ;
                vSys2PeArray [15][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][12].cb_test                                      ;
                vSys2PeArray [15][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][13].cb_test                                      ;
                vSys2PeArray [15][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][14].cb_test                                      ;
                vSys2PeArray [15][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][15].cb_test                                      ;
                vSys2PeArray [15][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][16].cb_test                                      ;
                vSys2PeArray [15][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][17].cb_test                                      ;
                vSys2PeArray [15][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][18].cb_test                                      ;
                vSys2PeArray [15][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][19].cb_test                                      ;
                vSys2PeArray [15][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][20].cb_test                                      ;
                vSys2PeArray [15][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][21].cb_test                                      ;
                vSys2PeArray [15][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][22].cb_test                                      ;
                vSys2PeArray [15][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][23].cb_test                                      ;
                vSys2PeArray [15][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][24].cb_test                                      ;
                vSys2PeArray [15][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][25].cb_test                                      ;
                vSys2PeArray [15][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][26].cb_test                                      ;
                vSys2PeArray [15][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][27].cb_test                                      ;
                vSys2PeArray [15][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][28].cb_test                                      ;
                vSys2PeArray [15][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][29].cb_test                                      ;
                vSys2PeArray [15][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][30].cb_test                                      ;
                vSys2PeArray [15][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[15][31].cb_test                                      ;
                vSys2PeArray [15][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [15][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[16][0].cb_test                                      ;
                vSys2PeArray [16][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][1].cb_test                                      ;
                vSys2PeArray [16][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][2].cb_test                                      ;
                vSys2PeArray [16][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][3].cb_test                                      ;
                vSys2PeArray [16][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][4].cb_test                                      ;
                vSys2PeArray [16][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][5].cb_test                                      ;
                vSys2PeArray [16][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][6].cb_test                                      ;
                vSys2PeArray [16][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][7].cb_test                                      ;
                vSys2PeArray [16][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][8].cb_test                                      ;
                vSys2PeArray [16][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][9].cb_test                                      ;
                vSys2PeArray [16][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][10].cb_test                                      ;
                vSys2PeArray [16][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][11].cb_test                                      ;
                vSys2PeArray [16][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][12].cb_test                                      ;
                vSys2PeArray [16][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][13].cb_test                                      ;
                vSys2PeArray [16][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][14].cb_test                                      ;
                vSys2PeArray [16][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][15].cb_test                                      ;
                vSys2PeArray [16][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][16].cb_test                                      ;
                vSys2PeArray [16][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][17].cb_test                                      ;
                vSys2PeArray [16][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][18].cb_test                                      ;
                vSys2PeArray [16][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][19].cb_test                                      ;
                vSys2PeArray [16][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][20].cb_test                                      ;
                vSys2PeArray [16][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][21].cb_test                                      ;
                vSys2PeArray [16][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][22].cb_test                                      ;
                vSys2PeArray [16][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][23].cb_test                                      ;
                vSys2PeArray [16][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][24].cb_test                                      ;
                vSys2PeArray [16][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][25].cb_test                                      ;
                vSys2PeArray [16][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][26].cb_test                                      ;
                vSys2PeArray [16][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][27].cb_test                                      ;
                vSys2PeArray [16][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][28].cb_test                                      ;
                vSys2PeArray [16][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][29].cb_test                                      ;
                vSys2PeArray [16][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][30].cb_test                                      ;
                vSys2PeArray [16][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[16][31].cb_test                                      ;
                vSys2PeArray [16][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [16][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[17][0].cb_test                                      ;
                vSys2PeArray [17][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][1].cb_test                                      ;
                vSys2PeArray [17][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][2].cb_test                                      ;
                vSys2PeArray [17][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][3].cb_test                                      ;
                vSys2PeArray [17][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][4].cb_test                                      ;
                vSys2PeArray [17][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][5].cb_test                                      ;
                vSys2PeArray [17][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][6].cb_test                                      ;
                vSys2PeArray [17][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][7].cb_test                                      ;
                vSys2PeArray [17][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][8].cb_test                                      ;
                vSys2PeArray [17][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][9].cb_test                                      ;
                vSys2PeArray [17][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][10].cb_test                                      ;
                vSys2PeArray [17][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][11].cb_test                                      ;
                vSys2PeArray [17][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][12].cb_test                                      ;
                vSys2PeArray [17][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][13].cb_test                                      ;
                vSys2PeArray [17][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][14].cb_test                                      ;
                vSys2PeArray [17][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][15].cb_test                                      ;
                vSys2PeArray [17][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][16].cb_test                                      ;
                vSys2PeArray [17][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][17].cb_test                                      ;
                vSys2PeArray [17][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][18].cb_test                                      ;
                vSys2PeArray [17][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][19].cb_test                                      ;
                vSys2PeArray [17][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][20].cb_test                                      ;
                vSys2PeArray [17][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][21].cb_test                                      ;
                vSys2PeArray [17][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][22].cb_test                                      ;
                vSys2PeArray [17][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][23].cb_test                                      ;
                vSys2PeArray [17][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][24].cb_test                                      ;
                vSys2PeArray [17][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][25].cb_test                                      ;
                vSys2PeArray [17][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][26].cb_test                                      ;
                vSys2PeArray [17][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][27].cb_test                                      ;
                vSys2PeArray [17][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][28].cb_test                                      ;
                vSys2PeArray [17][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][29].cb_test                                      ;
                vSys2PeArray [17][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][30].cb_test                                      ;
                vSys2PeArray [17][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[17][31].cb_test                                      ;
                vSys2PeArray [17][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [17][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[18][0].cb_test                                      ;
                vSys2PeArray [18][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][1].cb_test                                      ;
                vSys2PeArray [18][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][2].cb_test                                      ;
                vSys2PeArray [18][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][3].cb_test                                      ;
                vSys2PeArray [18][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][4].cb_test                                      ;
                vSys2PeArray [18][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][5].cb_test                                      ;
                vSys2PeArray [18][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][6].cb_test                                      ;
                vSys2PeArray [18][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][7].cb_test                                      ;
                vSys2PeArray [18][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][8].cb_test                                      ;
                vSys2PeArray [18][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][9].cb_test                                      ;
                vSys2PeArray [18][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][10].cb_test                                      ;
                vSys2PeArray [18][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][11].cb_test                                      ;
                vSys2PeArray [18][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][12].cb_test                                      ;
                vSys2PeArray [18][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][13].cb_test                                      ;
                vSys2PeArray [18][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][14].cb_test                                      ;
                vSys2PeArray [18][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][15].cb_test                                      ;
                vSys2PeArray [18][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][16].cb_test                                      ;
                vSys2PeArray [18][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][17].cb_test                                      ;
                vSys2PeArray [18][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][18].cb_test                                      ;
                vSys2PeArray [18][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][19].cb_test                                      ;
                vSys2PeArray [18][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][20].cb_test                                      ;
                vSys2PeArray [18][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][21].cb_test                                      ;
                vSys2PeArray [18][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][22].cb_test                                      ;
                vSys2PeArray [18][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][23].cb_test                                      ;
                vSys2PeArray [18][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][24].cb_test                                      ;
                vSys2PeArray [18][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][25].cb_test                                      ;
                vSys2PeArray [18][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][26].cb_test                                      ;
                vSys2PeArray [18][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][27].cb_test                                      ;
                vSys2PeArray [18][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][28].cb_test                                      ;
                vSys2PeArray [18][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][29].cb_test                                      ;
                vSys2PeArray [18][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][30].cb_test                                      ;
                vSys2PeArray [18][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[18][31].cb_test                                      ;
                vSys2PeArray [18][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [18][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[19][0].cb_test                                      ;
                vSys2PeArray [19][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][1].cb_test                                      ;
                vSys2PeArray [19][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][2].cb_test                                      ;
                vSys2PeArray [19][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][3].cb_test                                      ;
                vSys2PeArray [19][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][4].cb_test                                      ;
                vSys2PeArray [19][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][5].cb_test                                      ;
                vSys2PeArray [19][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][6].cb_test                                      ;
                vSys2PeArray [19][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][7].cb_test                                      ;
                vSys2PeArray [19][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][8].cb_test                                      ;
                vSys2PeArray [19][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][9].cb_test                                      ;
                vSys2PeArray [19][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][10].cb_test                                      ;
                vSys2PeArray [19][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][11].cb_test                                      ;
                vSys2PeArray [19][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][12].cb_test                                      ;
                vSys2PeArray [19][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][13].cb_test                                      ;
                vSys2PeArray [19][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][14].cb_test                                      ;
                vSys2PeArray [19][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][15].cb_test                                      ;
                vSys2PeArray [19][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][16].cb_test                                      ;
                vSys2PeArray [19][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][17].cb_test                                      ;
                vSys2PeArray [19][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][18].cb_test                                      ;
                vSys2PeArray [19][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][19].cb_test                                      ;
                vSys2PeArray [19][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][20].cb_test                                      ;
                vSys2PeArray [19][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][21].cb_test                                      ;
                vSys2PeArray [19][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][22].cb_test                                      ;
                vSys2PeArray [19][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][23].cb_test                                      ;
                vSys2PeArray [19][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][24].cb_test                                      ;
                vSys2PeArray [19][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][25].cb_test                                      ;
                vSys2PeArray [19][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][26].cb_test                                      ;
                vSys2PeArray [19][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][27].cb_test                                      ;
                vSys2PeArray [19][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][28].cb_test                                      ;
                vSys2PeArray [19][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][29].cb_test                                      ;
                vSys2PeArray [19][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][30].cb_test                                      ;
                vSys2PeArray [19][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[19][31].cb_test                                      ;
                vSys2PeArray [19][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [19][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[20][0].cb_test                                      ;
                vSys2PeArray [20][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][1].cb_test                                      ;
                vSys2PeArray [20][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][2].cb_test                                      ;
                vSys2PeArray [20][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][3].cb_test                                      ;
                vSys2PeArray [20][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][4].cb_test                                      ;
                vSys2PeArray [20][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][5].cb_test                                      ;
                vSys2PeArray [20][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][6].cb_test                                      ;
                vSys2PeArray [20][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][7].cb_test                                      ;
                vSys2PeArray [20][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][8].cb_test                                      ;
                vSys2PeArray [20][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][9].cb_test                                      ;
                vSys2PeArray [20][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][10].cb_test                                      ;
                vSys2PeArray [20][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][11].cb_test                                      ;
                vSys2PeArray [20][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][12].cb_test                                      ;
                vSys2PeArray [20][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][13].cb_test                                      ;
                vSys2PeArray [20][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][14].cb_test                                      ;
                vSys2PeArray [20][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][15].cb_test                                      ;
                vSys2PeArray [20][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][16].cb_test                                      ;
                vSys2PeArray [20][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][17].cb_test                                      ;
                vSys2PeArray [20][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][18].cb_test                                      ;
                vSys2PeArray [20][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][19].cb_test                                      ;
                vSys2PeArray [20][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][20].cb_test                                      ;
                vSys2PeArray [20][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][21].cb_test                                      ;
                vSys2PeArray [20][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][22].cb_test                                      ;
                vSys2PeArray [20][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][23].cb_test                                      ;
                vSys2PeArray [20][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][24].cb_test                                      ;
                vSys2PeArray [20][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][25].cb_test                                      ;
                vSys2PeArray [20][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][26].cb_test                                      ;
                vSys2PeArray [20][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][27].cb_test                                      ;
                vSys2PeArray [20][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][28].cb_test                                      ;
                vSys2PeArray [20][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][29].cb_test                                      ;
                vSys2PeArray [20][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][30].cb_test                                      ;
                vSys2PeArray [20][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[20][31].cb_test                                      ;
                vSys2PeArray [20][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [20][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[21][0].cb_test                                      ;
                vSys2PeArray [21][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][1].cb_test                                      ;
                vSys2PeArray [21][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][2].cb_test                                      ;
                vSys2PeArray [21][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][3].cb_test                                      ;
                vSys2PeArray [21][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][4].cb_test                                      ;
                vSys2PeArray [21][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][5].cb_test                                      ;
                vSys2PeArray [21][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][6].cb_test                                      ;
                vSys2PeArray [21][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][7].cb_test                                      ;
                vSys2PeArray [21][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][8].cb_test                                      ;
                vSys2PeArray [21][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][9].cb_test                                      ;
                vSys2PeArray [21][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][10].cb_test                                      ;
                vSys2PeArray [21][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][11].cb_test                                      ;
                vSys2PeArray [21][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][12].cb_test                                      ;
                vSys2PeArray [21][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][13].cb_test                                      ;
                vSys2PeArray [21][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][14].cb_test                                      ;
                vSys2PeArray [21][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][15].cb_test                                      ;
                vSys2PeArray [21][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][16].cb_test                                      ;
                vSys2PeArray [21][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][17].cb_test                                      ;
                vSys2PeArray [21][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][18].cb_test                                      ;
                vSys2PeArray [21][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][19].cb_test                                      ;
                vSys2PeArray [21][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][20].cb_test                                      ;
                vSys2PeArray [21][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][21].cb_test                                      ;
                vSys2PeArray [21][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][22].cb_test                                      ;
                vSys2PeArray [21][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][23].cb_test                                      ;
                vSys2PeArray [21][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][24].cb_test                                      ;
                vSys2PeArray [21][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][25].cb_test                                      ;
                vSys2PeArray [21][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][26].cb_test                                      ;
                vSys2PeArray [21][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][27].cb_test                                      ;
                vSys2PeArray [21][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][28].cb_test                                      ;
                vSys2PeArray [21][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][29].cb_test                                      ;
                vSys2PeArray [21][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][30].cb_test                                      ;
                vSys2PeArray [21][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[21][31].cb_test                                      ;
                vSys2PeArray [21][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [21][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[22][0].cb_test                                      ;
                vSys2PeArray [22][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][1].cb_test                                      ;
                vSys2PeArray [22][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][2].cb_test                                      ;
                vSys2PeArray [22][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][3].cb_test                                      ;
                vSys2PeArray [22][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][4].cb_test                                      ;
                vSys2PeArray [22][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][5].cb_test                                      ;
                vSys2PeArray [22][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][6].cb_test                                      ;
                vSys2PeArray [22][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][7].cb_test                                      ;
                vSys2PeArray [22][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][8].cb_test                                      ;
                vSys2PeArray [22][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][9].cb_test                                      ;
                vSys2PeArray [22][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][10].cb_test                                      ;
                vSys2PeArray [22][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][11].cb_test                                      ;
                vSys2PeArray [22][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][12].cb_test                                      ;
                vSys2PeArray [22][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][13].cb_test                                      ;
                vSys2PeArray [22][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][14].cb_test                                      ;
                vSys2PeArray [22][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][15].cb_test                                      ;
                vSys2PeArray [22][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][16].cb_test                                      ;
                vSys2PeArray [22][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][17].cb_test                                      ;
                vSys2PeArray [22][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][18].cb_test                                      ;
                vSys2PeArray [22][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][19].cb_test                                      ;
                vSys2PeArray [22][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][20].cb_test                                      ;
                vSys2PeArray [22][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][21].cb_test                                      ;
                vSys2PeArray [22][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][22].cb_test                                      ;
                vSys2PeArray [22][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][23].cb_test                                      ;
                vSys2PeArray [22][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][24].cb_test                                      ;
                vSys2PeArray [22][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][25].cb_test                                      ;
                vSys2PeArray [22][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][26].cb_test                                      ;
                vSys2PeArray [22][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][27].cb_test                                      ;
                vSys2PeArray [22][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][28].cb_test                                      ;
                vSys2PeArray [22][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][29].cb_test                                      ;
                vSys2PeArray [22][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][30].cb_test                                      ;
                vSys2PeArray [22][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[22][31].cb_test                                      ;
                vSys2PeArray [22][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [22][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[23][0].cb_test                                      ;
                vSys2PeArray [23][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][1].cb_test                                      ;
                vSys2PeArray [23][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][2].cb_test                                      ;
                vSys2PeArray [23][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][3].cb_test                                      ;
                vSys2PeArray [23][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][4].cb_test                                      ;
                vSys2PeArray [23][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][5].cb_test                                      ;
                vSys2PeArray [23][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][6].cb_test                                      ;
                vSys2PeArray [23][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][7].cb_test                                      ;
                vSys2PeArray [23][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][8].cb_test                                      ;
                vSys2PeArray [23][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][9].cb_test                                      ;
                vSys2PeArray [23][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][10].cb_test                                      ;
                vSys2PeArray [23][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][11].cb_test                                      ;
                vSys2PeArray [23][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][12].cb_test                                      ;
                vSys2PeArray [23][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][13].cb_test                                      ;
                vSys2PeArray [23][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][14].cb_test                                      ;
                vSys2PeArray [23][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][15].cb_test                                      ;
                vSys2PeArray [23][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][16].cb_test                                      ;
                vSys2PeArray [23][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][17].cb_test                                      ;
                vSys2PeArray [23][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][18].cb_test                                      ;
                vSys2PeArray [23][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][19].cb_test                                      ;
                vSys2PeArray [23][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][20].cb_test                                      ;
                vSys2PeArray [23][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][21].cb_test                                      ;
                vSys2PeArray [23][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][22].cb_test                                      ;
                vSys2PeArray [23][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][23].cb_test                                      ;
                vSys2PeArray [23][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][24].cb_test                                      ;
                vSys2PeArray [23][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][25].cb_test                                      ;
                vSys2PeArray [23][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][26].cb_test                                      ;
                vSys2PeArray [23][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][27].cb_test                                      ;
                vSys2PeArray [23][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][28].cb_test                                      ;
                vSys2PeArray [23][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][29].cb_test                                      ;
                vSys2PeArray [23][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][30].cb_test                                      ;
                vSys2PeArray [23][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[23][31].cb_test                                      ;
                vSys2PeArray [23][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [23][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[24][0].cb_test                                      ;
                vSys2PeArray [24][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][1].cb_test                                      ;
                vSys2PeArray [24][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][2].cb_test                                      ;
                vSys2PeArray [24][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][3].cb_test                                      ;
                vSys2PeArray [24][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][4].cb_test                                      ;
                vSys2PeArray [24][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][5].cb_test                                      ;
                vSys2PeArray [24][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][6].cb_test                                      ;
                vSys2PeArray [24][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][7].cb_test                                      ;
                vSys2PeArray [24][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][8].cb_test                                      ;
                vSys2PeArray [24][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][9].cb_test                                      ;
                vSys2PeArray [24][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][10].cb_test                                      ;
                vSys2PeArray [24][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][11].cb_test                                      ;
                vSys2PeArray [24][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][12].cb_test                                      ;
                vSys2PeArray [24][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][13].cb_test                                      ;
                vSys2PeArray [24][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][14].cb_test                                      ;
                vSys2PeArray [24][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][15].cb_test                                      ;
                vSys2PeArray [24][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][16].cb_test                                      ;
                vSys2PeArray [24][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][17].cb_test                                      ;
                vSys2PeArray [24][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][18].cb_test                                      ;
                vSys2PeArray [24][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][19].cb_test                                      ;
                vSys2PeArray [24][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][20].cb_test                                      ;
                vSys2PeArray [24][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][21].cb_test                                      ;
                vSys2PeArray [24][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][22].cb_test                                      ;
                vSys2PeArray [24][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][23].cb_test                                      ;
                vSys2PeArray [24][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][24].cb_test                                      ;
                vSys2PeArray [24][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][25].cb_test                                      ;
                vSys2PeArray [24][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][26].cb_test                                      ;
                vSys2PeArray [24][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][27].cb_test                                      ;
                vSys2PeArray [24][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][28].cb_test                                      ;
                vSys2PeArray [24][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][29].cb_test                                      ;
                vSys2PeArray [24][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][30].cb_test                                      ;
                vSys2PeArray [24][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[24][31].cb_test                                      ;
                vSys2PeArray [24][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [24][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[25][0].cb_test                                      ;
                vSys2PeArray [25][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][1].cb_test                                      ;
                vSys2PeArray [25][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][2].cb_test                                      ;
                vSys2PeArray [25][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][3].cb_test                                      ;
                vSys2PeArray [25][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][4].cb_test                                      ;
                vSys2PeArray [25][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][5].cb_test                                      ;
                vSys2PeArray [25][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][6].cb_test                                      ;
                vSys2PeArray [25][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][7].cb_test                                      ;
                vSys2PeArray [25][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][8].cb_test                                      ;
                vSys2PeArray [25][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][9].cb_test                                      ;
                vSys2PeArray [25][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][10].cb_test                                      ;
                vSys2PeArray [25][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][11].cb_test                                      ;
                vSys2PeArray [25][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][12].cb_test                                      ;
                vSys2PeArray [25][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][13].cb_test                                      ;
                vSys2PeArray [25][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][14].cb_test                                      ;
                vSys2PeArray [25][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][15].cb_test                                      ;
                vSys2PeArray [25][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][16].cb_test                                      ;
                vSys2PeArray [25][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][17].cb_test                                      ;
                vSys2PeArray [25][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][18].cb_test                                      ;
                vSys2PeArray [25][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][19].cb_test                                      ;
                vSys2PeArray [25][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][20].cb_test                                      ;
                vSys2PeArray [25][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][21].cb_test                                      ;
                vSys2PeArray [25][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][22].cb_test                                      ;
                vSys2PeArray [25][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][23].cb_test                                      ;
                vSys2PeArray [25][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][24].cb_test                                      ;
                vSys2PeArray [25][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][25].cb_test                                      ;
                vSys2PeArray [25][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][26].cb_test                                      ;
                vSys2PeArray [25][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][27].cb_test                                      ;
                vSys2PeArray [25][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][28].cb_test                                      ;
                vSys2PeArray [25][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][29].cb_test                                      ;
                vSys2PeArray [25][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][30].cb_test                                      ;
                vSys2PeArray [25][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[25][31].cb_test                                      ;
                vSys2PeArray [25][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [25][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[26][0].cb_test                                      ;
                vSys2PeArray [26][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][1].cb_test                                      ;
                vSys2PeArray [26][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][2].cb_test                                      ;
                vSys2PeArray [26][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][3].cb_test                                      ;
                vSys2PeArray [26][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][4].cb_test                                      ;
                vSys2PeArray [26][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][5].cb_test                                      ;
                vSys2PeArray [26][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][6].cb_test                                      ;
                vSys2PeArray [26][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][7].cb_test                                      ;
                vSys2PeArray [26][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][8].cb_test                                      ;
                vSys2PeArray [26][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][9].cb_test                                      ;
                vSys2PeArray [26][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][10].cb_test                                      ;
                vSys2PeArray [26][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][11].cb_test                                      ;
                vSys2PeArray [26][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][12].cb_test                                      ;
                vSys2PeArray [26][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][13].cb_test                                      ;
                vSys2PeArray [26][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][14].cb_test                                      ;
                vSys2PeArray [26][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][15].cb_test                                      ;
                vSys2PeArray [26][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][16].cb_test                                      ;
                vSys2PeArray [26][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][17].cb_test                                      ;
                vSys2PeArray [26][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][18].cb_test                                      ;
                vSys2PeArray [26][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][19].cb_test                                      ;
                vSys2PeArray [26][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][20].cb_test                                      ;
                vSys2PeArray [26][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][21].cb_test                                      ;
                vSys2PeArray [26][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][22].cb_test                                      ;
                vSys2PeArray [26][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][23].cb_test                                      ;
                vSys2PeArray [26][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][24].cb_test                                      ;
                vSys2PeArray [26][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][25].cb_test                                      ;
                vSys2PeArray [26][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][26].cb_test                                      ;
                vSys2PeArray [26][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][27].cb_test                                      ;
                vSys2PeArray [26][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][28].cb_test                                      ;
                vSys2PeArray [26][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][29].cb_test                                      ;
                vSys2PeArray [26][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][30].cb_test                                      ;
                vSys2PeArray [26][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[26][31].cb_test                                      ;
                vSys2PeArray [26][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [26][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[27][0].cb_test                                      ;
                vSys2PeArray [27][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][1].cb_test                                      ;
                vSys2PeArray [27][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][2].cb_test                                      ;
                vSys2PeArray [27][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][3].cb_test                                      ;
                vSys2PeArray [27][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][4].cb_test                                      ;
                vSys2PeArray [27][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][5].cb_test                                      ;
                vSys2PeArray [27][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][6].cb_test                                      ;
                vSys2PeArray [27][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][7].cb_test                                      ;
                vSys2PeArray [27][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][8].cb_test                                      ;
                vSys2PeArray [27][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][9].cb_test                                      ;
                vSys2PeArray [27][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][10].cb_test                                      ;
                vSys2PeArray [27][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][11].cb_test                                      ;
                vSys2PeArray [27][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][12].cb_test                                      ;
                vSys2PeArray [27][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][13].cb_test                                      ;
                vSys2PeArray [27][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][14].cb_test                                      ;
                vSys2PeArray [27][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][15].cb_test                                      ;
                vSys2PeArray [27][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][16].cb_test                                      ;
                vSys2PeArray [27][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][17].cb_test                                      ;
                vSys2PeArray [27][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][18].cb_test                                      ;
                vSys2PeArray [27][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][19].cb_test                                      ;
                vSys2PeArray [27][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][20].cb_test                                      ;
                vSys2PeArray [27][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][21].cb_test                                      ;
                vSys2PeArray [27][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][22].cb_test                                      ;
                vSys2PeArray [27][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][23].cb_test                                      ;
                vSys2PeArray [27][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][24].cb_test                                      ;
                vSys2PeArray [27][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][25].cb_test                                      ;
                vSys2PeArray [27][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][26].cb_test                                      ;
                vSys2PeArray [27][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][27].cb_test                                      ;
                vSys2PeArray [27][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][28].cb_test                                      ;
                vSys2PeArray [27][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][29].cb_test                                      ;
                vSys2PeArray [27][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][30].cb_test                                      ;
                vSys2PeArray [27][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[27][31].cb_test                                      ;
                vSys2PeArray [27][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [27][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[28][0].cb_test                                      ;
                vSys2PeArray [28][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][1].cb_test                                      ;
                vSys2PeArray [28][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][2].cb_test                                      ;
                vSys2PeArray [28][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][3].cb_test                                      ;
                vSys2PeArray [28][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][4].cb_test                                      ;
                vSys2PeArray [28][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][5].cb_test                                      ;
                vSys2PeArray [28][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][6].cb_test                                      ;
                vSys2PeArray [28][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][7].cb_test                                      ;
                vSys2PeArray [28][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][8].cb_test                                      ;
                vSys2PeArray [28][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][9].cb_test                                      ;
                vSys2PeArray [28][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][10].cb_test                                      ;
                vSys2PeArray [28][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][11].cb_test                                      ;
                vSys2PeArray [28][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][12].cb_test                                      ;
                vSys2PeArray [28][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][13].cb_test                                      ;
                vSys2PeArray [28][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][14].cb_test                                      ;
                vSys2PeArray [28][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][15].cb_test                                      ;
                vSys2PeArray [28][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][16].cb_test                                      ;
                vSys2PeArray [28][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][17].cb_test                                      ;
                vSys2PeArray [28][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][18].cb_test                                      ;
                vSys2PeArray [28][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][19].cb_test                                      ;
                vSys2PeArray [28][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][20].cb_test                                      ;
                vSys2PeArray [28][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][21].cb_test                                      ;
                vSys2PeArray [28][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][22].cb_test                                      ;
                vSys2PeArray [28][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][23].cb_test                                      ;
                vSys2PeArray [28][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][24].cb_test                                      ;
                vSys2PeArray [28][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][25].cb_test                                      ;
                vSys2PeArray [28][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][26].cb_test                                      ;
                vSys2PeArray [28][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][27].cb_test                                      ;
                vSys2PeArray [28][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][28].cb_test                                      ;
                vSys2PeArray [28][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][29].cb_test                                      ;
                vSys2PeArray [28][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][30].cb_test                                      ;
                vSys2PeArray [28][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[28][31].cb_test                                      ;
                vSys2PeArray [28][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [28][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[29][0].cb_test                                      ;
                vSys2PeArray [29][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][1].cb_test                                      ;
                vSys2PeArray [29][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][2].cb_test                                      ;
                vSys2PeArray [29][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][3].cb_test                                      ;
                vSys2PeArray [29][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][4].cb_test                                      ;
                vSys2PeArray [29][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][5].cb_test                                      ;
                vSys2PeArray [29][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][6].cb_test                                      ;
                vSys2PeArray [29][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][7].cb_test                                      ;
                vSys2PeArray [29][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][8].cb_test                                      ;
                vSys2PeArray [29][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][9].cb_test                                      ;
                vSys2PeArray [29][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][10].cb_test                                      ;
                vSys2PeArray [29][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][11].cb_test                                      ;
                vSys2PeArray [29][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][12].cb_test                                      ;
                vSys2PeArray [29][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][13].cb_test                                      ;
                vSys2PeArray [29][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][14].cb_test                                      ;
                vSys2PeArray [29][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][15].cb_test                                      ;
                vSys2PeArray [29][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][16].cb_test                                      ;
                vSys2PeArray [29][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][17].cb_test                                      ;
                vSys2PeArray [29][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][18].cb_test                                      ;
                vSys2PeArray [29][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][19].cb_test                                      ;
                vSys2PeArray [29][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][20].cb_test                                      ;
                vSys2PeArray [29][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][21].cb_test                                      ;
                vSys2PeArray [29][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][22].cb_test                                      ;
                vSys2PeArray [29][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][23].cb_test                                      ;
                vSys2PeArray [29][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][24].cb_test                                      ;
                vSys2PeArray [29][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][25].cb_test                                      ;
                vSys2PeArray [29][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][26].cb_test                                      ;
                vSys2PeArray [29][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][27].cb_test                                      ;
                vSys2PeArray [29][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][28].cb_test                                      ;
                vSys2PeArray [29][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][29].cb_test                                      ;
                vSys2PeArray [29][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][30].cb_test                                      ;
                vSys2PeArray [29][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[29][31].cb_test                                      ;
                vSys2PeArray [29][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [29][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[30][0].cb_test                                      ;
                vSys2PeArray [30][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][1].cb_test                                      ;
                vSys2PeArray [30][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][2].cb_test                                      ;
                vSys2PeArray [30][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][3].cb_test                                      ;
                vSys2PeArray [30][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][4].cb_test                                      ;
                vSys2PeArray [30][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][5].cb_test                                      ;
                vSys2PeArray [30][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][6].cb_test                                      ;
                vSys2PeArray [30][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][7].cb_test                                      ;
                vSys2PeArray [30][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][8].cb_test                                      ;
                vSys2PeArray [30][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][9].cb_test                                      ;
                vSys2PeArray [30][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][10].cb_test                                      ;
                vSys2PeArray [30][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][11].cb_test                                      ;
                vSys2PeArray [30][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][12].cb_test                                      ;
                vSys2PeArray [30][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][13].cb_test                                      ;
                vSys2PeArray [30][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][14].cb_test                                      ;
                vSys2PeArray [30][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][15].cb_test                                      ;
                vSys2PeArray [30][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][16].cb_test                                      ;
                vSys2PeArray [30][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][17].cb_test                                      ;
                vSys2PeArray [30][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][18].cb_test                                      ;
                vSys2PeArray [30][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][19].cb_test                                      ;
                vSys2PeArray [30][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][20].cb_test                                      ;
                vSys2PeArray [30][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][21].cb_test                                      ;
                vSys2PeArray [30][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][22].cb_test                                      ;
                vSys2PeArray [30][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][23].cb_test                                      ;
                vSys2PeArray [30][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][24].cb_test                                      ;
                vSys2PeArray [30][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][25].cb_test                                      ;
                vSys2PeArray [30][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][26].cb_test                                      ;
                vSys2PeArray [30][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][27].cb_test                                      ;
                vSys2PeArray [30][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][28].cb_test                                      ;
                vSys2PeArray [30][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][29].cb_test                                      ;
                vSys2PeArray [30][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][30].cb_test                                      ;
                vSys2PeArray [30][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[30][31].cb_test                                      ;
                vSys2PeArray [30][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [30][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[31][0].cb_test                                      ;
                vSys2PeArray [31][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][1].cb_test                                      ;
                vSys2PeArray [31][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][2].cb_test                                      ;
                vSys2PeArray [31][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][3].cb_test                                      ;
                vSys2PeArray [31][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][4].cb_test                                      ;
                vSys2PeArray [31][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][5].cb_test                                      ;
                vSys2PeArray [31][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][6].cb_test                                      ;
                vSys2PeArray [31][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][7].cb_test                                      ;
                vSys2PeArray [31][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][8].cb_test                                      ;
                vSys2PeArray [31][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][9].cb_test                                      ;
                vSys2PeArray [31][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][10].cb_test                                      ;
                vSys2PeArray [31][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][11].cb_test                                      ;
                vSys2PeArray [31][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][12].cb_test                                      ;
                vSys2PeArray [31][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][13].cb_test                                      ;
                vSys2PeArray [31][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][14].cb_test                                      ;
                vSys2PeArray [31][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][15].cb_test                                      ;
                vSys2PeArray [31][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][16].cb_test                                      ;
                vSys2PeArray [31][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][17].cb_test                                      ;
                vSys2PeArray [31][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][18].cb_test                                      ;
                vSys2PeArray [31][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][19].cb_test                                      ;
                vSys2PeArray [31][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][20].cb_test                                      ;
                vSys2PeArray [31][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][21].cb_test                                      ;
                vSys2PeArray [31][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][22].cb_test                                      ;
                vSys2PeArray [31][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][23].cb_test                                      ;
                vSys2PeArray [31][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][24].cb_test                                      ;
                vSys2PeArray [31][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][25].cb_test                                      ;
                vSys2PeArray [31][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][26].cb_test                                      ;
                vSys2PeArray [31][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][27].cb_test                                      ;
                vSys2PeArray [31][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][28].cb_test                                      ;
                vSys2PeArray [31][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][29].cb_test                                      ;
                vSys2PeArray [31][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][30].cb_test                                      ;
                vSys2PeArray [31][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[31][31].cb_test                                      ;
                vSys2PeArray [31][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [31][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[32][0].cb_test                                      ;
                vSys2PeArray [32][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][1].cb_test                                      ;
                vSys2PeArray [32][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][2].cb_test                                      ;
                vSys2PeArray [32][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][3].cb_test                                      ;
                vSys2PeArray [32][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][4].cb_test                                      ;
                vSys2PeArray [32][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][5].cb_test                                      ;
                vSys2PeArray [32][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][6].cb_test                                      ;
                vSys2PeArray [32][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][7].cb_test                                      ;
                vSys2PeArray [32][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][8].cb_test                                      ;
                vSys2PeArray [32][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][9].cb_test                                      ;
                vSys2PeArray [32][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][10].cb_test                                      ;
                vSys2PeArray [32][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][11].cb_test                                      ;
                vSys2PeArray [32][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][12].cb_test                                      ;
                vSys2PeArray [32][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][13].cb_test                                      ;
                vSys2PeArray [32][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][14].cb_test                                      ;
                vSys2PeArray [32][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][15].cb_test                                      ;
                vSys2PeArray [32][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][16].cb_test                                      ;
                vSys2PeArray [32][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][17].cb_test                                      ;
                vSys2PeArray [32][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][18].cb_test                                      ;
                vSys2PeArray [32][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][19].cb_test                                      ;
                vSys2PeArray [32][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][20].cb_test                                      ;
                vSys2PeArray [32][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][21].cb_test                                      ;
                vSys2PeArray [32][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][22].cb_test                                      ;
                vSys2PeArray [32][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][23].cb_test                                      ;
                vSys2PeArray [32][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][24].cb_test                                      ;
                vSys2PeArray [32][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][25].cb_test                                      ;
                vSys2PeArray [32][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][26].cb_test                                      ;
                vSys2PeArray [32][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][27].cb_test                                      ;
                vSys2PeArray [32][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][28].cb_test                                      ;
                vSys2PeArray [32][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][29].cb_test                                      ;
                vSys2PeArray [32][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][30].cb_test                                      ;
                vSys2PeArray [32][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[32][31].cb_test                                      ;
                vSys2PeArray [32][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [32][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[33][0].cb_test                                      ;
                vSys2PeArray [33][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][1].cb_test                                      ;
                vSys2PeArray [33][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][2].cb_test                                      ;
                vSys2PeArray [33][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][3].cb_test                                      ;
                vSys2PeArray [33][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][4].cb_test                                      ;
                vSys2PeArray [33][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][5].cb_test                                      ;
                vSys2PeArray [33][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][6].cb_test                                      ;
                vSys2PeArray [33][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][7].cb_test                                      ;
                vSys2PeArray [33][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][8].cb_test                                      ;
                vSys2PeArray [33][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][9].cb_test                                      ;
                vSys2PeArray [33][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][10].cb_test                                      ;
                vSys2PeArray [33][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][11].cb_test                                      ;
                vSys2PeArray [33][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][12].cb_test                                      ;
                vSys2PeArray [33][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][13].cb_test                                      ;
                vSys2PeArray [33][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][14].cb_test                                      ;
                vSys2PeArray [33][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][15].cb_test                                      ;
                vSys2PeArray [33][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][16].cb_test                                      ;
                vSys2PeArray [33][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][17].cb_test                                      ;
                vSys2PeArray [33][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][18].cb_test                                      ;
                vSys2PeArray [33][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][19].cb_test                                      ;
                vSys2PeArray [33][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][20].cb_test                                      ;
                vSys2PeArray [33][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][21].cb_test                                      ;
                vSys2PeArray [33][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][22].cb_test                                      ;
                vSys2PeArray [33][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][23].cb_test                                      ;
                vSys2PeArray [33][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][24].cb_test                                      ;
                vSys2PeArray [33][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][25].cb_test                                      ;
                vSys2PeArray [33][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][26].cb_test                                      ;
                vSys2PeArray [33][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][27].cb_test                                      ;
                vSys2PeArray [33][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][28].cb_test                                      ;
                vSys2PeArray [33][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][29].cb_test                                      ;
                vSys2PeArray [33][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][30].cb_test                                      ;
                vSys2PeArray [33][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[33][31].cb_test                                      ;
                vSys2PeArray [33][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [33][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[34][0].cb_test                                      ;
                vSys2PeArray [34][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][1].cb_test                                      ;
                vSys2PeArray [34][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][2].cb_test                                      ;
                vSys2PeArray [34][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][3].cb_test                                      ;
                vSys2PeArray [34][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][4].cb_test                                      ;
                vSys2PeArray [34][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][5].cb_test                                      ;
                vSys2PeArray [34][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][6].cb_test                                      ;
                vSys2PeArray [34][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][7].cb_test                                      ;
                vSys2PeArray [34][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][8].cb_test                                      ;
                vSys2PeArray [34][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][9].cb_test                                      ;
                vSys2PeArray [34][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][10].cb_test                                      ;
                vSys2PeArray [34][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][11].cb_test                                      ;
                vSys2PeArray [34][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][12].cb_test                                      ;
                vSys2PeArray [34][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][13].cb_test                                      ;
                vSys2PeArray [34][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][14].cb_test                                      ;
                vSys2PeArray [34][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][15].cb_test                                      ;
                vSys2PeArray [34][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][16].cb_test                                      ;
                vSys2PeArray [34][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][17].cb_test                                      ;
                vSys2PeArray [34][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][18].cb_test                                      ;
                vSys2PeArray [34][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][19].cb_test                                      ;
                vSys2PeArray [34][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][20].cb_test                                      ;
                vSys2PeArray [34][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][21].cb_test                                      ;
                vSys2PeArray [34][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][22].cb_test                                      ;
                vSys2PeArray [34][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][23].cb_test                                      ;
                vSys2PeArray [34][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][24].cb_test                                      ;
                vSys2PeArray [34][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][25].cb_test                                      ;
                vSys2PeArray [34][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][26].cb_test                                      ;
                vSys2PeArray [34][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][27].cb_test                                      ;
                vSys2PeArray [34][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][28].cb_test                                      ;
                vSys2PeArray [34][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][29].cb_test                                      ;
                vSys2PeArray [34][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][30].cb_test                                      ;
                vSys2PeArray [34][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[34][31].cb_test                                      ;
                vSys2PeArray [34][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [34][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[35][0].cb_test                                      ;
                vSys2PeArray [35][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][1].cb_test                                      ;
                vSys2PeArray [35][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][2].cb_test                                      ;
                vSys2PeArray [35][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][3].cb_test                                      ;
                vSys2PeArray [35][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][4].cb_test                                      ;
                vSys2PeArray [35][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][5].cb_test                                      ;
                vSys2PeArray [35][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][6].cb_test                                      ;
                vSys2PeArray [35][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][7].cb_test                                      ;
                vSys2PeArray [35][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][8].cb_test                                      ;
                vSys2PeArray [35][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][9].cb_test                                      ;
                vSys2PeArray [35][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][10].cb_test                                      ;
                vSys2PeArray [35][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][11].cb_test                                      ;
                vSys2PeArray [35][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][12].cb_test                                      ;
                vSys2PeArray [35][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][13].cb_test                                      ;
                vSys2PeArray [35][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][14].cb_test                                      ;
                vSys2PeArray [35][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][15].cb_test                                      ;
                vSys2PeArray [35][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][16].cb_test                                      ;
                vSys2PeArray [35][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][17].cb_test                                      ;
                vSys2PeArray [35][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][18].cb_test                                      ;
                vSys2PeArray [35][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][19].cb_test                                      ;
                vSys2PeArray [35][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][20].cb_test                                      ;
                vSys2PeArray [35][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][21].cb_test                                      ;
                vSys2PeArray [35][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][22].cb_test                                      ;
                vSys2PeArray [35][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][23].cb_test                                      ;
                vSys2PeArray [35][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][24].cb_test                                      ;
                vSys2PeArray [35][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][25].cb_test                                      ;
                vSys2PeArray [35][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][26].cb_test                                      ;
                vSys2PeArray [35][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][27].cb_test                                      ;
                vSys2PeArray [35][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][28].cb_test                                      ;
                vSys2PeArray [35][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][29].cb_test                                      ;
                vSys2PeArray [35][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][30].cb_test                                      ;
                vSys2PeArray [35][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[35][31].cb_test                                      ;
                vSys2PeArray [35][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [35][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[36][0].cb_test                                      ;
                vSys2PeArray [36][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][1].cb_test                                      ;
                vSys2PeArray [36][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][2].cb_test                                      ;
                vSys2PeArray [36][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][3].cb_test                                      ;
                vSys2PeArray [36][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][4].cb_test                                      ;
                vSys2PeArray [36][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][5].cb_test                                      ;
                vSys2PeArray [36][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][6].cb_test                                      ;
                vSys2PeArray [36][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][7].cb_test                                      ;
                vSys2PeArray [36][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][8].cb_test                                      ;
                vSys2PeArray [36][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][9].cb_test                                      ;
                vSys2PeArray [36][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][10].cb_test                                      ;
                vSys2PeArray [36][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][11].cb_test                                      ;
                vSys2PeArray [36][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][12].cb_test                                      ;
                vSys2PeArray [36][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][13].cb_test                                      ;
                vSys2PeArray [36][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][14].cb_test                                      ;
                vSys2PeArray [36][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][15].cb_test                                      ;
                vSys2PeArray [36][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][16].cb_test                                      ;
                vSys2PeArray [36][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][17].cb_test                                      ;
                vSys2PeArray [36][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][18].cb_test                                      ;
                vSys2PeArray [36][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][19].cb_test                                      ;
                vSys2PeArray [36][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][20].cb_test                                      ;
                vSys2PeArray [36][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][21].cb_test                                      ;
                vSys2PeArray [36][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][22].cb_test                                      ;
                vSys2PeArray [36][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][23].cb_test                                      ;
                vSys2PeArray [36][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][24].cb_test                                      ;
                vSys2PeArray [36][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][25].cb_test                                      ;
                vSys2PeArray [36][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][26].cb_test                                      ;
                vSys2PeArray [36][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][27].cb_test                                      ;
                vSys2PeArray [36][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][28].cb_test                                      ;
                vSys2PeArray [36][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][29].cb_test                                      ;
                vSys2PeArray [36][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][30].cb_test                                      ;
                vSys2PeArray [36][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[36][31].cb_test                                      ;
                vSys2PeArray [36][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [36][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[37][0].cb_test                                      ;
                vSys2PeArray [37][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][1].cb_test                                      ;
                vSys2PeArray [37][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][2].cb_test                                      ;
                vSys2PeArray [37][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][3].cb_test                                      ;
                vSys2PeArray [37][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][4].cb_test                                      ;
                vSys2PeArray [37][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][5].cb_test                                      ;
                vSys2PeArray [37][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][6].cb_test                                      ;
                vSys2PeArray [37][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][7].cb_test                                      ;
                vSys2PeArray [37][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][8].cb_test                                      ;
                vSys2PeArray [37][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][9].cb_test                                      ;
                vSys2PeArray [37][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][10].cb_test                                      ;
                vSys2PeArray [37][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][11].cb_test                                      ;
                vSys2PeArray [37][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][12].cb_test                                      ;
                vSys2PeArray [37][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][13].cb_test                                      ;
                vSys2PeArray [37][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][14].cb_test                                      ;
                vSys2PeArray [37][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][15].cb_test                                      ;
                vSys2PeArray [37][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][16].cb_test                                      ;
                vSys2PeArray [37][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][17].cb_test                                      ;
                vSys2PeArray [37][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][18].cb_test                                      ;
                vSys2PeArray [37][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][19].cb_test                                      ;
                vSys2PeArray [37][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][20].cb_test                                      ;
                vSys2PeArray [37][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][21].cb_test                                      ;
                vSys2PeArray [37][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][22].cb_test                                      ;
                vSys2PeArray [37][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][23].cb_test                                      ;
                vSys2PeArray [37][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][24].cb_test                                      ;
                vSys2PeArray [37][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][25].cb_test                                      ;
                vSys2PeArray [37][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][26].cb_test                                      ;
                vSys2PeArray [37][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][27].cb_test                                      ;
                vSys2PeArray [37][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][28].cb_test                                      ;
                vSys2PeArray [37][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][29].cb_test                                      ;
                vSys2PeArray [37][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][30].cb_test                                      ;
                vSys2PeArray [37][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[37][31].cb_test                                      ;
                vSys2PeArray [37][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [37][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[38][0].cb_test                                      ;
                vSys2PeArray [38][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][1].cb_test                                      ;
                vSys2PeArray [38][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][2].cb_test                                      ;
                vSys2PeArray [38][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][3].cb_test                                      ;
                vSys2PeArray [38][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][4].cb_test                                      ;
                vSys2PeArray [38][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][5].cb_test                                      ;
                vSys2PeArray [38][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][6].cb_test                                      ;
                vSys2PeArray [38][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][7].cb_test                                      ;
                vSys2PeArray [38][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][8].cb_test                                      ;
                vSys2PeArray [38][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][9].cb_test                                      ;
                vSys2PeArray [38][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][10].cb_test                                      ;
                vSys2PeArray [38][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][11].cb_test                                      ;
                vSys2PeArray [38][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][12].cb_test                                      ;
                vSys2PeArray [38][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][13].cb_test                                      ;
                vSys2PeArray [38][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][14].cb_test                                      ;
                vSys2PeArray [38][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][15].cb_test                                      ;
                vSys2PeArray [38][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][16].cb_test                                      ;
                vSys2PeArray [38][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][17].cb_test                                      ;
                vSys2PeArray [38][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][18].cb_test                                      ;
                vSys2PeArray [38][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][19].cb_test                                      ;
                vSys2PeArray [38][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][20].cb_test                                      ;
                vSys2PeArray [38][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][21].cb_test                                      ;
                vSys2PeArray [38][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][22].cb_test                                      ;
                vSys2PeArray [38][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][23].cb_test                                      ;
                vSys2PeArray [38][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][24].cb_test                                      ;
                vSys2PeArray [38][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][25].cb_test                                      ;
                vSys2PeArray [38][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][26].cb_test                                      ;
                vSys2PeArray [38][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][27].cb_test                                      ;
                vSys2PeArray [38][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][28].cb_test                                      ;
                vSys2PeArray [38][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][29].cb_test                                      ;
                vSys2PeArray [38][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][30].cb_test                                      ;
                vSys2PeArray [38][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[38][31].cb_test                                      ;
                vSys2PeArray [38][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [38][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[39][0].cb_test                                      ;
                vSys2PeArray [39][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][1].cb_test                                      ;
                vSys2PeArray [39][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][2].cb_test                                      ;
                vSys2PeArray [39][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][3].cb_test                                      ;
                vSys2PeArray [39][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][4].cb_test                                      ;
                vSys2PeArray [39][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][5].cb_test                                      ;
                vSys2PeArray [39][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][6].cb_test                                      ;
                vSys2PeArray [39][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][7].cb_test                                      ;
                vSys2PeArray [39][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][8].cb_test                                      ;
                vSys2PeArray [39][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][9].cb_test                                      ;
                vSys2PeArray [39][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][10].cb_test                                      ;
                vSys2PeArray [39][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][11].cb_test                                      ;
                vSys2PeArray [39][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][12].cb_test                                      ;
                vSys2PeArray [39][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][13].cb_test                                      ;
                vSys2PeArray [39][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][14].cb_test                                      ;
                vSys2PeArray [39][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][15].cb_test                                      ;
                vSys2PeArray [39][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][16].cb_test                                      ;
                vSys2PeArray [39][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][17].cb_test                                      ;
                vSys2PeArray [39][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][18].cb_test                                      ;
                vSys2PeArray [39][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][19].cb_test                                      ;
                vSys2PeArray [39][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][20].cb_test                                      ;
                vSys2PeArray [39][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][21].cb_test                                      ;
                vSys2PeArray [39][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][22].cb_test                                      ;
                vSys2PeArray [39][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][23].cb_test                                      ;
                vSys2PeArray [39][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][24].cb_test                                      ;
                vSys2PeArray [39][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][25].cb_test                                      ;
                vSys2PeArray [39][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][26].cb_test                                      ;
                vSys2PeArray [39][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][27].cb_test                                      ;
                vSys2PeArray [39][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][28].cb_test                                      ;
                vSys2PeArray [39][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][29].cb_test                                      ;
                vSys2PeArray [39][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][30].cb_test                                      ;
                vSys2PeArray [39][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[39][31].cb_test                                      ;
                vSys2PeArray [39][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [39][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[40][0].cb_test                                      ;
                vSys2PeArray [40][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][1].cb_test                                      ;
                vSys2PeArray [40][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][2].cb_test                                      ;
                vSys2PeArray [40][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][3].cb_test                                      ;
                vSys2PeArray [40][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][4].cb_test                                      ;
                vSys2PeArray [40][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][5].cb_test                                      ;
                vSys2PeArray [40][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][6].cb_test                                      ;
                vSys2PeArray [40][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][7].cb_test                                      ;
                vSys2PeArray [40][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][8].cb_test                                      ;
                vSys2PeArray [40][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][9].cb_test                                      ;
                vSys2PeArray [40][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][10].cb_test                                      ;
                vSys2PeArray [40][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][11].cb_test                                      ;
                vSys2PeArray [40][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][12].cb_test                                      ;
                vSys2PeArray [40][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][13].cb_test                                      ;
                vSys2PeArray [40][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][14].cb_test                                      ;
                vSys2PeArray [40][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][15].cb_test                                      ;
                vSys2PeArray [40][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][16].cb_test                                      ;
                vSys2PeArray [40][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][17].cb_test                                      ;
                vSys2PeArray [40][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][18].cb_test                                      ;
                vSys2PeArray [40][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][19].cb_test                                      ;
                vSys2PeArray [40][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][20].cb_test                                      ;
                vSys2PeArray [40][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][21].cb_test                                      ;
                vSys2PeArray [40][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][22].cb_test                                      ;
                vSys2PeArray [40][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][23].cb_test                                      ;
                vSys2PeArray [40][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][24].cb_test                                      ;
                vSys2PeArray [40][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][25].cb_test                                      ;
                vSys2PeArray [40][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][26].cb_test                                      ;
                vSys2PeArray [40][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][27].cb_test                                      ;
                vSys2PeArray [40][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][28].cb_test                                      ;
                vSys2PeArray [40][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][29].cb_test                                      ;
                vSys2PeArray [40][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][30].cb_test                                      ;
                vSys2PeArray [40][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[40][31].cb_test                                      ;
                vSys2PeArray [40][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [40][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[41][0].cb_test                                      ;
                vSys2PeArray [41][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][1].cb_test                                      ;
                vSys2PeArray [41][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][2].cb_test                                      ;
                vSys2PeArray [41][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][3].cb_test                                      ;
                vSys2PeArray [41][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][4].cb_test                                      ;
                vSys2PeArray [41][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][5].cb_test                                      ;
                vSys2PeArray [41][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][6].cb_test                                      ;
                vSys2PeArray [41][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][7].cb_test                                      ;
                vSys2PeArray [41][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][8].cb_test                                      ;
                vSys2PeArray [41][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][9].cb_test                                      ;
                vSys2PeArray [41][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][10].cb_test                                      ;
                vSys2PeArray [41][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][11].cb_test                                      ;
                vSys2PeArray [41][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][12].cb_test                                      ;
                vSys2PeArray [41][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][13].cb_test                                      ;
                vSys2PeArray [41][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][14].cb_test                                      ;
                vSys2PeArray [41][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][15].cb_test                                      ;
                vSys2PeArray [41][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][16].cb_test                                      ;
                vSys2PeArray [41][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][17].cb_test                                      ;
                vSys2PeArray [41][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][18].cb_test                                      ;
                vSys2PeArray [41][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][19].cb_test                                      ;
                vSys2PeArray [41][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][20].cb_test                                      ;
                vSys2PeArray [41][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][21].cb_test                                      ;
                vSys2PeArray [41][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][22].cb_test                                      ;
                vSys2PeArray [41][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][23].cb_test                                      ;
                vSys2PeArray [41][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][24].cb_test                                      ;
                vSys2PeArray [41][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][25].cb_test                                      ;
                vSys2PeArray [41][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][26].cb_test                                      ;
                vSys2PeArray [41][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][27].cb_test                                      ;
                vSys2PeArray [41][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][28].cb_test                                      ;
                vSys2PeArray [41][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][29].cb_test                                      ;
                vSys2PeArray [41][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][30].cb_test                                      ;
                vSys2PeArray [41][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[41][31].cb_test                                      ;
                vSys2PeArray [41][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [41][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[42][0].cb_test                                      ;
                vSys2PeArray [42][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][1].cb_test                                      ;
                vSys2PeArray [42][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][2].cb_test                                      ;
                vSys2PeArray [42][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][3].cb_test                                      ;
                vSys2PeArray [42][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][4].cb_test                                      ;
                vSys2PeArray [42][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][5].cb_test                                      ;
                vSys2PeArray [42][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][6].cb_test                                      ;
                vSys2PeArray [42][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][7].cb_test                                      ;
                vSys2PeArray [42][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][8].cb_test                                      ;
                vSys2PeArray [42][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][9].cb_test                                      ;
                vSys2PeArray [42][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][10].cb_test                                      ;
                vSys2PeArray [42][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][11].cb_test                                      ;
                vSys2PeArray [42][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][12].cb_test                                      ;
                vSys2PeArray [42][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][13].cb_test                                      ;
                vSys2PeArray [42][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][14].cb_test                                      ;
                vSys2PeArray [42][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][15].cb_test                                      ;
                vSys2PeArray [42][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][16].cb_test                                      ;
                vSys2PeArray [42][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][17].cb_test                                      ;
                vSys2PeArray [42][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][18].cb_test                                      ;
                vSys2PeArray [42][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][19].cb_test                                      ;
                vSys2PeArray [42][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][20].cb_test                                      ;
                vSys2PeArray [42][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][21].cb_test                                      ;
                vSys2PeArray [42][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][22].cb_test                                      ;
                vSys2PeArray [42][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][23].cb_test                                      ;
                vSys2PeArray [42][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][24].cb_test                                      ;
                vSys2PeArray [42][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][25].cb_test                                      ;
                vSys2PeArray [42][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][26].cb_test                                      ;
                vSys2PeArray [42][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][27].cb_test                                      ;
                vSys2PeArray [42][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][28].cb_test                                      ;
                vSys2PeArray [42][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][29].cb_test                                      ;
                vSys2PeArray [42][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][30].cb_test                                      ;
                vSys2PeArray [42][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[42][31].cb_test                                      ;
                vSys2PeArray [42][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [42][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[43][0].cb_test                                      ;
                vSys2PeArray [43][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][1].cb_test                                      ;
                vSys2PeArray [43][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][2].cb_test                                      ;
                vSys2PeArray [43][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][3].cb_test                                      ;
                vSys2PeArray [43][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][4].cb_test                                      ;
                vSys2PeArray [43][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][5].cb_test                                      ;
                vSys2PeArray [43][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][6].cb_test                                      ;
                vSys2PeArray [43][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][7].cb_test                                      ;
                vSys2PeArray [43][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][8].cb_test                                      ;
                vSys2PeArray [43][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][9].cb_test                                      ;
                vSys2PeArray [43][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][10].cb_test                                      ;
                vSys2PeArray [43][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][11].cb_test                                      ;
                vSys2PeArray [43][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][12].cb_test                                      ;
                vSys2PeArray [43][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][13].cb_test                                      ;
                vSys2PeArray [43][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][14].cb_test                                      ;
                vSys2PeArray [43][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][15].cb_test                                      ;
                vSys2PeArray [43][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][16].cb_test                                      ;
                vSys2PeArray [43][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][17].cb_test                                      ;
                vSys2PeArray [43][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][18].cb_test                                      ;
                vSys2PeArray [43][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][19].cb_test                                      ;
                vSys2PeArray [43][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][20].cb_test                                      ;
                vSys2PeArray [43][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][21].cb_test                                      ;
                vSys2PeArray [43][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][22].cb_test                                      ;
                vSys2PeArray [43][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][23].cb_test                                      ;
                vSys2PeArray [43][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][24].cb_test                                      ;
                vSys2PeArray [43][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][25].cb_test                                      ;
                vSys2PeArray [43][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][26].cb_test                                      ;
                vSys2PeArray [43][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][27].cb_test                                      ;
                vSys2PeArray [43][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][28].cb_test                                      ;
                vSys2PeArray [43][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][29].cb_test                                      ;
                vSys2PeArray [43][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][30].cb_test                                      ;
                vSys2PeArray [43][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[43][31].cb_test                                      ;
                vSys2PeArray [43][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [43][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[44][0].cb_test                                      ;
                vSys2PeArray [44][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][1].cb_test                                      ;
                vSys2PeArray [44][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][2].cb_test                                      ;
                vSys2PeArray [44][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][3].cb_test                                      ;
                vSys2PeArray [44][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][4].cb_test                                      ;
                vSys2PeArray [44][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][5].cb_test                                      ;
                vSys2PeArray [44][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][6].cb_test                                      ;
                vSys2PeArray [44][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][7].cb_test                                      ;
                vSys2PeArray [44][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][8].cb_test                                      ;
                vSys2PeArray [44][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][9].cb_test                                      ;
                vSys2PeArray [44][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][10].cb_test                                      ;
                vSys2PeArray [44][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][11].cb_test                                      ;
                vSys2PeArray [44][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][12].cb_test                                      ;
                vSys2PeArray [44][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][13].cb_test                                      ;
                vSys2PeArray [44][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][14].cb_test                                      ;
                vSys2PeArray [44][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][15].cb_test                                      ;
                vSys2PeArray [44][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][16].cb_test                                      ;
                vSys2PeArray [44][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][17].cb_test                                      ;
                vSys2PeArray [44][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][18].cb_test                                      ;
                vSys2PeArray [44][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][19].cb_test                                      ;
                vSys2PeArray [44][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][20].cb_test                                      ;
                vSys2PeArray [44][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][21].cb_test                                      ;
                vSys2PeArray [44][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][22].cb_test                                      ;
                vSys2PeArray [44][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][23].cb_test                                      ;
                vSys2PeArray [44][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][24].cb_test                                      ;
                vSys2PeArray [44][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][25].cb_test                                      ;
                vSys2PeArray [44][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][26].cb_test                                      ;
                vSys2PeArray [44][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][27].cb_test                                      ;
                vSys2PeArray [44][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][28].cb_test                                      ;
                vSys2PeArray [44][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][29].cb_test                                      ;
                vSys2PeArray [44][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][30].cb_test                                      ;
                vSys2PeArray [44][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[44][31].cb_test                                      ;
                vSys2PeArray [44][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [44][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[45][0].cb_test                                      ;
                vSys2PeArray [45][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][1].cb_test                                      ;
                vSys2PeArray [45][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][2].cb_test                                      ;
                vSys2PeArray [45][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][3].cb_test                                      ;
                vSys2PeArray [45][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][4].cb_test                                      ;
                vSys2PeArray [45][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][5].cb_test                                      ;
                vSys2PeArray [45][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][6].cb_test                                      ;
                vSys2PeArray [45][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][7].cb_test                                      ;
                vSys2PeArray [45][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][8].cb_test                                      ;
                vSys2PeArray [45][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][9].cb_test                                      ;
                vSys2PeArray [45][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][10].cb_test                                      ;
                vSys2PeArray [45][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][11].cb_test                                      ;
                vSys2PeArray [45][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][12].cb_test                                      ;
                vSys2PeArray [45][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][13].cb_test                                      ;
                vSys2PeArray [45][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][14].cb_test                                      ;
                vSys2PeArray [45][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][15].cb_test                                      ;
                vSys2PeArray [45][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][16].cb_test                                      ;
                vSys2PeArray [45][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][17].cb_test                                      ;
                vSys2PeArray [45][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][18].cb_test                                      ;
                vSys2PeArray [45][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][19].cb_test                                      ;
                vSys2PeArray [45][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][20].cb_test                                      ;
                vSys2PeArray [45][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][21].cb_test                                      ;
                vSys2PeArray [45][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][22].cb_test                                      ;
                vSys2PeArray [45][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][23].cb_test                                      ;
                vSys2PeArray [45][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][24].cb_test                                      ;
                vSys2PeArray [45][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][25].cb_test                                      ;
                vSys2PeArray [45][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][26].cb_test                                      ;
                vSys2PeArray [45][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][27].cb_test                                      ;
                vSys2PeArray [45][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][28].cb_test                                      ;
                vSys2PeArray [45][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][29].cb_test                                      ;
                vSys2PeArray [45][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][30].cb_test                                      ;
                vSys2PeArray [45][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[45][31].cb_test                                      ;
                vSys2PeArray [45][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [45][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[46][0].cb_test                                      ;
                vSys2PeArray [46][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][1].cb_test                                      ;
                vSys2PeArray [46][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][2].cb_test                                      ;
                vSys2PeArray [46][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][3].cb_test                                      ;
                vSys2PeArray [46][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][4].cb_test                                      ;
                vSys2PeArray [46][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][5].cb_test                                      ;
                vSys2PeArray [46][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][6].cb_test                                      ;
                vSys2PeArray [46][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][7].cb_test                                      ;
                vSys2PeArray [46][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][8].cb_test                                      ;
                vSys2PeArray [46][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][9].cb_test                                      ;
                vSys2PeArray [46][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][10].cb_test                                      ;
                vSys2PeArray [46][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][11].cb_test                                      ;
                vSys2PeArray [46][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][12].cb_test                                      ;
                vSys2PeArray [46][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][13].cb_test                                      ;
                vSys2PeArray [46][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][14].cb_test                                      ;
                vSys2PeArray [46][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][15].cb_test                                      ;
                vSys2PeArray [46][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][16].cb_test                                      ;
                vSys2PeArray [46][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][17].cb_test                                      ;
                vSys2PeArray [46][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][18].cb_test                                      ;
                vSys2PeArray [46][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][19].cb_test                                      ;
                vSys2PeArray [46][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][20].cb_test                                      ;
                vSys2PeArray [46][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][21].cb_test                                      ;
                vSys2PeArray [46][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][22].cb_test                                      ;
                vSys2PeArray [46][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][23].cb_test                                      ;
                vSys2PeArray [46][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][24].cb_test                                      ;
                vSys2PeArray [46][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][25].cb_test                                      ;
                vSys2PeArray [46][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][26].cb_test                                      ;
                vSys2PeArray [46][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][27].cb_test                                      ;
                vSys2PeArray [46][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][28].cb_test                                      ;
                vSys2PeArray [46][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][29].cb_test                                      ;
                vSys2PeArray [46][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][30].cb_test                                      ;
                vSys2PeArray [46][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[46][31].cb_test                                      ;
                vSys2PeArray [46][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [46][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[47][0].cb_test                                      ;
                vSys2PeArray [47][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][1].cb_test                                      ;
                vSys2PeArray [47][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][2].cb_test                                      ;
                vSys2PeArray [47][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][3].cb_test                                      ;
                vSys2PeArray [47][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][4].cb_test                                      ;
                vSys2PeArray [47][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][5].cb_test                                      ;
                vSys2PeArray [47][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][6].cb_test                                      ;
                vSys2PeArray [47][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][7].cb_test                                      ;
                vSys2PeArray [47][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][8].cb_test                                      ;
                vSys2PeArray [47][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][9].cb_test                                      ;
                vSys2PeArray [47][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][10].cb_test                                      ;
                vSys2PeArray [47][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][11].cb_test                                      ;
                vSys2PeArray [47][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][12].cb_test                                      ;
                vSys2PeArray [47][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][13].cb_test                                      ;
                vSys2PeArray [47][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][14].cb_test                                      ;
                vSys2PeArray [47][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][15].cb_test                                      ;
                vSys2PeArray [47][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][16].cb_test                                      ;
                vSys2PeArray [47][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][17].cb_test                                      ;
                vSys2PeArray [47][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][18].cb_test                                      ;
                vSys2PeArray [47][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][19].cb_test                                      ;
                vSys2PeArray [47][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][20].cb_test                                      ;
                vSys2PeArray [47][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][21].cb_test                                      ;
                vSys2PeArray [47][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][22].cb_test                                      ;
                vSys2PeArray [47][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][23].cb_test                                      ;
                vSys2PeArray [47][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][24].cb_test                                      ;
                vSys2PeArray [47][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][25].cb_test                                      ;
                vSys2PeArray [47][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][26].cb_test                                      ;
                vSys2PeArray [47][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][27].cb_test                                      ;
                vSys2PeArray [47][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][28].cb_test                                      ;
                vSys2PeArray [47][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][29].cb_test                                      ;
                vSys2PeArray [47][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][30].cb_test                                      ;
                vSys2PeArray [47][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[47][31].cb_test                                      ;
                vSys2PeArray [47][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [47][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[48][0].cb_test                                      ;
                vSys2PeArray [48][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][1].cb_test                                      ;
                vSys2PeArray [48][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][2].cb_test                                      ;
                vSys2PeArray [48][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][3].cb_test                                      ;
                vSys2PeArray [48][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][4].cb_test                                      ;
                vSys2PeArray [48][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][5].cb_test                                      ;
                vSys2PeArray [48][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][6].cb_test                                      ;
                vSys2PeArray [48][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][7].cb_test                                      ;
                vSys2PeArray [48][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][8].cb_test                                      ;
                vSys2PeArray [48][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][9].cb_test                                      ;
                vSys2PeArray [48][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][10].cb_test                                      ;
                vSys2PeArray [48][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][11].cb_test                                      ;
                vSys2PeArray [48][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][12].cb_test                                      ;
                vSys2PeArray [48][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][13].cb_test                                      ;
                vSys2PeArray [48][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][14].cb_test                                      ;
                vSys2PeArray [48][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][15].cb_test                                      ;
                vSys2PeArray [48][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][16].cb_test                                      ;
                vSys2PeArray [48][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][17].cb_test                                      ;
                vSys2PeArray [48][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][18].cb_test                                      ;
                vSys2PeArray [48][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][19].cb_test                                      ;
                vSys2PeArray [48][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][20].cb_test                                      ;
                vSys2PeArray [48][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][21].cb_test                                      ;
                vSys2PeArray [48][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][22].cb_test                                      ;
                vSys2PeArray [48][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][23].cb_test                                      ;
                vSys2PeArray [48][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][24].cb_test                                      ;
                vSys2PeArray [48][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][25].cb_test                                      ;
                vSys2PeArray [48][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][26].cb_test                                      ;
                vSys2PeArray [48][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][27].cb_test                                      ;
                vSys2PeArray [48][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][28].cb_test                                      ;
                vSys2PeArray [48][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][29].cb_test                                      ;
                vSys2PeArray [48][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][30].cb_test                                      ;
                vSys2PeArray [48][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[48][31].cb_test                                      ;
                vSys2PeArray [48][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [48][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[49][0].cb_test                                      ;
                vSys2PeArray [49][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][1].cb_test                                      ;
                vSys2PeArray [49][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][2].cb_test                                      ;
                vSys2PeArray [49][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][3].cb_test                                      ;
                vSys2PeArray [49][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][4].cb_test                                      ;
                vSys2PeArray [49][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][5].cb_test                                      ;
                vSys2PeArray [49][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][6].cb_test                                      ;
                vSys2PeArray [49][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][7].cb_test                                      ;
                vSys2PeArray [49][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][8].cb_test                                      ;
                vSys2PeArray [49][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][9].cb_test                                      ;
                vSys2PeArray [49][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][10].cb_test                                      ;
                vSys2PeArray [49][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][11].cb_test                                      ;
                vSys2PeArray [49][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][12].cb_test                                      ;
                vSys2PeArray [49][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][13].cb_test                                      ;
                vSys2PeArray [49][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][14].cb_test                                      ;
                vSys2PeArray [49][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][15].cb_test                                      ;
                vSys2PeArray [49][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][16].cb_test                                      ;
                vSys2PeArray [49][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][17].cb_test                                      ;
                vSys2PeArray [49][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][18].cb_test                                      ;
                vSys2PeArray [49][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][19].cb_test                                      ;
                vSys2PeArray [49][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][20].cb_test                                      ;
                vSys2PeArray [49][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][21].cb_test                                      ;
                vSys2PeArray [49][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][22].cb_test                                      ;
                vSys2PeArray [49][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][23].cb_test                                      ;
                vSys2PeArray [49][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][24].cb_test                                      ;
                vSys2PeArray [49][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][25].cb_test                                      ;
                vSys2PeArray [49][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][26].cb_test                                      ;
                vSys2PeArray [49][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][27].cb_test                                      ;
                vSys2PeArray [49][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][28].cb_test                                      ;
                vSys2PeArray [49][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][29].cb_test                                      ;
                vSys2PeArray [49][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][30].cb_test                                      ;
                vSys2PeArray [49][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[49][31].cb_test                                      ;
                vSys2PeArray [49][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [49][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[50][0].cb_test                                      ;
                vSys2PeArray [50][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][1].cb_test                                      ;
                vSys2PeArray [50][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][2].cb_test                                      ;
                vSys2PeArray [50][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][3].cb_test                                      ;
                vSys2PeArray [50][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][4].cb_test                                      ;
                vSys2PeArray [50][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][5].cb_test                                      ;
                vSys2PeArray [50][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][6].cb_test                                      ;
                vSys2PeArray [50][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][7].cb_test                                      ;
                vSys2PeArray [50][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][8].cb_test                                      ;
                vSys2PeArray [50][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][9].cb_test                                      ;
                vSys2PeArray [50][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][10].cb_test                                      ;
                vSys2PeArray [50][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][11].cb_test                                      ;
                vSys2PeArray [50][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][12].cb_test                                      ;
                vSys2PeArray [50][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][13].cb_test                                      ;
                vSys2PeArray [50][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][14].cb_test                                      ;
                vSys2PeArray [50][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][15].cb_test                                      ;
                vSys2PeArray [50][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][16].cb_test                                      ;
                vSys2PeArray [50][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][17].cb_test                                      ;
                vSys2PeArray [50][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][18].cb_test                                      ;
                vSys2PeArray [50][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][19].cb_test                                      ;
                vSys2PeArray [50][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][20].cb_test                                      ;
                vSys2PeArray [50][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][21].cb_test                                      ;
                vSys2PeArray [50][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][22].cb_test                                      ;
                vSys2PeArray [50][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][23].cb_test                                      ;
                vSys2PeArray [50][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][24].cb_test                                      ;
                vSys2PeArray [50][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][25].cb_test                                      ;
                vSys2PeArray [50][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][26].cb_test                                      ;
                vSys2PeArray [50][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][27].cb_test                                      ;
                vSys2PeArray [50][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][28].cb_test                                      ;
                vSys2PeArray [50][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][29].cb_test                                      ;
                vSys2PeArray [50][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][30].cb_test                                      ;
                vSys2PeArray [50][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[50][31].cb_test                                      ;
                vSys2PeArray [50][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [50][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[51][0].cb_test                                      ;
                vSys2PeArray [51][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][1].cb_test                                      ;
                vSys2PeArray [51][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][2].cb_test                                      ;
                vSys2PeArray [51][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][3].cb_test                                      ;
                vSys2PeArray [51][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][4].cb_test                                      ;
                vSys2PeArray [51][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][5].cb_test                                      ;
                vSys2PeArray [51][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][6].cb_test                                      ;
                vSys2PeArray [51][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][7].cb_test                                      ;
                vSys2PeArray [51][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][8].cb_test                                      ;
                vSys2PeArray [51][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][9].cb_test                                      ;
                vSys2PeArray [51][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][10].cb_test                                      ;
                vSys2PeArray [51][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][11].cb_test                                      ;
                vSys2PeArray [51][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][12].cb_test                                      ;
                vSys2PeArray [51][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][13].cb_test                                      ;
                vSys2PeArray [51][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][14].cb_test                                      ;
                vSys2PeArray [51][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][15].cb_test                                      ;
                vSys2PeArray [51][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][16].cb_test                                      ;
                vSys2PeArray [51][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][17].cb_test                                      ;
                vSys2PeArray [51][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][18].cb_test                                      ;
                vSys2PeArray [51][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][19].cb_test                                      ;
                vSys2PeArray [51][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][20].cb_test                                      ;
                vSys2PeArray [51][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][21].cb_test                                      ;
                vSys2PeArray [51][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][22].cb_test                                      ;
                vSys2PeArray [51][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][23].cb_test                                      ;
                vSys2PeArray [51][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][24].cb_test                                      ;
                vSys2PeArray [51][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][25].cb_test                                      ;
                vSys2PeArray [51][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][26].cb_test                                      ;
                vSys2PeArray [51][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][27].cb_test                                      ;
                vSys2PeArray [51][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][28].cb_test                                      ;
                vSys2PeArray [51][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][29].cb_test                                      ;
                vSys2PeArray [51][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][30].cb_test                                      ;
                vSys2PeArray [51][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[51][31].cb_test                                      ;
                vSys2PeArray [51][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [51][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[52][0].cb_test                                      ;
                vSys2PeArray [52][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][1].cb_test                                      ;
                vSys2PeArray [52][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][2].cb_test                                      ;
                vSys2PeArray [52][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][3].cb_test                                      ;
                vSys2PeArray [52][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][4].cb_test                                      ;
                vSys2PeArray [52][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][5].cb_test                                      ;
                vSys2PeArray [52][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][6].cb_test                                      ;
                vSys2PeArray [52][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][7].cb_test                                      ;
                vSys2PeArray [52][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][8].cb_test                                      ;
                vSys2PeArray [52][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][9].cb_test                                      ;
                vSys2PeArray [52][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][10].cb_test                                      ;
                vSys2PeArray [52][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][11].cb_test                                      ;
                vSys2PeArray [52][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][12].cb_test                                      ;
                vSys2PeArray [52][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][13].cb_test                                      ;
                vSys2PeArray [52][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][14].cb_test                                      ;
                vSys2PeArray [52][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][15].cb_test                                      ;
                vSys2PeArray [52][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][16].cb_test                                      ;
                vSys2PeArray [52][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][17].cb_test                                      ;
                vSys2PeArray [52][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][18].cb_test                                      ;
                vSys2PeArray [52][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][19].cb_test                                      ;
                vSys2PeArray [52][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][20].cb_test                                      ;
                vSys2PeArray [52][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][21].cb_test                                      ;
                vSys2PeArray [52][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][22].cb_test                                      ;
                vSys2PeArray [52][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][23].cb_test                                      ;
                vSys2PeArray [52][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][24].cb_test                                      ;
                vSys2PeArray [52][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][25].cb_test                                      ;
                vSys2PeArray [52][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][26].cb_test                                      ;
                vSys2PeArray [52][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][27].cb_test                                      ;
                vSys2PeArray [52][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][28].cb_test                                      ;
                vSys2PeArray [52][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][29].cb_test                                      ;
                vSys2PeArray [52][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][30].cb_test                                      ;
                vSys2PeArray [52][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[52][31].cb_test                                      ;
                vSys2PeArray [52][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [52][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[53][0].cb_test                                      ;
                vSys2PeArray [53][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][1].cb_test                                      ;
                vSys2PeArray [53][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][2].cb_test                                      ;
                vSys2PeArray [53][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][3].cb_test                                      ;
                vSys2PeArray [53][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][4].cb_test                                      ;
                vSys2PeArray [53][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][5].cb_test                                      ;
                vSys2PeArray [53][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][6].cb_test                                      ;
                vSys2PeArray [53][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][7].cb_test                                      ;
                vSys2PeArray [53][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][8].cb_test                                      ;
                vSys2PeArray [53][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][9].cb_test                                      ;
                vSys2PeArray [53][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][10].cb_test                                      ;
                vSys2PeArray [53][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][11].cb_test                                      ;
                vSys2PeArray [53][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][12].cb_test                                      ;
                vSys2PeArray [53][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][13].cb_test                                      ;
                vSys2PeArray [53][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][14].cb_test                                      ;
                vSys2PeArray [53][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][15].cb_test                                      ;
                vSys2PeArray [53][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][16].cb_test                                      ;
                vSys2PeArray [53][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][17].cb_test                                      ;
                vSys2PeArray [53][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][18].cb_test                                      ;
                vSys2PeArray [53][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][19].cb_test                                      ;
                vSys2PeArray [53][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][20].cb_test                                      ;
                vSys2PeArray [53][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][21].cb_test                                      ;
                vSys2PeArray [53][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][22].cb_test                                      ;
                vSys2PeArray [53][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][23].cb_test                                      ;
                vSys2PeArray [53][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][24].cb_test                                      ;
                vSys2PeArray [53][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][25].cb_test                                      ;
                vSys2PeArray [53][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][26].cb_test                                      ;
                vSys2PeArray [53][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][27].cb_test                                      ;
                vSys2PeArray [53][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][28].cb_test                                      ;
                vSys2PeArray [53][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][29].cb_test                                      ;
                vSys2PeArray [53][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][30].cb_test                                      ;
                vSys2PeArray [53][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[53][31].cb_test                                      ;
                vSys2PeArray [53][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [53][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[54][0].cb_test                                      ;
                vSys2PeArray [54][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][1].cb_test                                      ;
                vSys2PeArray [54][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][2].cb_test                                      ;
                vSys2PeArray [54][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][3].cb_test                                      ;
                vSys2PeArray [54][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][4].cb_test                                      ;
                vSys2PeArray [54][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][5].cb_test                                      ;
                vSys2PeArray [54][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][6].cb_test                                      ;
                vSys2PeArray [54][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][7].cb_test                                      ;
                vSys2PeArray [54][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][8].cb_test                                      ;
                vSys2PeArray [54][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][9].cb_test                                      ;
                vSys2PeArray [54][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][10].cb_test                                      ;
                vSys2PeArray [54][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][11].cb_test                                      ;
                vSys2PeArray [54][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][12].cb_test                                      ;
                vSys2PeArray [54][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][13].cb_test                                      ;
                vSys2PeArray [54][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][14].cb_test                                      ;
                vSys2PeArray [54][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][15].cb_test                                      ;
                vSys2PeArray [54][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][16].cb_test                                      ;
                vSys2PeArray [54][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][17].cb_test                                      ;
                vSys2PeArray [54][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][18].cb_test                                      ;
                vSys2PeArray [54][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][19].cb_test                                      ;
                vSys2PeArray [54][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][20].cb_test                                      ;
                vSys2PeArray [54][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][21].cb_test                                      ;
                vSys2PeArray [54][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][22].cb_test                                      ;
                vSys2PeArray [54][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][23].cb_test                                      ;
                vSys2PeArray [54][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][24].cb_test                                      ;
                vSys2PeArray [54][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][25].cb_test                                      ;
                vSys2PeArray [54][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][26].cb_test                                      ;
                vSys2PeArray [54][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][27].cb_test                                      ;
                vSys2PeArray [54][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][28].cb_test                                      ;
                vSys2PeArray [54][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][29].cb_test                                      ;
                vSys2PeArray [54][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][30].cb_test                                      ;
                vSys2PeArray [54][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[54][31].cb_test                                      ;
                vSys2PeArray [54][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [54][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[55][0].cb_test                                      ;
                vSys2PeArray [55][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][1].cb_test                                      ;
                vSys2PeArray [55][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][2].cb_test                                      ;
                vSys2PeArray [55][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][3].cb_test                                      ;
                vSys2PeArray [55][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][4].cb_test                                      ;
                vSys2PeArray [55][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][5].cb_test                                      ;
                vSys2PeArray [55][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][6].cb_test                                      ;
                vSys2PeArray [55][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][7].cb_test                                      ;
                vSys2PeArray [55][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][8].cb_test                                      ;
                vSys2PeArray [55][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][9].cb_test                                      ;
                vSys2PeArray [55][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][10].cb_test                                      ;
                vSys2PeArray [55][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][11].cb_test                                      ;
                vSys2PeArray [55][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][12].cb_test                                      ;
                vSys2PeArray [55][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][13].cb_test                                      ;
                vSys2PeArray [55][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][14].cb_test                                      ;
                vSys2PeArray [55][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][15].cb_test                                      ;
                vSys2PeArray [55][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][16].cb_test                                      ;
                vSys2PeArray [55][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][17].cb_test                                      ;
                vSys2PeArray [55][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][18].cb_test                                      ;
                vSys2PeArray [55][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][19].cb_test                                      ;
                vSys2PeArray [55][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][20].cb_test                                      ;
                vSys2PeArray [55][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][21].cb_test                                      ;
                vSys2PeArray [55][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][22].cb_test                                      ;
                vSys2PeArray [55][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][23].cb_test                                      ;
                vSys2PeArray [55][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][24].cb_test                                      ;
                vSys2PeArray [55][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][25].cb_test                                      ;
                vSys2PeArray [55][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][26].cb_test                                      ;
                vSys2PeArray [55][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][27].cb_test                                      ;
                vSys2PeArray [55][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][28].cb_test                                      ;
                vSys2PeArray [55][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][29].cb_test                                      ;
                vSys2PeArray [55][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][30].cb_test                                      ;
                vSys2PeArray [55][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[55][31].cb_test                                      ;
                vSys2PeArray [55][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [55][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[56][0].cb_test                                      ;
                vSys2PeArray [56][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][1].cb_test                                      ;
                vSys2PeArray [56][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][2].cb_test                                      ;
                vSys2PeArray [56][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][3].cb_test                                      ;
                vSys2PeArray [56][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][4].cb_test                                      ;
                vSys2PeArray [56][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][5].cb_test                                      ;
                vSys2PeArray [56][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][6].cb_test                                      ;
                vSys2PeArray [56][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][7].cb_test                                      ;
                vSys2PeArray [56][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][8].cb_test                                      ;
                vSys2PeArray [56][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][9].cb_test                                      ;
                vSys2PeArray [56][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][10].cb_test                                      ;
                vSys2PeArray [56][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][11].cb_test                                      ;
                vSys2PeArray [56][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][12].cb_test                                      ;
                vSys2PeArray [56][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][13].cb_test                                      ;
                vSys2PeArray [56][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][14].cb_test                                      ;
                vSys2PeArray [56][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][15].cb_test                                      ;
                vSys2PeArray [56][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][16].cb_test                                      ;
                vSys2PeArray [56][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][17].cb_test                                      ;
                vSys2PeArray [56][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][18].cb_test                                      ;
                vSys2PeArray [56][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][19].cb_test                                      ;
                vSys2PeArray [56][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][20].cb_test                                      ;
                vSys2PeArray [56][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][21].cb_test                                      ;
                vSys2PeArray [56][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][22].cb_test                                      ;
                vSys2PeArray [56][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][23].cb_test                                      ;
                vSys2PeArray [56][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][24].cb_test                                      ;
                vSys2PeArray [56][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][25].cb_test                                      ;
                vSys2PeArray [56][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][26].cb_test                                      ;
                vSys2PeArray [56][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][27].cb_test                                      ;
                vSys2PeArray [56][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][28].cb_test                                      ;
                vSys2PeArray [56][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][29].cb_test                                      ;
                vSys2PeArray [56][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][30].cb_test                                      ;
                vSys2PeArray [56][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[56][31].cb_test                                      ;
                vSys2PeArray [56][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [56][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[57][0].cb_test                                      ;
                vSys2PeArray [57][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][1].cb_test                                      ;
                vSys2PeArray [57][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][2].cb_test                                      ;
                vSys2PeArray [57][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][3].cb_test                                      ;
                vSys2PeArray [57][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][4].cb_test                                      ;
                vSys2PeArray [57][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][5].cb_test                                      ;
                vSys2PeArray [57][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][6].cb_test                                      ;
                vSys2PeArray [57][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][7].cb_test                                      ;
                vSys2PeArray [57][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][8].cb_test                                      ;
                vSys2PeArray [57][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][9].cb_test                                      ;
                vSys2PeArray [57][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][10].cb_test                                      ;
                vSys2PeArray [57][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][11].cb_test                                      ;
                vSys2PeArray [57][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][12].cb_test                                      ;
                vSys2PeArray [57][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][13].cb_test                                      ;
                vSys2PeArray [57][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][14].cb_test                                      ;
                vSys2PeArray [57][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][15].cb_test                                      ;
                vSys2PeArray [57][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][16].cb_test                                      ;
                vSys2PeArray [57][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][17].cb_test                                      ;
                vSys2PeArray [57][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][18].cb_test                                      ;
                vSys2PeArray [57][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][19].cb_test                                      ;
                vSys2PeArray [57][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][20].cb_test                                      ;
                vSys2PeArray [57][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][21].cb_test                                      ;
                vSys2PeArray [57][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][22].cb_test                                      ;
                vSys2PeArray [57][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][23].cb_test                                      ;
                vSys2PeArray [57][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][24].cb_test                                      ;
                vSys2PeArray [57][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][25].cb_test                                      ;
                vSys2PeArray [57][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][26].cb_test                                      ;
                vSys2PeArray [57][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][27].cb_test                                      ;
                vSys2PeArray [57][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][28].cb_test                                      ;
                vSys2PeArray [57][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][29].cb_test                                      ;
                vSys2PeArray [57][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][30].cb_test                                      ;
                vSys2PeArray [57][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[57][31].cb_test                                      ;
                vSys2PeArray [57][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [57][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[58][0].cb_test                                      ;
                vSys2PeArray [58][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][1].cb_test                                      ;
                vSys2PeArray [58][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][2].cb_test                                      ;
                vSys2PeArray [58][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][3].cb_test                                      ;
                vSys2PeArray [58][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][4].cb_test                                      ;
                vSys2PeArray [58][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][5].cb_test                                      ;
                vSys2PeArray [58][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][6].cb_test                                      ;
                vSys2PeArray [58][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][7].cb_test                                      ;
                vSys2PeArray [58][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][8].cb_test                                      ;
                vSys2PeArray [58][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][9].cb_test                                      ;
                vSys2PeArray [58][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][10].cb_test                                      ;
                vSys2PeArray [58][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][11].cb_test                                      ;
                vSys2PeArray [58][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][12].cb_test                                      ;
                vSys2PeArray [58][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][13].cb_test                                      ;
                vSys2PeArray [58][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][14].cb_test                                      ;
                vSys2PeArray [58][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][15].cb_test                                      ;
                vSys2PeArray [58][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][16].cb_test                                      ;
                vSys2PeArray [58][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][17].cb_test                                      ;
                vSys2PeArray [58][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][18].cb_test                                      ;
                vSys2PeArray [58][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][19].cb_test                                      ;
                vSys2PeArray [58][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][20].cb_test                                      ;
                vSys2PeArray [58][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][21].cb_test                                      ;
                vSys2PeArray [58][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][22].cb_test                                      ;
                vSys2PeArray [58][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][23].cb_test                                      ;
                vSys2PeArray [58][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][24].cb_test                                      ;
                vSys2PeArray [58][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][25].cb_test                                      ;
                vSys2PeArray [58][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][26].cb_test                                      ;
                vSys2PeArray [58][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][27].cb_test                                      ;
                vSys2PeArray [58][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][28].cb_test                                      ;
                vSys2PeArray [58][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][29].cb_test                                      ;
                vSys2PeArray [58][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][30].cb_test                                      ;
                vSys2PeArray [58][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[58][31].cb_test                                      ;
                vSys2PeArray [58][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [58][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[59][0].cb_test                                      ;
                vSys2PeArray [59][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][1].cb_test                                      ;
                vSys2PeArray [59][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][2].cb_test                                      ;
                vSys2PeArray [59][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][3].cb_test                                      ;
                vSys2PeArray [59][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][4].cb_test                                      ;
                vSys2PeArray [59][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][5].cb_test                                      ;
                vSys2PeArray [59][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][6].cb_test                                      ;
                vSys2PeArray [59][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][7].cb_test                                      ;
                vSys2PeArray [59][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][8].cb_test                                      ;
                vSys2PeArray [59][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][9].cb_test                                      ;
                vSys2PeArray [59][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][10].cb_test                                      ;
                vSys2PeArray [59][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][11].cb_test                                      ;
                vSys2PeArray [59][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][12].cb_test                                      ;
                vSys2PeArray [59][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][13].cb_test                                      ;
                vSys2PeArray [59][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][14].cb_test                                      ;
                vSys2PeArray [59][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][15].cb_test                                      ;
                vSys2PeArray [59][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][16].cb_test                                      ;
                vSys2PeArray [59][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][17].cb_test                                      ;
                vSys2PeArray [59][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][18].cb_test                                      ;
                vSys2PeArray [59][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][19].cb_test                                      ;
                vSys2PeArray [59][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][20].cb_test                                      ;
                vSys2PeArray [59][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][21].cb_test                                      ;
                vSys2PeArray [59][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][22].cb_test                                      ;
                vSys2PeArray [59][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][23].cb_test                                      ;
                vSys2PeArray [59][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][24].cb_test                                      ;
                vSys2PeArray [59][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][25].cb_test                                      ;
                vSys2PeArray [59][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][26].cb_test                                      ;
                vSys2PeArray [59][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][27].cb_test                                      ;
                vSys2PeArray [59][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][28].cb_test                                      ;
                vSys2PeArray [59][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][29].cb_test                                      ;
                vSys2PeArray [59][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][30].cb_test                                      ;
                vSys2PeArray [59][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[59][31].cb_test                                      ;
                vSys2PeArray [59][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [59][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[60][0].cb_test                                      ;
                vSys2PeArray [60][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][1].cb_test                                      ;
                vSys2PeArray [60][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][2].cb_test                                      ;
                vSys2PeArray [60][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][3].cb_test                                      ;
                vSys2PeArray [60][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][4].cb_test                                      ;
                vSys2PeArray [60][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][5].cb_test                                      ;
                vSys2PeArray [60][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][6].cb_test                                      ;
                vSys2PeArray [60][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][7].cb_test                                      ;
                vSys2PeArray [60][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][8].cb_test                                      ;
                vSys2PeArray [60][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][9].cb_test                                      ;
                vSys2PeArray [60][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][10].cb_test                                      ;
                vSys2PeArray [60][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][11].cb_test                                      ;
                vSys2PeArray [60][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][12].cb_test                                      ;
                vSys2PeArray [60][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][13].cb_test                                      ;
                vSys2PeArray [60][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][14].cb_test                                      ;
                vSys2PeArray [60][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][15].cb_test                                      ;
                vSys2PeArray [60][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][16].cb_test                                      ;
                vSys2PeArray [60][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][17].cb_test                                      ;
                vSys2PeArray [60][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][18].cb_test                                      ;
                vSys2PeArray [60][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][19].cb_test                                      ;
                vSys2PeArray [60][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][20].cb_test                                      ;
                vSys2PeArray [60][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][21].cb_test                                      ;
                vSys2PeArray [60][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][22].cb_test                                      ;
                vSys2PeArray [60][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][23].cb_test                                      ;
                vSys2PeArray [60][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][24].cb_test                                      ;
                vSys2PeArray [60][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][25].cb_test                                      ;
                vSys2PeArray [60][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][26].cb_test                                      ;
                vSys2PeArray [60][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][27].cb_test                                      ;
                vSys2PeArray [60][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][28].cb_test                                      ;
                vSys2PeArray [60][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][29].cb_test                                      ;
                vSys2PeArray [60][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][30].cb_test                                      ;
                vSys2PeArray [60][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[60][31].cb_test                                      ;
                vSys2PeArray [60][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [60][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[61][0].cb_test                                      ;
                vSys2PeArray [61][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][1].cb_test                                      ;
                vSys2PeArray [61][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][2].cb_test                                      ;
                vSys2PeArray [61][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][3].cb_test                                      ;
                vSys2PeArray [61][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][4].cb_test                                      ;
                vSys2PeArray [61][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][5].cb_test                                      ;
                vSys2PeArray [61][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][6].cb_test                                      ;
                vSys2PeArray [61][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][7].cb_test                                      ;
                vSys2PeArray [61][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][8].cb_test                                      ;
                vSys2PeArray [61][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][9].cb_test                                      ;
                vSys2PeArray [61][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][10].cb_test                                      ;
                vSys2PeArray [61][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][11].cb_test                                      ;
                vSys2PeArray [61][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][12].cb_test                                      ;
                vSys2PeArray [61][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][13].cb_test                                      ;
                vSys2PeArray [61][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][14].cb_test                                      ;
                vSys2PeArray [61][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][15].cb_test                                      ;
                vSys2PeArray [61][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][16].cb_test                                      ;
                vSys2PeArray [61][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][17].cb_test                                      ;
                vSys2PeArray [61][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][18].cb_test                                      ;
                vSys2PeArray [61][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][19].cb_test                                      ;
                vSys2PeArray [61][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][20].cb_test                                      ;
                vSys2PeArray [61][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][21].cb_test                                      ;
                vSys2PeArray [61][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][22].cb_test                                      ;
                vSys2PeArray [61][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][23].cb_test                                      ;
                vSys2PeArray [61][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][24].cb_test                                      ;
                vSys2PeArray [61][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][25].cb_test                                      ;
                vSys2PeArray [61][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][26].cb_test                                      ;
                vSys2PeArray [61][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][27].cb_test                                      ;
                vSys2PeArray [61][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][28].cb_test                                      ;
                vSys2PeArray [61][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][29].cb_test                                      ;
                vSys2PeArray [61][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][30].cb_test                                      ;
                vSys2PeArray [61][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[61][31].cb_test                                      ;
                vSys2PeArray [61][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [61][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[62][0].cb_test                                      ;
                vSys2PeArray [62][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][1].cb_test                                      ;
                vSys2PeArray [62][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][2].cb_test                                      ;
                vSys2PeArray [62][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][3].cb_test                                      ;
                vSys2PeArray [62][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][4].cb_test                                      ;
                vSys2PeArray [62][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][5].cb_test                                      ;
                vSys2PeArray [62][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][6].cb_test                                      ;
                vSys2PeArray [62][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][7].cb_test                                      ;
                vSys2PeArray [62][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][8].cb_test                                      ;
                vSys2PeArray [62][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][9].cb_test                                      ;
                vSys2PeArray [62][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][10].cb_test                                      ;
                vSys2PeArray [62][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][11].cb_test                                      ;
                vSys2PeArray [62][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][12].cb_test                                      ;
                vSys2PeArray [62][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][13].cb_test                                      ;
                vSys2PeArray [62][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][14].cb_test                                      ;
                vSys2PeArray [62][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][15].cb_test                                      ;
                vSys2PeArray [62][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][16].cb_test                                      ;
                vSys2PeArray [62][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][17].cb_test                                      ;
                vSys2PeArray [62][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][18].cb_test                                      ;
                vSys2PeArray [62][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][19].cb_test                                      ;
                vSys2PeArray [62][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][20].cb_test                                      ;
                vSys2PeArray [62][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][21].cb_test                                      ;
                vSys2PeArray [62][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][22].cb_test                                      ;
                vSys2PeArray [62][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][23].cb_test                                      ;
                vSys2PeArray [62][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][24].cb_test                                      ;
                vSys2PeArray [62][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][25].cb_test                                      ;
                vSys2PeArray [62][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][26].cb_test                                      ;
                vSys2PeArray [62][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][27].cb_test                                      ;
                vSys2PeArray [62][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][28].cb_test                                      ;
                vSys2PeArray [62][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][29].cb_test                                      ;
                vSys2PeArray [62][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][30].cb_test                                      ;
                vSys2PeArray [62][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[62][31].cb_test                                      ;
                vSys2PeArray [62][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [62][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end

            begin
                @vSys2PeArray[63][0].cb_test                                      ;
                vSys2PeArray [63][0].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][0].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][1].cb_test                                      ;
                vSys2PeArray [63][1].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][1].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][2].cb_test                                      ;
                vSys2PeArray [63][2].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][2].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][3].cb_test                                      ;
                vSys2PeArray [63][3].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][3].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][4].cb_test                                      ;
                vSys2PeArray [63][4].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][4].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][5].cb_test                                      ;
                vSys2PeArray [63][5].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][5].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][6].cb_test                                      ;
                vSys2PeArray [63][6].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][6].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][7].cb_test                                      ;
                vSys2PeArray [63][7].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][7].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][8].cb_test                                      ;
                vSys2PeArray [63][8].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][8].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][9].cb_test                                      ;
                vSys2PeArray [63][9].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][9].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][10].cb_test                                      ;
                vSys2PeArray [63][10].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][10].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][11].cb_test                                      ;
                vSys2PeArray [63][11].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][11].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][12].cb_test                                      ;
                vSys2PeArray [63][12].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][12].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][13].cb_test                                      ;
                vSys2PeArray [63][13].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][13].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][14].cb_test                                      ;
                vSys2PeArray [63][14].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][14].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][15].cb_test                                      ;
                vSys2PeArray [63][15].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][15].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][16].cb_test                                      ;
                vSys2PeArray [63][16].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][16].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][17].cb_test                                      ;
                vSys2PeArray [63][17].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][17].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][18].cb_test                                      ;
                vSys2PeArray [63][18].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][18].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][19].cb_test                                      ;
                vSys2PeArray [63][19].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][19].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][20].cb_test                                      ;
                vSys2PeArray [63][20].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][20].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][21].cb_test                                      ;
                vSys2PeArray [63][21].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][21].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][22].cb_test                                      ;
                vSys2PeArray [63][22].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][22].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][23].cb_test                                      ;
                vSys2PeArray [63][23].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][23].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][24].cb_test                                      ;
                vSys2PeArray [63][24].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][24].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][25].cb_test                                      ;
                vSys2PeArray [63][25].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][25].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][26].cb_test                                      ;
                vSys2PeArray [63][26].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][26].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][27].cb_test                                      ;
                vSys2PeArray [63][27].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][27].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][28].cb_test                                      ;
                vSys2PeArray [63][28].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][28].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][29].cb_test                                      ;
                vSys2PeArray [63][29].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][29].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][30].cb_test                                      ;
                vSys2PeArray [63][30].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][30].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
            begin
                @vSys2PeArray[63][31].cb_test                                      ;
                vSys2PeArray [63][31].cb_test.std__pe__lane_strm0_data_valid  <= 0  ;
                vSys2PeArray [63][31].cb_test.std__pe__lane_strm1_data_valid  <= 0  ;
            end
