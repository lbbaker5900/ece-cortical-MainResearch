
       // lane0 NoC to stOp 
      .sdp__cntl__lane0_strm_ready          ( sdp__cntl__lane0_strm_ready         ), 
      .cntl__sdp__lane0_strm_cntl           ( cntl__sdp__lane0_strm_cntl          ), 
      .cntl__sdp__lane0_strm_id             ( cntl__sdp__lane0_strm_id            ), 
      .cntl__sdp__lane0_strm_data           ( cntl__sdp__lane0_strm_data          ), 
      .cntl__sdp__lane0_strm_data_valid     ( cntl__sdp__lane0_strm_data_valid    ), 
       // lane0 stOp to NoC 
      .cntl__sdp__lane0_strm_ready          ( cntl__sdp__lane0_strm_ready         ), 
      .sdp__cntl__lane0_strm_cntl           ( sdp__cntl__lane0_strm_cntl          ), 
      .sdp__cntl__lane0_strm_id             ( sdp__cntl__lane0_strm_id            ), 
      .sdp__cntl__lane0_strm_data           ( sdp__cntl__lane0_strm_data          ), 
      .sdp__cntl__lane0_strm_data_valid     ( sdp__cntl__lane0_strm_data_valid    ), 
       // lane1 NoC to stOp 
      .sdp__cntl__lane1_strm_ready          ( sdp__cntl__lane1_strm_ready         ), 
      .cntl__sdp__lane1_strm_cntl           ( cntl__sdp__lane1_strm_cntl          ), 
      .cntl__sdp__lane1_strm_id             ( cntl__sdp__lane1_strm_id            ), 
      .cntl__sdp__lane1_strm_data           ( cntl__sdp__lane1_strm_data          ), 
      .cntl__sdp__lane1_strm_data_valid     ( cntl__sdp__lane1_strm_data_valid    ), 
       // lane1 stOp to NoC 
      .cntl__sdp__lane1_strm_ready          ( cntl__sdp__lane1_strm_ready         ), 
      .sdp__cntl__lane1_strm_cntl           ( sdp__cntl__lane1_strm_cntl          ), 
      .sdp__cntl__lane1_strm_id             ( sdp__cntl__lane1_strm_id            ), 
      .sdp__cntl__lane1_strm_data           ( sdp__cntl__lane1_strm_data          ), 
      .sdp__cntl__lane1_strm_data_valid     ( sdp__cntl__lane1_strm_data_valid    ), 
       // lane2 NoC to stOp 
      .sdp__cntl__lane2_strm_ready          ( sdp__cntl__lane2_strm_ready         ), 
      .cntl__sdp__lane2_strm_cntl           ( cntl__sdp__lane2_strm_cntl          ), 
      .cntl__sdp__lane2_strm_id             ( cntl__sdp__lane2_strm_id            ), 
      .cntl__sdp__lane2_strm_data           ( cntl__sdp__lane2_strm_data          ), 
      .cntl__sdp__lane2_strm_data_valid     ( cntl__sdp__lane2_strm_data_valid    ), 
       // lane2 stOp to NoC 
      .cntl__sdp__lane2_strm_ready          ( cntl__sdp__lane2_strm_ready         ), 
      .sdp__cntl__lane2_strm_cntl           ( sdp__cntl__lane2_strm_cntl          ), 
      .sdp__cntl__lane2_strm_id             ( sdp__cntl__lane2_strm_id            ), 
      .sdp__cntl__lane2_strm_data           ( sdp__cntl__lane2_strm_data          ), 
      .sdp__cntl__lane2_strm_data_valid     ( sdp__cntl__lane2_strm_data_valid    ), 
       // lane3 NoC to stOp 
      .sdp__cntl__lane3_strm_ready          ( sdp__cntl__lane3_strm_ready         ), 
      .cntl__sdp__lane3_strm_cntl           ( cntl__sdp__lane3_strm_cntl          ), 
      .cntl__sdp__lane3_strm_id             ( cntl__sdp__lane3_strm_id            ), 
      .cntl__sdp__lane3_strm_data           ( cntl__sdp__lane3_strm_data          ), 
      .cntl__sdp__lane3_strm_data_valid     ( cntl__sdp__lane3_strm_data_valid    ), 
       // lane3 stOp to NoC 
      .cntl__sdp__lane3_strm_ready          ( cntl__sdp__lane3_strm_ready         ), 
      .sdp__cntl__lane3_strm_cntl           ( sdp__cntl__lane3_strm_cntl          ), 
      .sdp__cntl__lane3_strm_id             ( sdp__cntl__lane3_strm_id            ), 
      .sdp__cntl__lane3_strm_data           ( sdp__cntl__lane3_strm_data          ), 
      .sdp__cntl__lane3_strm_data_valid     ( sdp__cntl__lane3_strm_data_valid    ), 
       // lane4 NoC to stOp 
      .sdp__cntl__lane4_strm_ready          ( sdp__cntl__lane4_strm_ready         ), 
      .cntl__sdp__lane4_strm_cntl           ( cntl__sdp__lane4_strm_cntl          ), 
      .cntl__sdp__lane4_strm_id             ( cntl__sdp__lane4_strm_id            ), 
      .cntl__sdp__lane4_strm_data           ( cntl__sdp__lane4_strm_data          ), 
      .cntl__sdp__lane4_strm_data_valid     ( cntl__sdp__lane4_strm_data_valid    ), 
       // lane4 stOp to NoC 
      .cntl__sdp__lane4_strm_ready          ( cntl__sdp__lane4_strm_ready         ), 
      .sdp__cntl__lane4_strm_cntl           ( sdp__cntl__lane4_strm_cntl          ), 
      .sdp__cntl__lane4_strm_id             ( sdp__cntl__lane4_strm_id            ), 
      .sdp__cntl__lane4_strm_data           ( sdp__cntl__lane4_strm_data          ), 
      .sdp__cntl__lane4_strm_data_valid     ( sdp__cntl__lane4_strm_data_valid    ), 
       // lane5 NoC to stOp 
      .sdp__cntl__lane5_strm_ready          ( sdp__cntl__lane5_strm_ready         ), 
      .cntl__sdp__lane5_strm_cntl           ( cntl__sdp__lane5_strm_cntl          ), 
      .cntl__sdp__lane5_strm_id             ( cntl__sdp__lane5_strm_id            ), 
      .cntl__sdp__lane5_strm_data           ( cntl__sdp__lane5_strm_data          ), 
      .cntl__sdp__lane5_strm_data_valid     ( cntl__sdp__lane5_strm_data_valid    ), 
       // lane5 stOp to NoC 
      .cntl__sdp__lane5_strm_ready          ( cntl__sdp__lane5_strm_ready         ), 
      .sdp__cntl__lane5_strm_cntl           ( sdp__cntl__lane5_strm_cntl          ), 
      .sdp__cntl__lane5_strm_id             ( sdp__cntl__lane5_strm_id            ), 
      .sdp__cntl__lane5_strm_data           ( sdp__cntl__lane5_strm_data          ), 
      .sdp__cntl__lane5_strm_data_valid     ( sdp__cntl__lane5_strm_data_valid    ), 
       // lane6 NoC to stOp 
      .sdp__cntl__lane6_strm_ready          ( sdp__cntl__lane6_strm_ready         ), 
      .cntl__sdp__lane6_strm_cntl           ( cntl__sdp__lane6_strm_cntl          ), 
      .cntl__sdp__lane6_strm_id             ( cntl__sdp__lane6_strm_id            ), 
      .cntl__sdp__lane6_strm_data           ( cntl__sdp__lane6_strm_data          ), 
      .cntl__sdp__lane6_strm_data_valid     ( cntl__sdp__lane6_strm_data_valid    ), 
       // lane6 stOp to NoC 
      .cntl__sdp__lane6_strm_ready          ( cntl__sdp__lane6_strm_ready         ), 
      .sdp__cntl__lane6_strm_cntl           ( sdp__cntl__lane6_strm_cntl          ), 
      .sdp__cntl__lane6_strm_id             ( sdp__cntl__lane6_strm_id            ), 
      .sdp__cntl__lane6_strm_data           ( sdp__cntl__lane6_strm_data          ), 
      .sdp__cntl__lane6_strm_data_valid     ( sdp__cntl__lane6_strm_data_valid    ), 
       // lane7 NoC to stOp 
      .sdp__cntl__lane7_strm_ready          ( sdp__cntl__lane7_strm_ready         ), 
      .cntl__sdp__lane7_strm_cntl           ( cntl__sdp__lane7_strm_cntl          ), 
      .cntl__sdp__lane7_strm_id             ( cntl__sdp__lane7_strm_id            ), 
      .cntl__sdp__lane7_strm_data           ( cntl__sdp__lane7_strm_data          ), 
      .cntl__sdp__lane7_strm_data_valid     ( cntl__sdp__lane7_strm_data_valid    ), 
       // lane7 stOp to NoC 
      .cntl__sdp__lane7_strm_ready          ( cntl__sdp__lane7_strm_ready         ), 
      .sdp__cntl__lane7_strm_cntl           ( sdp__cntl__lane7_strm_cntl          ), 
      .sdp__cntl__lane7_strm_id             ( sdp__cntl__lane7_strm_id            ), 
      .sdp__cntl__lane7_strm_data           ( sdp__cntl__lane7_strm_data          ), 
      .sdp__cntl__lane7_strm_data_valid     ( sdp__cntl__lane7_strm_data_valid    ), 
       // lane8 NoC to stOp 
      .sdp__cntl__lane8_strm_ready          ( sdp__cntl__lane8_strm_ready         ), 
      .cntl__sdp__lane8_strm_cntl           ( cntl__sdp__lane8_strm_cntl          ), 
      .cntl__sdp__lane8_strm_id             ( cntl__sdp__lane8_strm_id            ), 
      .cntl__sdp__lane8_strm_data           ( cntl__sdp__lane8_strm_data          ), 
      .cntl__sdp__lane8_strm_data_valid     ( cntl__sdp__lane8_strm_data_valid    ), 
       // lane8 stOp to NoC 
      .cntl__sdp__lane8_strm_ready          ( cntl__sdp__lane8_strm_ready         ), 
      .sdp__cntl__lane8_strm_cntl           ( sdp__cntl__lane8_strm_cntl          ), 
      .sdp__cntl__lane8_strm_id             ( sdp__cntl__lane8_strm_id            ), 
      .sdp__cntl__lane8_strm_data           ( sdp__cntl__lane8_strm_data          ), 
      .sdp__cntl__lane8_strm_data_valid     ( sdp__cntl__lane8_strm_data_valid    ), 
       // lane9 NoC to stOp 
      .sdp__cntl__lane9_strm_ready          ( sdp__cntl__lane9_strm_ready         ), 
      .cntl__sdp__lane9_strm_cntl           ( cntl__sdp__lane9_strm_cntl          ), 
      .cntl__sdp__lane9_strm_id             ( cntl__sdp__lane9_strm_id            ), 
      .cntl__sdp__lane9_strm_data           ( cntl__sdp__lane9_strm_data          ), 
      .cntl__sdp__lane9_strm_data_valid     ( cntl__sdp__lane9_strm_data_valid    ), 
       // lane9 stOp to NoC 
      .cntl__sdp__lane9_strm_ready          ( cntl__sdp__lane9_strm_ready         ), 
      .sdp__cntl__lane9_strm_cntl           ( sdp__cntl__lane9_strm_cntl          ), 
      .sdp__cntl__lane9_strm_id             ( sdp__cntl__lane9_strm_id            ), 
      .sdp__cntl__lane9_strm_data           ( sdp__cntl__lane9_strm_data          ), 
      .sdp__cntl__lane9_strm_data_valid     ( sdp__cntl__lane9_strm_data_valid    ), 
       // lane10 NoC to stOp 
      .sdp__cntl__lane10_strm_ready          ( sdp__cntl__lane10_strm_ready         ), 
      .cntl__sdp__lane10_strm_cntl           ( cntl__sdp__lane10_strm_cntl          ), 
      .cntl__sdp__lane10_strm_id             ( cntl__sdp__lane10_strm_id            ), 
      .cntl__sdp__lane10_strm_data           ( cntl__sdp__lane10_strm_data          ), 
      .cntl__sdp__lane10_strm_data_valid     ( cntl__sdp__lane10_strm_data_valid    ), 
       // lane10 stOp to NoC 
      .cntl__sdp__lane10_strm_ready          ( cntl__sdp__lane10_strm_ready         ), 
      .sdp__cntl__lane10_strm_cntl           ( sdp__cntl__lane10_strm_cntl          ), 
      .sdp__cntl__lane10_strm_id             ( sdp__cntl__lane10_strm_id            ), 
      .sdp__cntl__lane10_strm_data           ( sdp__cntl__lane10_strm_data          ), 
      .sdp__cntl__lane10_strm_data_valid     ( sdp__cntl__lane10_strm_data_valid    ), 
       // lane11 NoC to stOp 
      .sdp__cntl__lane11_strm_ready          ( sdp__cntl__lane11_strm_ready         ), 
      .cntl__sdp__lane11_strm_cntl           ( cntl__sdp__lane11_strm_cntl          ), 
      .cntl__sdp__lane11_strm_id             ( cntl__sdp__lane11_strm_id            ), 
      .cntl__sdp__lane11_strm_data           ( cntl__sdp__lane11_strm_data          ), 
      .cntl__sdp__lane11_strm_data_valid     ( cntl__sdp__lane11_strm_data_valid    ), 
       // lane11 stOp to NoC 
      .cntl__sdp__lane11_strm_ready          ( cntl__sdp__lane11_strm_ready         ), 
      .sdp__cntl__lane11_strm_cntl           ( sdp__cntl__lane11_strm_cntl          ), 
      .sdp__cntl__lane11_strm_id             ( sdp__cntl__lane11_strm_id            ), 
      .sdp__cntl__lane11_strm_data           ( sdp__cntl__lane11_strm_data          ), 
      .sdp__cntl__lane11_strm_data_valid     ( sdp__cntl__lane11_strm_data_valid    ), 
       // lane12 NoC to stOp 
      .sdp__cntl__lane12_strm_ready          ( sdp__cntl__lane12_strm_ready         ), 
      .cntl__sdp__lane12_strm_cntl           ( cntl__sdp__lane12_strm_cntl          ), 
      .cntl__sdp__lane12_strm_id             ( cntl__sdp__lane12_strm_id            ), 
      .cntl__sdp__lane12_strm_data           ( cntl__sdp__lane12_strm_data          ), 
      .cntl__sdp__lane12_strm_data_valid     ( cntl__sdp__lane12_strm_data_valid    ), 
       // lane12 stOp to NoC 
      .cntl__sdp__lane12_strm_ready          ( cntl__sdp__lane12_strm_ready         ), 
      .sdp__cntl__lane12_strm_cntl           ( sdp__cntl__lane12_strm_cntl          ), 
      .sdp__cntl__lane12_strm_id             ( sdp__cntl__lane12_strm_id            ), 
      .sdp__cntl__lane12_strm_data           ( sdp__cntl__lane12_strm_data          ), 
      .sdp__cntl__lane12_strm_data_valid     ( sdp__cntl__lane12_strm_data_valid    ), 
       // lane13 NoC to stOp 
      .sdp__cntl__lane13_strm_ready          ( sdp__cntl__lane13_strm_ready         ), 
      .cntl__sdp__lane13_strm_cntl           ( cntl__sdp__lane13_strm_cntl          ), 
      .cntl__sdp__lane13_strm_id             ( cntl__sdp__lane13_strm_id            ), 
      .cntl__sdp__lane13_strm_data           ( cntl__sdp__lane13_strm_data          ), 
      .cntl__sdp__lane13_strm_data_valid     ( cntl__sdp__lane13_strm_data_valid    ), 
       // lane13 stOp to NoC 
      .cntl__sdp__lane13_strm_ready          ( cntl__sdp__lane13_strm_ready         ), 
      .sdp__cntl__lane13_strm_cntl           ( sdp__cntl__lane13_strm_cntl          ), 
      .sdp__cntl__lane13_strm_id             ( sdp__cntl__lane13_strm_id            ), 
      .sdp__cntl__lane13_strm_data           ( sdp__cntl__lane13_strm_data          ), 
      .sdp__cntl__lane13_strm_data_valid     ( sdp__cntl__lane13_strm_data_valid    ), 
       // lane14 NoC to stOp 
      .sdp__cntl__lane14_strm_ready          ( sdp__cntl__lane14_strm_ready         ), 
      .cntl__sdp__lane14_strm_cntl           ( cntl__sdp__lane14_strm_cntl          ), 
      .cntl__sdp__lane14_strm_id             ( cntl__sdp__lane14_strm_id            ), 
      .cntl__sdp__lane14_strm_data           ( cntl__sdp__lane14_strm_data          ), 
      .cntl__sdp__lane14_strm_data_valid     ( cntl__sdp__lane14_strm_data_valid    ), 
       // lane14 stOp to NoC 
      .cntl__sdp__lane14_strm_ready          ( cntl__sdp__lane14_strm_ready         ), 
      .sdp__cntl__lane14_strm_cntl           ( sdp__cntl__lane14_strm_cntl          ), 
      .sdp__cntl__lane14_strm_id             ( sdp__cntl__lane14_strm_id            ), 
      .sdp__cntl__lane14_strm_data           ( sdp__cntl__lane14_strm_data          ), 
      .sdp__cntl__lane14_strm_data_valid     ( sdp__cntl__lane14_strm_data_valid    ), 
       // lane15 NoC to stOp 
      .sdp__cntl__lane15_strm_ready          ( sdp__cntl__lane15_strm_ready         ), 
      .cntl__sdp__lane15_strm_cntl           ( cntl__sdp__lane15_strm_cntl          ), 
      .cntl__sdp__lane15_strm_id             ( cntl__sdp__lane15_strm_id            ), 
      .cntl__sdp__lane15_strm_data           ( cntl__sdp__lane15_strm_data          ), 
      .cntl__sdp__lane15_strm_data_valid     ( cntl__sdp__lane15_strm_data_valid    ), 
       // lane15 stOp to NoC 
      .cntl__sdp__lane15_strm_ready          ( cntl__sdp__lane15_strm_ready         ), 
      .sdp__cntl__lane15_strm_cntl           ( sdp__cntl__lane15_strm_cntl          ), 
      .sdp__cntl__lane15_strm_id             ( sdp__cntl__lane15_strm_id            ), 
      .sdp__cntl__lane15_strm_data           ( sdp__cntl__lane15_strm_data          ), 
      .sdp__cntl__lane15_strm_data_valid     ( sdp__cntl__lane15_strm_data_valid    ), 
       // lane16 NoC to stOp 
      .sdp__cntl__lane16_strm_ready          ( sdp__cntl__lane16_strm_ready         ), 
      .cntl__sdp__lane16_strm_cntl           ( cntl__sdp__lane16_strm_cntl          ), 
      .cntl__sdp__lane16_strm_id             ( cntl__sdp__lane16_strm_id            ), 
      .cntl__sdp__lane16_strm_data           ( cntl__sdp__lane16_strm_data          ), 
      .cntl__sdp__lane16_strm_data_valid     ( cntl__sdp__lane16_strm_data_valid    ), 
       // lane16 stOp to NoC 
      .cntl__sdp__lane16_strm_ready          ( cntl__sdp__lane16_strm_ready         ), 
      .sdp__cntl__lane16_strm_cntl           ( sdp__cntl__lane16_strm_cntl          ), 
      .sdp__cntl__lane16_strm_id             ( sdp__cntl__lane16_strm_id            ), 
      .sdp__cntl__lane16_strm_data           ( sdp__cntl__lane16_strm_data          ), 
      .sdp__cntl__lane16_strm_data_valid     ( sdp__cntl__lane16_strm_data_valid    ), 
       // lane17 NoC to stOp 
      .sdp__cntl__lane17_strm_ready          ( sdp__cntl__lane17_strm_ready         ), 
      .cntl__sdp__lane17_strm_cntl           ( cntl__sdp__lane17_strm_cntl          ), 
      .cntl__sdp__lane17_strm_id             ( cntl__sdp__lane17_strm_id            ), 
      .cntl__sdp__lane17_strm_data           ( cntl__sdp__lane17_strm_data          ), 
      .cntl__sdp__lane17_strm_data_valid     ( cntl__sdp__lane17_strm_data_valid    ), 
       // lane17 stOp to NoC 
      .cntl__sdp__lane17_strm_ready          ( cntl__sdp__lane17_strm_ready         ), 
      .sdp__cntl__lane17_strm_cntl           ( sdp__cntl__lane17_strm_cntl          ), 
      .sdp__cntl__lane17_strm_id             ( sdp__cntl__lane17_strm_id            ), 
      .sdp__cntl__lane17_strm_data           ( sdp__cntl__lane17_strm_data          ), 
      .sdp__cntl__lane17_strm_data_valid     ( sdp__cntl__lane17_strm_data_valid    ), 
       // lane18 NoC to stOp 
      .sdp__cntl__lane18_strm_ready          ( sdp__cntl__lane18_strm_ready         ), 
      .cntl__sdp__lane18_strm_cntl           ( cntl__sdp__lane18_strm_cntl          ), 
      .cntl__sdp__lane18_strm_id             ( cntl__sdp__lane18_strm_id            ), 
      .cntl__sdp__lane18_strm_data           ( cntl__sdp__lane18_strm_data          ), 
      .cntl__sdp__lane18_strm_data_valid     ( cntl__sdp__lane18_strm_data_valid    ), 
       // lane18 stOp to NoC 
      .cntl__sdp__lane18_strm_ready          ( cntl__sdp__lane18_strm_ready         ), 
      .sdp__cntl__lane18_strm_cntl           ( sdp__cntl__lane18_strm_cntl          ), 
      .sdp__cntl__lane18_strm_id             ( sdp__cntl__lane18_strm_id            ), 
      .sdp__cntl__lane18_strm_data           ( sdp__cntl__lane18_strm_data          ), 
      .sdp__cntl__lane18_strm_data_valid     ( sdp__cntl__lane18_strm_data_valid    ), 
       // lane19 NoC to stOp 
      .sdp__cntl__lane19_strm_ready          ( sdp__cntl__lane19_strm_ready         ), 
      .cntl__sdp__lane19_strm_cntl           ( cntl__sdp__lane19_strm_cntl          ), 
      .cntl__sdp__lane19_strm_id             ( cntl__sdp__lane19_strm_id            ), 
      .cntl__sdp__lane19_strm_data           ( cntl__sdp__lane19_strm_data          ), 
      .cntl__sdp__lane19_strm_data_valid     ( cntl__sdp__lane19_strm_data_valid    ), 
       // lane19 stOp to NoC 
      .cntl__sdp__lane19_strm_ready          ( cntl__sdp__lane19_strm_ready         ), 
      .sdp__cntl__lane19_strm_cntl           ( sdp__cntl__lane19_strm_cntl          ), 
      .sdp__cntl__lane19_strm_id             ( sdp__cntl__lane19_strm_id            ), 
      .sdp__cntl__lane19_strm_data           ( sdp__cntl__lane19_strm_data          ), 
      .sdp__cntl__lane19_strm_data_valid     ( sdp__cntl__lane19_strm_data_valid    ), 
       // lane20 NoC to stOp 
      .sdp__cntl__lane20_strm_ready          ( sdp__cntl__lane20_strm_ready         ), 
      .cntl__sdp__lane20_strm_cntl           ( cntl__sdp__lane20_strm_cntl          ), 
      .cntl__sdp__lane20_strm_id             ( cntl__sdp__lane20_strm_id            ), 
      .cntl__sdp__lane20_strm_data           ( cntl__sdp__lane20_strm_data          ), 
      .cntl__sdp__lane20_strm_data_valid     ( cntl__sdp__lane20_strm_data_valid    ), 
       // lane20 stOp to NoC 
      .cntl__sdp__lane20_strm_ready          ( cntl__sdp__lane20_strm_ready         ), 
      .sdp__cntl__lane20_strm_cntl           ( sdp__cntl__lane20_strm_cntl          ), 
      .sdp__cntl__lane20_strm_id             ( sdp__cntl__lane20_strm_id            ), 
      .sdp__cntl__lane20_strm_data           ( sdp__cntl__lane20_strm_data          ), 
      .sdp__cntl__lane20_strm_data_valid     ( sdp__cntl__lane20_strm_data_valid    ), 
       // lane21 NoC to stOp 
      .sdp__cntl__lane21_strm_ready          ( sdp__cntl__lane21_strm_ready         ), 
      .cntl__sdp__lane21_strm_cntl           ( cntl__sdp__lane21_strm_cntl          ), 
      .cntl__sdp__lane21_strm_id             ( cntl__sdp__lane21_strm_id            ), 
      .cntl__sdp__lane21_strm_data           ( cntl__sdp__lane21_strm_data          ), 
      .cntl__sdp__lane21_strm_data_valid     ( cntl__sdp__lane21_strm_data_valid    ), 
       // lane21 stOp to NoC 
      .cntl__sdp__lane21_strm_ready          ( cntl__sdp__lane21_strm_ready         ), 
      .sdp__cntl__lane21_strm_cntl           ( sdp__cntl__lane21_strm_cntl          ), 
      .sdp__cntl__lane21_strm_id             ( sdp__cntl__lane21_strm_id            ), 
      .sdp__cntl__lane21_strm_data           ( sdp__cntl__lane21_strm_data          ), 
      .sdp__cntl__lane21_strm_data_valid     ( sdp__cntl__lane21_strm_data_valid    ), 
       // lane22 NoC to stOp 
      .sdp__cntl__lane22_strm_ready          ( sdp__cntl__lane22_strm_ready         ), 
      .cntl__sdp__lane22_strm_cntl           ( cntl__sdp__lane22_strm_cntl          ), 
      .cntl__sdp__lane22_strm_id             ( cntl__sdp__lane22_strm_id            ), 
      .cntl__sdp__lane22_strm_data           ( cntl__sdp__lane22_strm_data          ), 
      .cntl__sdp__lane22_strm_data_valid     ( cntl__sdp__lane22_strm_data_valid    ), 
       // lane22 stOp to NoC 
      .cntl__sdp__lane22_strm_ready          ( cntl__sdp__lane22_strm_ready         ), 
      .sdp__cntl__lane22_strm_cntl           ( sdp__cntl__lane22_strm_cntl          ), 
      .sdp__cntl__lane22_strm_id             ( sdp__cntl__lane22_strm_id            ), 
      .sdp__cntl__lane22_strm_data           ( sdp__cntl__lane22_strm_data          ), 
      .sdp__cntl__lane22_strm_data_valid     ( sdp__cntl__lane22_strm_data_valid    ), 
       // lane23 NoC to stOp 
      .sdp__cntl__lane23_strm_ready          ( sdp__cntl__lane23_strm_ready         ), 
      .cntl__sdp__lane23_strm_cntl           ( cntl__sdp__lane23_strm_cntl          ), 
      .cntl__sdp__lane23_strm_id             ( cntl__sdp__lane23_strm_id            ), 
      .cntl__sdp__lane23_strm_data           ( cntl__sdp__lane23_strm_data          ), 
      .cntl__sdp__lane23_strm_data_valid     ( cntl__sdp__lane23_strm_data_valid    ), 
       // lane23 stOp to NoC 
      .cntl__sdp__lane23_strm_ready          ( cntl__sdp__lane23_strm_ready         ), 
      .sdp__cntl__lane23_strm_cntl           ( sdp__cntl__lane23_strm_cntl          ), 
      .sdp__cntl__lane23_strm_id             ( sdp__cntl__lane23_strm_id            ), 
      .sdp__cntl__lane23_strm_data           ( sdp__cntl__lane23_strm_data          ), 
      .sdp__cntl__lane23_strm_data_valid     ( sdp__cntl__lane23_strm_data_valid    ), 
       // lane24 NoC to stOp 
      .sdp__cntl__lane24_strm_ready          ( sdp__cntl__lane24_strm_ready         ), 
      .cntl__sdp__lane24_strm_cntl           ( cntl__sdp__lane24_strm_cntl          ), 
      .cntl__sdp__lane24_strm_id             ( cntl__sdp__lane24_strm_id            ), 
      .cntl__sdp__lane24_strm_data           ( cntl__sdp__lane24_strm_data          ), 
      .cntl__sdp__lane24_strm_data_valid     ( cntl__sdp__lane24_strm_data_valid    ), 
       // lane24 stOp to NoC 
      .cntl__sdp__lane24_strm_ready          ( cntl__sdp__lane24_strm_ready         ), 
      .sdp__cntl__lane24_strm_cntl           ( sdp__cntl__lane24_strm_cntl          ), 
      .sdp__cntl__lane24_strm_id             ( sdp__cntl__lane24_strm_id            ), 
      .sdp__cntl__lane24_strm_data           ( sdp__cntl__lane24_strm_data          ), 
      .sdp__cntl__lane24_strm_data_valid     ( sdp__cntl__lane24_strm_data_valid    ), 
       // lane25 NoC to stOp 
      .sdp__cntl__lane25_strm_ready          ( sdp__cntl__lane25_strm_ready         ), 
      .cntl__sdp__lane25_strm_cntl           ( cntl__sdp__lane25_strm_cntl          ), 
      .cntl__sdp__lane25_strm_id             ( cntl__sdp__lane25_strm_id            ), 
      .cntl__sdp__lane25_strm_data           ( cntl__sdp__lane25_strm_data          ), 
      .cntl__sdp__lane25_strm_data_valid     ( cntl__sdp__lane25_strm_data_valid    ), 
       // lane25 stOp to NoC 
      .cntl__sdp__lane25_strm_ready          ( cntl__sdp__lane25_strm_ready         ), 
      .sdp__cntl__lane25_strm_cntl           ( sdp__cntl__lane25_strm_cntl          ), 
      .sdp__cntl__lane25_strm_id             ( sdp__cntl__lane25_strm_id            ), 
      .sdp__cntl__lane25_strm_data           ( sdp__cntl__lane25_strm_data          ), 
      .sdp__cntl__lane25_strm_data_valid     ( sdp__cntl__lane25_strm_data_valid    ), 
       // lane26 NoC to stOp 
      .sdp__cntl__lane26_strm_ready          ( sdp__cntl__lane26_strm_ready         ), 
      .cntl__sdp__lane26_strm_cntl           ( cntl__sdp__lane26_strm_cntl          ), 
      .cntl__sdp__lane26_strm_id             ( cntl__sdp__lane26_strm_id            ), 
      .cntl__sdp__lane26_strm_data           ( cntl__sdp__lane26_strm_data          ), 
      .cntl__sdp__lane26_strm_data_valid     ( cntl__sdp__lane26_strm_data_valid    ), 
       // lane26 stOp to NoC 
      .cntl__sdp__lane26_strm_ready          ( cntl__sdp__lane26_strm_ready         ), 
      .sdp__cntl__lane26_strm_cntl           ( sdp__cntl__lane26_strm_cntl          ), 
      .sdp__cntl__lane26_strm_id             ( sdp__cntl__lane26_strm_id            ), 
      .sdp__cntl__lane26_strm_data           ( sdp__cntl__lane26_strm_data          ), 
      .sdp__cntl__lane26_strm_data_valid     ( sdp__cntl__lane26_strm_data_valid    ), 
       // lane27 NoC to stOp 
      .sdp__cntl__lane27_strm_ready          ( sdp__cntl__lane27_strm_ready         ), 
      .cntl__sdp__lane27_strm_cntl           ( cntl__sdp__lane27_strm_cntl          ), 
      .cntl__sdp__lane27_strm_id             ( cntl__sdp__lane27_strm_id            ), 
      .cntl__sdp__lane27_strm_data           ( cntl__sdp__lane27_strm_data          ), 
      .cntl__sdp__lane27_strm_data_valid     ( cntl__sdp__lane27_strm_data_valid    ), 
       // lane27 stOp to NoC 
      .cntl__sdp__lane27_strm_ready          ( cntl__sdp__lane27_strm_ready         ), 
      .sdp__cntl__lane27_strm_cntl           ( sdp__cntl__lane27_strm_cntl          ), 
      .sdp__cntl__lane27_strm_id             ( sdp__cntl__lane27_strm_id            ), 
      .sdp__cntl__lane27_strm_data           ( sdp__cntl__lane27_strm_data          ), 
      .sdp__cntl__lane27_strm_data_valid     ( sdp__cntl__lane27_strm_data_valid    ), 
       // lane28 NoC to stOp 
      .sdp__cntl__lane28_strm_ready          ( sdp__cntl__lane28_strm_ready         ), 
      .cntl__sdp__lane28_strm_cntl           ( cntl__sdp__lane28_strm_cntl          ), 
      .cntl__sdp__lane28_strm_id             ( cntl__sdp__lane28_strm_id            ), 
      .cntl__sdp__lane28_strm_data           ( cntl__sdp__lane28_strm_data          ), 
      .cntl__sdp__lane28_strm_data_valid     ( cntl__sdp__lane28_strm_data_valid    ), 
       // lane28 stOp to NoC 
      .cntl__sdp__lane28_strm_ready          ( cntl__sdp__lane28_strm_ready         ), 
      .sdp__cntl__lane28_strm_cntl           ( sdp__cntl__lane28_strm_cntl          ), 
      .sdp__cntl__lane28_strm_id             ( sdp__cntl__lane28_strm_id            ), 
      .sdp__cntl__lane28_strm_data           ( sdp__cntl__lane28_strm_data          ), 
      .sdp__cntl__lane28_strm_data_valid     ( sdp__cntl__lane28_strm_data_valid    ), 
       // lane29 NoC to stOp 
      .sdp__cntl__lane29_strm_ready          ( sdp__cntl__lane29_strm_ready         ), 
      .cntl__sdp__lane29_strm_cntl           ( cntl__sdp__lane29_strm_cntl          ), 
      .cntl__sdp__lane29_strm_id             ( cntl__sdp__lane29_strm_id            ), 
      .cntl__sdp__lane29_strm_data           ( cntl__sdp__lane29_strm_data          ), 
      .cntl__sdp__lane29_strm_data_valid     ( cntl__sdp__lane29_strm_data_valid    ), 
       // lane29 stOp to NoC 
      .cntl__sdp__lane29_strm_ready          ( cntl__sdp__lane29_strm_ready         ), 
      .sdp__cntl__lane29_strm_cntl           ( sdp__cntl__lane29_strm_cntl          ), 
      .sdp__cntl__lane29_strm_id             ( sdp__cntl__lane29_strm_id            ), 
      .sdp__cntl__lane29_strm_data           ( sdp__cntl__lane29_strm_data          ), 
      .sdp__cntl__lane29_strm_data_valid     ( sdp__cntl__lane29_strm_data_valid    ), 
       // lane30 NoC to stOp 
      .sdp__cntl__lane30_strm_ready          ( sdp__cntl__lane30_strm_ready         ), 
      .cntl__sdp__lane30_strm_cntl           ( cntl__sdp__lane30_strm_cntl          ), 
      .cntl__sdp__lane30_strm_id             ( cntl__sdp__lane30_strm_id            ), 
      .cntl__sdp__lane30_strm_data           ( cntl__sdp__lane30_strm_data          ), 
      .cntl__sdp__lane30_strm_data_valid     ( cntl__sdp__lane30_strm_data_valid    ), 
       // lane30 stOp to NoC 
      .cntl__sdp__lane30_strm_ready          ( cntl__sdp__lane30_strm_ready         ), 
      .sdp__cntl__lane30_strm_cntl           ( sdp__cntl__lane30_strm_cntl          ), 
      .sdp__cntl__lane30_strm_id             ( sdp__cntl__lane30_strm_id            ), 
      .sdp__cntl__lane30_strm_data           ( sdp__cntl__lane30_strm_data          ), 
      .sdp__cntl__lane30_strm_data_valid     ( sdp__cntl__lane30_strm_data_valid    ), 
       // lane31 NoC to stOp 
      .sdp__cntl__lane31_strm_ready          ( sdp__cntl__lane31_strm_ready         ), 
      .cntl__sdp__lane31_strm_cntl           ( cntl__sdp__lane31_strm_cntl          ), 
      .cntl__sdp__lane31_strm_id             ( cntl__sdp__lane31_strm_id            ), 
      .cntl__sdp__lane31_strm_data           ( cntl__sdp__lane31_strm_data          ), 
      .cntl__sdp__lane31_strm_data_valid     ( cntl__sdp__lane31_strm_data_valid    ), 
       // lane31 stOp to NoC 
      .cntl__sdp__lane31_strm_ready          ( cntl__sdp__lane31_strm_ready         ), 
      .sdp__cntl__lane31_strm_cntl           ( sdp__cntl__lane31_strm_cntl          ), 
      .sdp__cntl__lane31_strm_id             ( sdp__cntl__lane31_strm_id            ), 
      .sdp__cntl__lane31_strm_data           ( sdp__cntl__lane31_strm_data          ), 
      .sdp__cntl__lane31_strm_data_valid     ( sdp__cntl__lane31_strm_data_valid    ), 
