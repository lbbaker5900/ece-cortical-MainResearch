
  // OOB controls how the lanes are interpreted                                  
 assign    std__pe0__oob_cntl    =    mgr0__std__oob_cntl            ;
 assign    std__pe0__oob_valid   =    mgr0__std__oob_valid           ;
 assign    std__mgr0__oob_ready  =    pe0__std__oob_ready            ;
 assign    std__pe0__oob_type    =    mgr0__std__oob_type            ;
 assign    std__pe0__oob_data    =    mgr0__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe1__oob_cntl    =    mgr1__std__oob_cntl            ;
 assign    std__pe1__oob_valid   =    mgr1__std__oob_valid           ;
 assign    std__mgr1__oob_ready  =    pe1__std__oob_ready            ;
 assign    std__pe1__oob_type    =    mgr1__std__oob_type            ;
 assign    std__pe1__oob_data    =    mgr1__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe2__oob_cntl    =    mgr2__std__oob_cntl            ;
 assign    std__pe2__oob_valid   =    mgr2__std__oob_valid           ;
 assign    std__mgr2__oob_ready  =    pe2__std__oob_ready            ;
 assign    std__pe2__oob_type    =    mgr2__std__oob_type            ;
 assign    std__pe2__oob_data    =    mgr2__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe3__oob_cntl    =    mgr3__std__oob_cntl            ;
 assign    std__pe3__oob_valid   =    mgr3__std__oob_valid           ;
 assign    std__mgr3__oob_ready  =    pe3__std__oob_ready            ;
 assign    std__pe3__oob_type    =    mgr3__std__oob_type            ;
 assign    std__pe3__oob_data    =    mgr3__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe4__oob_cntl    =    mgr4__std__oob_cntl            ;
 assign    std__pe4__oob_valid   =    mgr4__std__oob_valid           ;
 assign    std__mgr4__oob_ready  =    pe4__std__oob_ready            ;
 assign    std__pe4__oob_type    =    mgr4__std__oob_type            ;
 assign    std__pe4__oob_data    =    mgr4__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe5__oob_cntl    =    mgr5__std__oob_cntl            ;
 assign    std__pe5__oob_valid   =    mgr5__std__oob_valid           ;
 assign    std__mgr5__oob_ready  =    pe5__std__oob_ready            ;
 assign    std__pe5__oob_type    =    mgr5__std__oob_type            ;
 assign    std__pe5__oob_data    =    mgr5__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe6__oob_cntl    =    mgr6__std__oob_cntl            ;
 assign    std__pe6__oob_valid   =    mgr6__std__oob_valid           ;
 assign    std__mgr6__oob_ready  =    pe6__std__oob_ready            ;
 assign    std__pe6__oob_type    =    mgr6__std__oob_type            ;
 assign    std__pe6__oob_data    =    mgr6__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe7__oob_cntl    =    mgr7__std__oob_cntl            ;
 assign    std__pe7__oob_valid   =    mgr7__std__oob_valid           ;
 assign    std__mgr7__oob_ready  =    pe7__std__oob_ready            ;
 assign    std__pe7__oob_type    =    mgr7__std__oob_type            ;
 assign    std__pe7__oob_data    =    mgr7__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe8__oob_cntl    =    mgr8__std__oob_cntl            ;
 assign    std__pe8__oob_valid   =    mgr8__std__oob_valid           ;
 assign    std__mgr8__oob_ready  =    pe8__std__oob_ready            ;
 assign    std__pe8__oob_type    =    mgr8__std__oob_type            ;
 assign    std__pe8__oob_data    =    mgr8__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe9__oob_cntl    =    mgr9__std__oob_cntl            ;
 assign    std__pe9__oob_valid   =    mgr9__std__oob_valid           ;
 assign    std__mgr9__oob_ready  =    pe9__std__oob_ready            ;
 assign    std__pe9__oob_type    =    mgr9__std__oob_type            ;
 assign    std__pe9__oob_data    =    mgr9__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe10__oob_cntl    =    mgr10__std__oob_cntl            ;
 assign    std__pe10__oob_valid   =    mgr10__std__oob_valid           ;
 assign    std__mgr10__oob_ready  =    pe10__std__oob_ready            ;
 assign    std__pe10__oob_type    =    mgr10__std__oob_type            ;
 assign    std__pe10__oob_data    =    mgr10__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe11__oob_cntl    =    mgr11__std__oob_cntl            ;
 assign    std__pe11__oob_valid   =    mgr11__std__oob_valid           ;
 assign    std__mgr11__oob_ready  =    pe11__std__oob_ready            ;
 assign    std__pe11__oob_type    =    mgr11__std__oob_type            ;
 assign    std__pe11__oob_data    =    mgr11__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe12__oob_cntl    =    mgr12__std__oob_cntl            ;
 assign    std__pe12__oob_valid   =    mgr12__std__oob_valid           ;
 assign    std__mgr12__oob_ready  =    pe12__std__oob_ready            ;
 assign    std__pe12__oob_type    =    mgr12__std__oob_type            ;
 assign    std__pe12__oob_data    =    mgr12__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe13__oob_cntl    =    mgr13__std__oob_cntl            ;
 assign    std__pe13__oob_valid   =    mgr13__std__oob_valid           ;
 assign    std__mgr13__oob_ready  =    pe13__std__oob_ready            ;
 assign    std__pe13__oob_type    =    mgr13__std__oob_type            ;
 assign    std__pe13__oob_data    =    mgr13__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe14__oob_cntl    =    mgr14__std__oob_cntl            ;
 assign    std__pe14__oob_valid   =    mgr14__std__oob_valid           ;
 assign    std__mgr14__oob_ready  =    pe14__std__oob_ready            ;
 assign    std__pe14__oob_type    =    mgr14__std__oob_type            ;
 assign    std__pe14__oob_data    =    mgr14__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe15__oob_cntl    =    mgr15__std__oob_cntl            ;
 assign    std__pe15__oob_valid   =    mgr15__std__oob_valid           ;
 assign    std__mgr15__oob_ready  =    pe15__std__oob_ready            ;
 assign    std__pe15__oob_type    =    mgr15__std__oob_type            ;
 assign    std__pe15__oob_data    =    mgr15__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe16__oob_cntl    =    mgr16__std__oob_cntl            ;
 assign    std__pe16__oob_valid   =    mgr16__std__oob_valid           ;
 assign    std__mgr16__oob_ready  =    pe16__std__oob_ready            ;
 assign    std__pe16__oob_type    =    mgr16__std__oob_type            ;
 assign    std__pe16__oob_data    =    mgr16__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe17__oob_cntl    =    mgr17__std__oob_cntl            ;
 assign    std__pe17__oob_valid   =    mgr17__std__oob_valid           ;
 assign    std__mgr17__oob_ready  =    pe17__std__oob_ready            ;
 assign    std__pe17__oob_type    =    mgr17__std__oob_type            ;
 assign    std__pe17__oob_data    =    mgr17__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe18__oob_cntl    =    mgr18__std__oob_cntl            ;
 assign    std__pe18__oob_valid   =    mgr18__std__oob_valid           ;
 assign    std__mgr18__oob_ready  =    pe18__std__oob_ready            ;
 assign    std__pe18__oob_type    =    mgr18__std__oob_type            ;
 assign    std__pe18__oob_data    =    mgr18__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe19__oob_cntl    =    mgr19__std__oob_cntl            ;
 assign    std__pe19__oob_valid   =    mgr19__std__oob_valid           ;
 assign    std__mgr19__oob_ready  =    pe19__std__oob_ready            ;
 assign    std__pe19__oob_type    =    mgr19__std__oob_type            ;
 assign    std__pe19__oob_data    =    mgr19__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe20__oob_cntl    =    mgr20__std__oob_cntl            ;
 assign    std__pe20__oob_valid   =    mgr20__std__oob_valid           ;
 assign    std__mgr20__oob_ready  =    pe20__std__oob_ready            ;
 assign    std__pe20__oob_type    =    mgr20__std__oob_type            ;
 assign    std__pe20__oob_data    =    mgr20__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe21__oob_cntl    =    mgr21__std__oob_cntl            ;
 assign    std__pe21__oob_valid   =    mgr21__std__oob_valid           ;
 assign    std__mgr21__oob_ready  =    pe21__std__oob_ready            ;
 assign    std__pe21__oob_type    =    mgr21__std__oob_type            ;
 assign    std__pe21__oob_data    =    mgr21__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe22__oob_cntl    =    mgr22__std__oob_cntl            ;
 assign    std__pe22__oob_valid   =    mgr22__std__oob_valid           ;
 assign    std__mgr22__oob_ready  =    pe22__std__oob_ready            ;
 assign    std__pe22__oob_type    =    mgr22__std__oob_type            ;
 assign    std__pe22__oob_data    =    mgr22__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe23__oob_cntl    =    mgr23__std__oob_cntl            ;
 assign    std__pe23__oob_valid   =    mgr23__std__oob_valid           ;
 assign    std__mgr23__oob_ready  =    pe23__std__oob_ready            ;
 assign    std__pe23__oob_type    =    mgr23__std__oob_type            ;
 assign    std__pe23__oob_data    =    mgr23__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe24__oob_cntl    =    mgr24__std__oob_cntl            ;
 assign    std__pe24__oob_valid   =    mgr24__std__oob_valid           ;
 assign    std__mgr24__oob_ready  =    pe24__std__oob_ready            ;
 assign    std__pe24__oob_type    =    mgr24__std__oob_type            ;
 assign    std__pe24__oob_data    =    mgr24__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe25__oob_cntl    =    mgr25__std__oob_cntl            ;
 assign    std__pe25__oob_valid   =    mgr25__std__oob_valid           ;
 assign    std__mgr25__oob_ready  =    pe25__std__oob_ready            ;
 assign    std__pe25__oob_type    =    mgr25__std__oob_type            ;
 assign    std__pe25__oob_data    =    mgr25__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe26__oob_cntl    =    mgr26__std__oob_cntl            ;
 assign    std__pe26__oob_valid   =    mgr26__std__oob_valid           ;
 assign    std__mgr26__oob_ready  =    pe26__std__oob_ready            ;
 assign    std__pe26__oob_type    =    mgr26__std__oob_type            ;
 assign    std__pe26__oob_data    =    mgr26__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe27__oob_cntl    =    mgr27__std__oob_cntl            ;
 assign    std__pe27__oob_valid   =    mgr27__std__oob_valid           ;
 assign    std__mgr27__oob_ready  =    pe27__std__oob_ready            ;
 assign    std__pe27__oob_type    =    mgr27__std__oob_type            ;
 assign    std__pe27__oob_data    =    mgr27__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe28__oob_cntl    =    mgr28__std__oob_cntl            ;
 assign    std__pe28__oob_valid   =    mgr28__std__oob_valid           ;
 assign    std__mgr28__oob_ready  =    pe28__std__oob_ready            ;
 assign    std__pe28__oob_type    =    mgr28__std__oob_type            ;
 assign    std__pe28__oob_data    =    mgr28__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe29__oob_cntl    =    mgr29__std__oob_cntl            ;
 assign    std__pe29__oob_valid   =    mgr29__std__oob_valid           ;
 assign    std__mgr29__oob_ready  =    pe29__std__oob_ready            ;
 assign    std__pe29__oob_type    =    mgr29__std__oob_type            ;
 assign    std__pe29__oob_data    =    mgr29__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe30__oob_cntl    =    mgr30__std__oob_cntl            ;
 assign    std__pe30__oob_valid   =    mgr30__std__oob_valid           ;
 assign    std__mgr30__oob_ready  =    pe30__std__oob_ready            ;
 assign    std__pe30__oob_type    =    mgr30__std__oob_type            ;
 assign    std__pe30__oob_data    =    mgr30__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe31__oob_cntl    =    mgr31__std__oob_cntl            ;
 assign    std__pe31__oob_valid   =    mgr31__std__oob_valid           ;
 assign    std__mgr31__oob_ready  =    pe31__std__oob_ready            ;
 assign    std__pe31__oob_type    =    mgr31__std__oob_type            ;
 assign    std__pe31__oob_data    =    mgr31__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe32__oob_cntl    =    mgr32__std__oob_cntl            ;
 assign    std__pe32__oob_valid   =    mgr32__std__oob_valid           ;
 assign    std__mgr32__oob_ready  =    pe32__std__oob_ready            ;
 assign    std__pe32__oob_type    =    mgr32__std__oob_type            ;
 assign    std__pe32__oob_data    =    mgr32__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe33__oob_cntl    =    mgr33__std__oob_cntl            ;
 assign    std__pe33__oob_valid   =    mgr33__std__oob_valid           ;
 assign    std__mgr33__oob_ready  =    pe33__std__oob_ready            ;
 assign    std__pe33__oob_type    =    mgr33__std__oob_type            ;
 assign    std__pe33__oob_data    =    mgr33__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe34__oob_cntl    =    mgr34__std__oob_cntl            ;
 assign    std__pe34__oob_valid   =    mgr34__std__oob_valid           ;
 assign    std__mgr34__oob_ready  =    pe34__std__oob_ready            ;
 assign    std__pe34__oob_type    =    mgr34__std__oob_type            ;
 assign    std__pe34__oob_data    =    mgr34__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe35__oob_cntl    =    mgr35__std__oob_cntl            ;
 assign    std__pe35__oob_valid   =    mgr35__std__oob_valid           ;
 assign    std__mgr35__oob_ready  =    pe35__std__oob_ready            ;
 assign    std__pe35__oob_type    =    mgr35__std__oob_type            ;
 assign    std__pe35__oob_data    =    mgr35__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe36__oob_cntl    =    mgr36__std__oob_cntl            ;
 assign    std__pe36__oob_valid   =    mgr36__std__oob_valid           ;
 assign    std__mgr36__oob_ready  =    pe36__std__oob_ready            ;
 assign    std__pe36__oob_type    =    mgr36__std__oob_type            ;
 assign    std__pe36__oob_data    =    mgr36__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe37__oob_cntl    =    mgr37__std__oob_cntl            ;
 assign    std__pe37__oob_valid   =    mgr37__std__oob_valid           ;
 assign    std__mgr37__oob_ready  =    pe37__std__oob_ready            ;
 assign    std__pe37__oob_type    =    mgr37__std__oob_type            ;
 assign    std__pe37__oob_data    =    mgr37__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe38__oob_cntl    =    mgr38__std__oob_cntl            ;
 assign    std__pe38__oob_valid   =    mgr38__std__oob_valid           ;
 assign    std__mgr38__oob_ready  =    pe38__std__oob_ready            ;
 assign    std__pe38__oob_type    =    mgr38__std__oob_type            ;
 assign    std__pe38__oob_data    =    mgr38__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe39__oob_cntl    =    mgr39__std__oob_cntl            ;
 assign    std__pe39__oob_valid   =    mgr39__std__oob_valid           ;
 assign    std__mgr39__oob_ready  =    pe39__std__oob_ready            ;
 assign    std__pe39__oob_type    =    mgr39__std__oob_type            ;
 assign    std__pe39__oob_data    =    mgr39__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe40__oob_cntl    =    mgr40__std__oob_cntl            ;
 assign    std__pe40__oob_valid   =    mgr40__std__oob_valid           ;
 assign    std__mgr40__oob_ready  =    pe40__std__oob_ready            ;
 assign    std__pe40__oob_type    =    mgr40__std__oob_type            ;
 assign    std__pe40__oob_data    =    mgr40__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe41__oob_cntl    =    mgr41__std__oob_cntl            ;
 assign    std__pe41__oob_valid   =    mgr41__std__oob_valid           ;
 assign    std__mgr41__oob_ready  =    pe41__std__oob_ready            ;
 assign    std__pe41__oob_type    =    mgr41__std__oob_type            ;
 assign    std__pe41__oob_data    =    mgr41__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe42__oob_cntl    =    mgr42__std__oob_cntl            ;
 assign    std__pe42__oob_valid   =    mgr42__std__oob_valid           ;
 assign    std__mgr42__oob_ready  =    pe42__std__oob_ready            ;
 assign    std__pe42__oob_type    =    mgr42__std__oob_type            ;
 assign    std__pe42__oob_data    =    mgr42__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe43__oob_cntl    =    mgr43__std__oob_cntl            ;
 assign    std__pe43__oob_valid   =    mgr43__std__oob_valid           ;
 assign    std__mgr43__oob_ready  =    pe43__std__oob_ready            ;
 assign    std__pe43__oob_type    =    mgr43__std__oob_type            ;
 assign    std__pe43__oob_data    =    mgr43__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe44__oob_cntl    =    mgr44__std__oob_cntl            ;
 assign    std__pe44__oob_valid   =    mgr44__std__oob_valid           ;
 assign    std__mgr44__oob_ready  =    pe44__std__oob_ready            ;
 assign    std__pe44__oob_type    =    mgr44__std__oob_type            ;
 assign    std__pe44__oob_data    =    mgr44__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe45__oob_cntl    =    mgr45__std__oob_cntl            ;
 assign    std__pe45__oob_valid   =    mgr45__std__oob_valid           ;
 assign    std__mgr45__oob_ready  =    pe45__std__oob_ready            ;
 assign    std__pe45__oob_type    =    mgr45__std__oob_type            ;
 assign    std__pe45__oob_data    =    mgr45__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe46__oob_cntl    =    mgr46__std__oob_cntl            ;
 assign    std__pe46__oob_valid   =    mgr46__std__oob_valid           ;
 assign    std__mgr46__oob_ready  =    pe46__std__oob_ready            ;
 assign    std__pe46__oob_type    =    mgr46__std__oob_type            ;
 assign    std__pe46__oob_data    =    mgr46__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe47__oob_cntl    =    mgr47__std__oob_cntl            ;
 assign    std__pe47__oob_valid   =    mgr47__std__oob_valid           ;
 assign    std__mgr47__oob_ready  =    pe47__std__oob_ready            ;
 assign    std__pe47__oob_type    =    mgr47__std__oob_type            ;
 assign    std__pe47__oob_data    =    mgr47__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe48__oob_cntl    =    mgr48__std__oob_cntl            ;
 assign    std__pe48__oob_valid   =    mgr48__std__oob_valid           ;
 assign    std__mgr48__oob_ready  =    pe48__std__oob_ready            ;
 assign    std__pe48__oob_type    =    mgr48__std__oob_type            ;
 assign    std__pe48__oob_data    =    mgr48__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe49__oob_cntl    =    mgr49__std__oob_cntl            ;
 assign    std__pe49__oob_valid   =    mgr49__std__oob_valid           ;
 assign    std__mgr49__oob_ready  =    pe49__std__oob_ready            ;
 assign    std__pe49__oob_type    =    mgr49__std__oob_type            ;
 assign    std__pe49__oob_data    =    mgr49__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe50__oob_cntl    =    mgr50__std__oob_cntl            ;
 assign    std__pe50__oob_valid   =    mgr50__std__oob_valid           ;
 assign    std__mgr50__oob_ready  =    pe50__std__oob_ready            ;
 assign    std__pe50__oob_type    =    mgr50__std__oob_type            ;
 assign    std__pe50__oob_data    =    mgr50__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe51__oob_cntl    =    mgr51__std__oob_cntl            ;
 assign    std__pe51__oob_valid   =    mgr51__std__oob_valid           ;
 assign    std__mgr51__oob_ready  =    pe51__std__oob_ready            ;
 assign    std__pe51__oob_type    =    mgr51__std__oob_type            ;
 assign    std__pe51__oob_data    =    mgr51__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe52__oob_cntl    =    mgr52__std__oob_cntl            ;
 assign    std__pe52__oob_valid   =    mgr52__std__oob_valid           ;
 assign    std__mgr52__oob_ready  =    pe52__std__oob_ready            ;
 assign    std__pe52__oob_type    =    mgr52__std__oob_type            ;
 assign    std__pe52__oob_data    =    mgr52__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe53__oob_cntl    =    mgr53__std__oob_cntl            ;
 assign    std__pe53__oob_valid   =    mgr53__std__oob_valid           ;
 assign    std__mgr53__oob_ready  =    pe53__std__oob_ready            ;
 assign    std__pe53__oob_type    =    mgr53__std__oob_type            ;
 assign    std__pe53__oob_data    =    mgr53__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe54__oob_cntl    =    mgr54__std__oob_cntl            ;
 assign    std__pe54__oob_valid   =    mgr54__std__oob_valid           ;
 assign    std__mgr54__oob_ready  =    pe54__std__oob_ready            ;
 assign    std__pe54__oob_type    =    mgr54__std__oob_type            ;
 assign    std__pe54__oob_data    =    mgr54__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe55__oob_cntl    =    mgr55__std__oob_cntl            ;
 assign    std__pe55__oob_valid   =    mgr55__std__oob_valid           ;
 assign    std__mgr55__oob_ready  =    pe55__std__oob_ready            ;
 assign    std__pe55__oob_type    =    mgr55__std__oob_type            ;
 assign    std__pe55__oob_data    =    mgr55__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe56__oob_cntl    =    mgr56__std__oob_cntl            ;
 assign    std__pe56__oob_valid   =    mgr56__std__oob_valid           ;
 assign    std__mgr56__oob_ready  =    pe56__std__oob_ready            ;
 assign    std__pe56__oob_type    =    mgr56__std__oob_type            ;
 assign    std__pe56__oob_data    =    mgr56__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe57__oob_cntl    =    mgr57__std__oob_cntl            ;
 assign    std__pe57__oob_valid   =    mgr57__std__oob_valid           ;
 assign    std__mgr57__oob_ready  =    pe57__std__oob_ready            ;
 assign    std__pe57__oob_type    =    mgr57__std__oob_type            ;
 assign    std__pe57__oob_data    =    mgr57__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe58__oob_cntl    =    mgr58__std__oob_cntl            ;
 assign    std__pe58__oob_valid   =    mgr58__std__oob_valid           ;
 assign    std__mgr58__oob_ready  =    pe58__std__oob_ready            ;
 assign    std__pe58__oob_type    =    mgr58__std__oob_type            ;
 assign    std__pe58__oob_data    =    mgr58__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe59__oob_cntl    =    mgr59__std__oob_cntl            ;
 assign    std__pe59__oob_valid   =    mgr59__std__oob_valid           ;
 assign    std__mgr59__oob_ready  =    pe59__std__oob_ready            ;
 assign    std__pe59__oob_type    =    mgr59__std__oob_type            ;
 assign    std__pe59__oob_data    =    mgr59__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe60__oob_cntl    =    mgr60__std__oob_cntl            ;
 assign    std__pe60__oob_valid   =    mgr60__std__oob_valid           ;
 assign    std__mgr60__oob_ready  =    pe60__std__oob_ready            ;
 assign    std__pe60__oob_type    =    mgr60__std__oob_type            ;
 assign    std__pe60__oob_data    =    mgr60__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe61__oob_cntl    =    mgr61__std__oob_cntl            ;
 assign    std__pe61__oob_valid   =    mgr61__std__oob_valid           ;
 assign    std__mgr61__oob_ready  =    pe61__std__oob_ready            ;
 assign    std__pe61__oob_type    =    mgr61__std__oob_type            ;
 assign    std__pe61__oob_data    =    mgr61__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe62__oob_cntl    =    mgr62__std__oob_cntl            ;
 assign    std__pe62__oob_valid   =    mgr62__std__oob_valid           ;
 assign    std__mgr62__oob_ready  =    pe62__std__oob_ready            ;
 assign    std__pe62__oob_type    =    mgr62__std__oob_type            ;
 assign    std__pe62__oob_data    =    mgr62__std__oob_data            ;

  // OOB controls how the lanes are interpreted                                  
 assign    std__pe63__oob_cntl    =    mgr63__std__oob_cntl            ;
 assign    std__pe63__oob_valid   =    mgr63__std__oob_valid           ;
 assign    std__mgr63__oob_ready  =    pe63__std__oob_ready            ;
 assign    std__pe63__oob_type    =    mgr63__std__oob_type            ;
 assign    std__pe63__oob_data    =    mgr63__std__oob_data            ;
