
                // Stream 2                 
                .dma__memc__write_valid2       ( 1'd0  ),
                .dma__memc__write_address2     (17'd0  ),
                .dma__memc__write_data2        (32'd0  ),
                .memc__dma__write_ready2       (  ),
                .dma__memc__read_valid2        ( 1'd0  ),
                .dma__memc__read_address2      (17'd0  ),
                .memc__dma__read_data2         (  ),
                .memc__dma__read_data_valid2   (  ),
                .memc__dma__read_ready2        (  ),
                .dma__memc__read_pause2        ( 1'd0  ),
                // Stream 3                 
                .dma__memc__write_valid3       ( 1'd0  ),
                .dma__memc__write_address3     (17'd0  ),
                .dma__memc__write_data3        (32'd0  ),
                .memc__dma__write_ready3       (  ),
                .dma__memc__read_valid3        ( 1'd0  ),
                .dma__memc__read_address3      (17'd0  ),
                .memc__dma__read_data3         (  ),
                .memc__dma__read_data_valid3   (  ),
                .memc__dma__read_ready3        (  ),
                .dma__memc__read_pause3        ( 1'd0  ),
                // Stream 4                 
                .dma__memc__write_valid4       ( 1'd0  ),
                .dma__memc__write_address4     (17'd0  ),
                .dma__memc__write_data4        (32'd0  ),
                .memc__dma__write_ready4       (  ),
                .dma__memc__read_valid4        ( 1'd0  ),
                .dma__memc__read_address4      (17'd0  ),
                .memc__dma__read_data4         (  ),
                .memc__dma__read_data_valid4   (  ),
                .memc__dma__read_ready4        (  ),
                .dma__memc__read_pause4        ( 1'd0  ),
                // Stream 5                 
                .dma__memc__write_valid5       ( 1'd0  ),
                .dma__memc__write_address5     (17'd0  ),
                .dma__memc__write_data5        (32'd0  ),
                .memc__dma__write_ready5       (  ),
                .dma__memc__read_valid5        ( 1'd0  ),
                .dma__memc__read_address5      (17'd0  ),
                .memc__dma__read_data5         (  ),
                .memc__dma__read_data_valid5   (  ),
                .memc__dma__read_ready5        (  ),
                .dma__memc__read_pause5        ( 1'd0  ),
                // Stream 6                 
                .dma__memc__write_valid6       ( 1'd0  ),
                .dma__memc__write_address6     (17'd0  ),
                .dma__memc__write_data6        (32'd0  ),
                .memc__dma__write_ready6       (  ),
                .dma__memc__read_valid6        ( 1'd0  ),
                .dma__memc__read_address6      (17'd0  ),
                .memc__dma__read_data6         (  ),
                .memc__dma__read_data_valid6   (  ),
                .memc__dma__read_ready6        (  ),
                .dma__memc__read_pause6        ( 1'd0  ),
                // Stream 7                 
                .dma__memc__write_valid7       ( 1'd0  ),
                .dma__memc__write_address7     (17'd0  ),
                .dma__memc__write_data7        (32'd0  ),
                .memc__dma__write_ready7       (  ),
                .dma__memc__read_valid7        ( 1'd0  ),
                .dma__memc__read_address7      (17'd0  ),
                .memc__dma__read_data7         (  ),
                .memc__dma__read_data_valid7   (  ),
                .memc__dma__read_ready7        (  ),
                .dma__memc__read_pause7        ( 1'd0  ),
                // Stream 8                 
                .dma__memc__write_valid8       ( 1'd0  ),
                .dma__memc__write_address8     (17'd0  ),
                .dma__memc__write_data8        (32'd0  ),
                .memc__dma__write_ready8       (  ),
                .dma__memc__read_valid8        ( 1'd0  ),
                .dma__memc__read_address8      (17'd0  ),
                .memc__dma__read_data8         (  ),
                .memc__dma__read_data_valid8   (  ),
                .memc__dma__read_ready8        (  ),
                .dma__memc__read_pause8        ( 1'd0  ),
                // Stream 9                 
                .dma__memc__write_valid9       ( 1'd0  ),
                .dma__memc__write_address9     (17'd0  ),
                .dma__memc__write_data9        (32'd0  ),
                .memc__dma__write_ready9       (  ),
                .dma__memc__read_valid9        ( 1'd0  ),
                .dma__memc__read_address9      (17'd0  ),
                .memc__dma__read_data9         (  ),
                .memc__dma__read_data_valid9   (  ),
                .memc__dma__read_ready9        (  ),
                .dma__memc__read_pause9        ( 1'd0  ),
                // Stream 10                 
                .dma__memc__write_valid10       ( 1'd0  ),
                .dma__memc__write_address10     (17'd0  ),
                .dma__memc__write_data10        (32'd0  ),
                .memc__dma__write_ready10       (  ),
                .dma__memc__read_valid10        ( 1'd0  ),
                .dma__memc__read_address10      (17'd0  ),
                .memc__dma__read_data10         (  ),
                .memc__dma__read_data_valid10   (  ),
                .memc__dma__read_ready10        (  ),
                .dma__memc__read_pause10        ( 1'd0  ),
                // Stream 11                 
                .dma__memc__write_valid11       ( 1'd0  ),
                .dma__memc__write_address11     (17'd0  ),
                .dma__memc__write_data11        (32'd0  ),
                .memc__dma__write_ready11       (  ),
                .dma__memc__read_valid11        ( 1'd0  ),
                .dma__memc__read_address11      (17'd0  ),
                .memc__dma__read_data11         (  ),
                .memc__dma__read_data_valid11   (  ),
                .memc__dma__read_ready11        (  ),
                .dma__memc__read_pause11        ( 1'd0  ),
                // Stream 12                 
                .dma__memc__write_valid12       ( 1'd0  ),
                .dma__memc__write_address12     (17'd0  ),
                .dma__memc__write_data12        (32'd0  ),
                .memc__dma__write_ready12       (  ),
                .dma__memc__read_valid12        ( 1'd0  ),
                .dma__memc__read_address12      (17'd0  ),
                .memc__dma__read_data12         (  ),
                .memc__dma__read_data_valid12   (  ),
                .memc__dma__read_ready12        (  ),
                .dma__memc__read_pause12        ( 1'd0  ),
                // Stream 13                 
                .dma__memc__write_valid13       ( 1'd0  ),
                .dma__memc__write_address13     (17'd0  ),
                .dma__memc__write_data13        (32'd0  ),
                .memc__dma__write_ready13       (  ),
                .dma__memc__read_valid13        ( 1'd0  ),
                .dma__memc__read_address13      (17'd0  ),
                .memc__dma__read_data13         (  ),
                .memc__dma__read_data_valid13   (  ),
                .memc__dma__read_ready13        (  ),
                .dma__memc__read_pause13        ( 1'd0  ),
                // Stream 14                 
                .dma__memc__write_valid14       ( 1'd0  ),
                .dma__memc__write_address14     (17'd0  ),
                .dma__memc__write_data14        (32'd0  ),
                .memc__dma__write_ready14       (  ),
                .dma__memc__read_valid14        ( 1'd0  ),
                .dma__memc__read_address14      (17'd0  ),
                .memc__dma__read_data14         (  ),
                .memc__dma__read_data_valid14   (  ),
                .memc__dma__read_ready14        (  ),
                .dma__memc__read_pause14        ( 1'd0  ),
                // Stream 15                 
                .dma__memc__write_valid15       ( 1'd0  ),
                .dma__memc__write_address15     (17'd0  ),
                .dma__memc__write_data15        (32'd0  ),
                .memc__dma__write_ready15       (  ),
                .dma__memc__read_valid15        ( 1'd0  ),
                .dma__memc__read_address15      (17'd0  ),
                .memc__dma__read_data15         (  ),
                .memc__dma__read_data_valid15   (  ),
                .memc__dma__read_ready15        (  ),
                .dma__memc__read_pause15        ( 1'd0  ),
                // Stream 16                 
                .dma__memc__write_valid16       ( 1'd0  ),
                .dma__memc__write_address16     (17'd0  ),
                .dma__memc__write_data16        (32'd0  ),
                .memc__dma__write_ready16       (  ),
                .dma__memc__read_valid16        ( 1'd0  ),
                .dma__memc__read_address16      (17'd0  ),
                .memc__dma__read_data16         (  ),
                .memc__dma__read_data_valid16   (  ),
                .memc__dma__read_ready16        (  ),
                .dma__memc__read_pause16        ( 1'd0  ),
                // Stream 17                 
                .dma__memc__write_valid17       ( 1'd0  ),
                .dma__memc__write_address17     (17'd0  ),
                .dma__memc__write_data17        (32'd0  ),
                .memc__dma__write_ready17       (  ),
                .dma__memc__read_valid17        ( 1'd0  ),
                .dma__memc__read_address17      (17'd0  ),
                .memc__dma__read_data17         (  ),
                .memc__dma__read_data_valid17   (  ),
                .memc__dma__read_ready17        (  ),
                .dma__memc__read_pause17        ( 1'd0  ),
                // Stream 18                 
                .dma__memc__write_valid18       ( 1'd0  ),
                .dma__memc__write_address18     (17'd0  ),
                .dma__memc__write_data18        (32'd0  ),
                .memc__dma__write_ready18       (  ),
                .dma__memc__read_valid18        ( 1'd0  ),
                .dma__memc__read_address18      (17'd0  ),
                .memc__dma__read_data18         (  ),
                .memc__dma__read_data_valid18   (  ),
                .memc__dma__read_ready18        (  ),
                .dma__memc__read_pause18        ( 1'd0  ),
                // Stream 19                 
                .dma__memc__write_valid19       ( 1'd0  ),
                .dma__memc__write_address19     (17'd0  ),
                .dma__memc__write_data19        (32'd0  ),
                .memc__dma__write_ready19       (  ),
                .dma__memc__read_valid19        ( 1'd0  ),
                .dma__memc__read_address19      (17'd0  ),
                .memc__dma__read_data19         (  ),
                .memc__dma__read_data_valid19   (  ),
                .memc__dma__read_ready19        (  ),
                .dma__memc__read_pause19        ( 1'd0  ),
                // Stream 20                 
                .dma__memc__write_valid20       ( 1'd0  ),
                .dma__memc__write_address20     (17'd0  ),
                .dma__memc__write_data20        (32'd0  ),
                .memc__dma__write_ready20       (  ),
                .dma__memc__read_valid20        ( 1'd0  ),
                .dma__memc__read_address20      (17'd0  ),
                .memc__dma__read_data20         (  ),
                .memc__dma__read_data_valid20   (  ),
                .memc__dma__read_ready20        (  ),
                .dma__memc__read_pause20        ( 1'd0  ),
                // Stream 21                 
                .dma__memc__write_valid21       ( 1'd0  ),
                .dma__memc__write_address21     (17'd0  ),
                .dma__memc__write_data21        (32'd0  ),
                .memc__dma__write_ready21       (  ),
                .dma__memc__read_valid21        ( 1'd0  ),
                .dma__memc__read_address21      (17'd0  ),
                .memc__dma__read_data21         (  ),
                .memc__dma__read_data_valid21   (  ),
                .memc__dma__read_ready21        (  ),
                .dma__memc__read_pause21        ( 1'd0  ),
                // Stream 22                 
                .dma__memc__write_valid22       ( 1'd0  ),
                .dma__memc__write_address22     (17'd0  ),
                .dma__memc__write_data22        (32'd0  ),
                .memc__dma__write_ready22       (  ),
                .dma__memc__read_valid22        ( 1'd0  ),
                .dma__memc__read_address22      (17'd0  ),
                .memc__dma__read_data22         (  ),
                .memc__dma__read_data_valid22   (  ),
                .memc__dma__read_ready22        (  ),
                .dma__memc__read_pause22        ( 1'd0  ),
                // Stream 23                 
                .dma__memc__write_valid23       ( 1'd0  ),
                .dma__memc__write_address23     (17'd0  ),
                .dma__memc__write_data23        (32'd0  ),
                .memc__dma__write_ready23       (  ),
                .dma__memc__read_valid23        ( 1'd0  ),
                .dma__memc__read_address23      (17'd0  ),
                .memc__dma__read_data23         (  ),
                .memc__dma__read_data_valid23   (  ),
                .memc__dma__read_ready23        (  ),
                .dma__memc__read_pause23        ( 1'd0  ),
                // Stream 24                 
                .dma__memc__write_valid24       ( 1'd0  ),
                .dma__memc__write_address24     (17'd0  ),
                .dma__memc__write_data24        (32'd0  ),
                .memc__dma__write_ready24       (  ),
                .dma__memc__read_valid24        ( 1'd0  ),
                .dma__memc__read_address24      (17'd0  ),
                .memc__dma__read_data24         (  ),
                .memc__dma__read_data_valid24   (  ),
                .memc__dma__read_ready24        (  ),
                .dma__memc__read_pause24        ( 1'd0  ),
                // Stream 25                 
                .dma__memc__write_valid25       ( 1'd0  ),
                .dma__memc__write_address25     (17'd0  ),
                .dma__memc__write_data25        (32'd0  ),
                .memc__dma__write_ready25       (  ),
                .dma__memc__read_valid25        ( 1'd0  ),
                .dma__memc__read_address25      (17'd0  ),
                .memc__dma__read_data25         (  ),
                .memc__dma__read_data_valid25   (  ),
                .memc__dma__read_ready25        (  ),
                .dma__memc__read_pause25        ( 1'd0  ),
                // Stream 26                 
                .dma__memc__write_valid26       ( 1'd0  ),
                .dma__memc__write_address26     (17'd0  ),
                .dma__memc__write_data26        (32'd0  ),
                .memc__dma__write_ready26       (  ),
                .dma__memc__read_valid26        ( 1'd0  ),
                .dma__memc__read_address26      (17'd0  ),
                .memc__dma__read_data26         (  ),
                .memc__dma__read_data_valid26   (  ),
                .memc__dma__read_ready26        (  ),
                .dma__memc__read_pause26        ( 1'd0  ),
                // Stream 27                 
                .dma__memc__write_valid27       ( 1'd0  ),
                .dma__memc__write_address27     (17'd0  ),
                .dma__memc__write_data27        (32'd0  ),
                .memc__dma__write_ready27       (  ),
                .dma__memc__read_valid27        ( 1'd0  ),
                .dma__memc__read_address27      (17'd0  ),
                .memc__dma__read_data27         (  ),
                .memc__dma__read_data_valid27   (  ),
                .memc__dma__read_ready27        (  ),
                .dma__memc__read_pause27        ( 1'd0  ),
                // Stream 28                 
                .dma__memc__write_valid28       ( 1'd0  ),
                .dma__memc__write_address28     (17'd0  ),
                .dma__memc__write_data28        (32'd0  ),
                .memc__dma__write_ready28       (  ),
                .dma__memc__read_valid28        ( 1'd0  ),
                .dma__memc__read_address28      (17'd0  ),
                .memc__dma__read_data28         (  ),
                .memc__dma__read_data_valid28   (  ),
                .memc__dma__read_ready28        (  ),
                .dma__memc__read_pause28        ( 1'd0  ),
                // Stream 29                 
                .dma__memc__write_valid29       ( 1'd0  ),
                .dma__memc__write_address29     (17'd0  ),
                .dma__memc__write_data29        (32'd0  ),
                .memc__dma__write_ready29       (  ),
                .dma__memc__read_valid29        ( 1'd0  ),
                .dma__memc__read_address29      (17'd0  ),
                .memc__dma__read_data29         (  ),
                .memc__dma__read_data_valid29   (  ),
                .memc__dma__read_ready29        (  ),
                .dma__memc__read_pause29        ( 1'd0  ),
                // Stream 30                 
                .dma__memc__write_valid30       ( 1'd0  ),
                .dma__memc__write_address30     (17'd0  ),
                .dma__memc__write_data30        (32'd0  ),
                .memc__dma__write_ready30       (  ),
                .dma__memc__read_valid30        ( 1'd0  ),
                .dma__memc__read_address30      (17'd0  ),
                .memc__dma__read_data30         (  ),
                .memc__dma__read_data_valid30   (  ),
                .memc__dma__read_ready30        (  ),
                .dma__memc__read_pause30        ( 1'd0  ),
                // Stream 31                 
                .dma__memc__write_valid31       ( 1'd0  ),
                .dma__memc__write_address31     (17'd0  ),
                .dma__memc__write_data31        (32'd0  ),
                .memc__dma__write_ready31       (  ),
                .dma__memc__read_valid31        ( 1'd0  ),
                .dma__memc__read_address31      (17'd0  ),
                .memc__dma__read_data31         (  ),
                .memc__dma__read_data_valid31   (  ),
                .memc__dma__read_ready31        (  ),
                .dma__memc__read_pause31        ( 1'd0  ),