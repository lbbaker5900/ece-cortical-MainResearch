
    .reg__sdp__lane0_ready    ( reg__sdp__lane0_ready  ),
    .sdp__reg__lane0_valid    ( sdp__reg__lane0_valid  ),
    .sdp__reg__lane0_data     ( sdp__reg__lane0_data   ),

    .reg__sdp__lane1_ready    ( reg__sdp__lane1_ready  ),
    .sdp__reg__lane1_valid    ( sdp__reg__lane1_valid  ),
    .sdp__reg__lane1_data     ( sdp__reg__lane1_data   ),

    .reg__sdp__lane2_ready    ( reg__sdp__lane2_ready  ),
    .sdp__reg__lane2_valid    ( sdp__reg__lane2_valid  ),
    .sdp__reg__lane2_data     ( sdp__reg__lane2_data   ),

    .reg__sdp__lane3_ready    ( reg__sdp__lane3_ready  ),
    .sdp__reg__lane3_valid    ( sdp__reg__lane3_valid  ),
    .sdp__reg__lane3_data     ( sdp__reg__lane3_data   ),

    .reg__sdp__lane4_ready    ( reg__sdp__lane4_ready  ),
    .sdp__reg__lane4_valid    ( sdp__reg__lane4_valid  ),
    .sdp__reg__lane4_data     ( sdp__reg__lane4_data   ),

    .reg__sdp__lane5_ready    ( reg__sdp__lane5_ready  ),
    .sdp__reg__lane5_valid    ( sdp__reg__lane5_valid  ),
    .sdp__reg__lane5_data     ( sdp__reg__lane5_data   ),

    .reg__sdp__lane6_ready    ( reg__sdp__lane6_ready  ),
    .sdp__reg__lane6_valid    ( sdp__reg__lane6_valid  ),
    .sdp__reg__lane6_data     ( sdp__reg__lane6_data   ),

    .reg__sdp__lane7_ready    ( reg__sdp__lane7_ready  ),
    .sdp__reg__lane7_valid    ( sdp__reg__lane7_valid  ),
    .sdp__reg__lane7_data     ( sdp__reg__lane7_data   ),

    .reg__sdp__lane8_ready    ( reg__sdp__lane8_ready  ),
    .sdp__reg__lane8_valid    ( sdp__reg__lane8_valid  ),
    .sdp__reg__lane8_data     ( sdp__reg__lane8_data   ),

    .reg__sdp__lane9_ready    ( reg__sdp__lane9_ready  ),
    .sdp__reg__lane9_valid    ( sdp__reg__lane9_valid  ),
    .sdp__reg__lane9_data     ( sdp__reg__lane9_data   ),

    .reg__sdp__lane10_ready    ( reg__sdp__lane10_ready  ),
    .sdp__reg__lane10_valid    ( sdp__reg__lane10_valid  ),
    .sdp__reg__lane10_data     ( sdp__reg__lane10_data   ),

    .reg__sdp__lane11_ready    ( reg__sdp__lane11_ready  ),
    .sdp__reg__lane11_valid    ( sdp__reg__lane11_valid  ),
    .sdp__reg__lane11_data     ( sdp__reg__lane11_data   ),

    .reg__sdp__lane12_ready    ( reg__sdp__lane12_ready  ),
    .sdp__reg__lane12_valid    ( sdp__reg__lane12_valid  ),
    .sdp__reg__lane12_data     ( sdp__reg__lane12_data   ),

    .reg__sdp__lane13_ready    ( reg__sdp__lane13_ready  ),
    .sdp__reg__lane13_valid    ( sdp__reg__lane13_valid  ),
    .sdp__reg__lane13_data     ( sdp__reg__lane13_data   ),

    .reg__sdp__lane14_ready    ( reg__sdp__lane14_ready  ),
    .sdp__reg__lane14_valid    ( sdp__reg__lane14_valid  ),
    .sdp__reg__lane14_data     ( sdp__reg__lane14_data   ),

    .reg__sdp__lane15_ready    ( reg__sdp__lane15_ready  ),
    .sdp__reg__lane15_valid    ( sdp__reg__lane15_valid  ),
    .sdp__reg__lane15_data     ( sdp__reg__lane15_data   ),

    .reg__sdp__lane16_ready    ( reg__sdp__lane16_ready  ),
    .sdp__reg__lane16_valid    ( sdp__reg__lane16_valid  ),
    .sdp__reg__lane16_data     ( sdp__reg__lane16_data   ),

    .reg__sdp__lane17_ready    ( reg__sdp__lane17_ready  ),
    .sdp__reg__lane17_valid    ( sdp__reg__lane17_valid  ),
    .sdp__reg__lane17_data     ( sdp__reg__lane17_data   ),

    .reg__sdp__lane18_ready    ( reg__sdp__lane18_ready  ),
    .sdp__reg__lane18_valid    ( sdp__reg__lane18_valid  ),
    .sdp__reg__lane18_data     ( sdp__reg__lane18_data   ),

    .reg__sdp__lane19_ready    ( reg__sdp__lane19_ready  ),
    .sdp__reg__lane19_valid    ( sdp__reg__lane19_valid  ),
    .sdp__reg__lane19_data     ( sdp__reg__lane19_data   ),

    .reg__sdp__lane20_ready    ( reg__sdp__lane20_ready  ),
    .sdp__reg__lane20_valid    ( sdp__reg__lane20_valid  ),
    .sdp__reg__lane20_data     ( sdp__reg__lane20_data   ),

    .reg__sdp__lane21_ready    ( reg__sdp__lane21_ready  ),
    .sdp__reg__lane21_valid    ( sdp__reg__lane21_valid  ),
    .sdp__reg__lane21_data     ( sdp__reg__lane21_data   ),

    .reg__sdp__lane22_ready    ( reg__sdp__lane22_ready  ),
    .sdp__reg__lane22_valid    ( sdp__reg__lane22_valid  ),
    .sdp__reg__lane22_data     ( sdp__reg__lane22_data   ),

    .reg__sdp__lane23_ready    ( reg__sdp__lane23_ready  ),
    .sdp__reg__lane23_valid    ( sdp__reg__lane23_valid  ),
    .sdp__reg__lane23_data     ( sdp__reg__lane23_data   ),

    .reg__sdp__lane24_ready    ( reg__sdp__lane24_ready  ),
    .sdp__reg__lane24_valid    ( sdp__reg__lane24_valid  ),
    .sdp__reg__lane24_data     ( sdp__reg__lane24_data   ),

    .reg__sdp__lane25_ready    ( reg__sdp__lane25_ready  ),
    .sdp__reg__lane25_valid    ( sdp__reg__lane25_valid  ),
    .sdp__reg__lane25_data     ( sdp__reg__lane25_data   ),

    .reg__sdp__lane26_ready    ( reg__sdp__lane26_ready  ),
    .sdp__reg__lane26_valid    ( sdp__reg__lane26_valid  ),
    .sdp__reg__lane26_data     ( sdp__reg__lane26_data   ),

    .reg__sdp__lane27_ready    ( reg__sdp__lane27_ready  ),
    .sdp__reg__lane27_valid    ( sdp__reg__lane27_valid  ),
    .sdp__reg__lane27_data     ( sdp__reg__lane27_data   ),

    .reg__sdp__lane28_ready    ( reg__sdp__lane28_ready  ),
    .sdp__reg__lane28_valid    ( sdp__reg__lane28_valid  ),
    .sdp__reg__lane28_data     ( sdp__reg__lane28_data   ),

    .reg__sdp__lane29_ready    ( reg__sdp__lane29_ready  ),
    .sdp__reg__lane29_valid    ( sdp__reg__lane29_valid  ),
    .sdp__reg__lane29_data     ( sdp__reg__lane29_data   ),

    .reg__sdp__lane30_ready    ( reg__sdp__lane30_ready  ),
    .sdp__reg__lane30_valid    ( sdp__reg__lane30_valid  ),
    .sdp__reg__lane30_data     ( sdp__reg__lane30_data   ),

    .reg__sdp__lane31_ready    ( reg__sdp__lane31_ready  ),
    .sdp__reg__lane31_valid    ( sdp__reg__lane31_valid  ),
    .sdp__reg__lane31_data     ( sdp__reg__lane31_data   ),

