
  assign   mgr_inst[0].stu__mgr__valid     =   stu__mgr0__valid               ;
  assign   mgr_inst[0].stu__mgr__cntl      =   stu__mgr0__cntl                ;
  assign   mgr__stu0__ready                =   mgr_inst[0].mgr__stu__ready    ;
  assign   mgr_inst[0].stu__mgr__type      =   stu__mgr0__type                ;
  assign   mgr_inst[0].stu__mgr__data      =   stu__mgr0__data                ;
  assign   mgr_inst[0].stu__mgr__oob_data  =   stu__mgr0__oob_data            ;

  assign   mgr_inst[1].stu__mgr__valid     =   stu__mgr1__valid               ;
  assign   mgr_inst[1].stu__mgr__cntl      =   stu__mgr1__cntl                ;
  assign   mgr__stu1__ready                =   mgr_inst[1].mgr__stu__ready    ;
  assign   mgr_inst[1].stu__mgr__type      =   stu__mgr1__type                ;
  assign   mgr_inst[1].stu__mgr__data      =   stu__mgr1__data                ;
  assign   mgr_inst[1].stu__mgr__oob_data  =   stu__mgr1__oob_data            ;

  assign   mgr_inst[2].stu__mgr__valid     =   stu__mgr2__valid               ;
  assign   mgr_inst[2].stu__mgr__cntl      =   stu__mgr2__cntl                ;
  assign   mgr__stu2__ready                =   mgr_inst[2].mgr__stu__ready    ;
  assign   mgr_inst[2].stu__mgr__type      =   stu__mgr2__type                ;
  assign   mgr_inst[2].stu__mgr__data      =   stu__mgr2__data                ;
  assign   mgr_inst[2].stu__mgr__oob_data  =   stu__mgr2__oob_data            ;

  assign   mgr_inst[3].stu__mgr__valid     =   stu__mgr3__valid               ;
  assign   mgr_inst[3].stu__mgr__cntl      =   stu__mgr3__cntl                ;
  assign   mgr__stu3__ready                =   mgr_inst[3].mgr__stu__ready    ;
  assign   mgr_inst[3].stu__mgr__type      =   stu__mgr3__type                ;
  assign   mgr_inst[3].stu__mgr__data      =   stu__mgr3__data                ;
  assign   mgr_inst[3].stu__mgr__oob_data  =   stu__mgr3__oob_data            ;

  assign   mgr_inst[4].stu__mgr__valid     =   stu__mgr4__valid               ;
  assign   mgr_inst[4].stu__mgr__cntl      =   stu__mgr4__cntl                ;
  assign   mgr__stu4__ready                =   mgr_inst[4].mgr__stu__ready    ;
  assign   mgr_inst[4].stu__mgr__type      =   stu__mgr4__type                ;
  assign   mgr_inst[4].stu__mgr__data      =   stu__mgr4__data                ;
  assign   mgr_inst[4].stu__mgr__oob_data  =   stu__mgr4__oob_data            ;

  assign   mgr_inst[5].stu__mgr__valid     =   stu__mgr5__valid               ;
  assign   mgr_inst[5].stu__mgr__cntl      =   stu__mgr5__cntl                ;
  assign   mgr__stu5__ready                =   mgr_inst[5].mgr__stu__ready    ;
  assign   mgr_inst[5].stu__mgr__type      =   stu__mgr5__type                ;
  assign   mgr_inst[5].stu__mgr__data      =   stu__mgr5__data                ;
  assign   mgr_inst[5].stu__mgr__oob_data  =   stu__mgr5__oob_data            ;

  assign   mgr_inst[6].stu__mgr__valid     =   stu__mgr6__valid               ;
  assign   mgr_inst[6].stu__mgr__cntl      =   stu__mgr6__cntl                ;
  assign   mgr__stu6__ready                =   mgr_inst[6].mgr__stu__ready    ;
  assign   mgr_inst[6].stu__mgr__type      =   stu__mgr6__type                ;
  assign   mgr_inst[6].stu__mgr__data      =   stu__mgr6__data                ;
  assign   mgr_inst[6].stu__mgr__oob_data  =   stu__mgr6__oob_data            ;

  assign   mgr_inst[7].stu__mgr__valid     =   stu__mgr7__valid               ;
  assign   mgr_inst[7].stu__mgr__cntl      =   stu__mgr7__cntl                ;
  assign   mgr__stu7__ready                =   mgr_inst[7].mgr__stu__ready    ;
  assign   mgr_inst[7].stu__mgr__type      =   stu__mgr7__type                ;
  assign   mgr_inst[7].stu__mgr__data      =   stu__mgr7__data                ;
  assign   mgr_inst[7].stu__mgr__oob_data  =   stu__mgr7__oob_data            ;

  assign   mgr_inst[8].stu__mgr__valid     =   stu__mgr8__valid               ;
  assign   mgr_inst[8].stu__mgr__cntl      =   stu__mgr8__cntl                ;
  assign   mgr__stu8__ready                =   mgr_inst[8].mgr__stu__ready    ;
  assign   mgr_inst[8].stu__mgr__type      =   stu__mgr8__type                ;
  assign   mgr_inst[8].stu__mgr__data      =   stu__mgr8__data                ;
  assign   mgr_inst[8].stu__mgr__oob_data  =   stu__mgr8__oob_data            ;

  assign   mgr_inst[9].stu__mgr__valid     =   stu__mgr9__valid               ;
  assign   mgr_inst[9].stu__mgr__cntl      =   stu__mgr9__cntl                ;
  assign   mgr__stu9__ready                =   mgr_inst[9].mgr__stu__ready    ;
  assign   mgr_inst[9].stu__mgr__type      =   stu__mgr9__type                ;
  assign   mgr_inst[9].stu__mgr__data      =   stu__mgr9__data                ;
  assign   mgr_inst[9].stu__mgr__oob_data  =   stu__mgr9__oob_data            ;

  assign   mgr_inst[10].stu__mgr__valid     =   stu__mgr10__valid               ;
  assign   mgr_inst[10].stu__mgr__cntl      =   stu__mgr10__cntl                ;
  assign   mgr__stu10__ready                =   mgr_inst[10].mgr__stu__ready    ;
  assign   mgr_inst[10].stu__mgr__type      =   stu__mgr10__type                ;
  assign   mgr_inst[10].stu__mgr__data      =   stu__mgr10__data                ;
  assign   mgr_inst[10].stu__mgr__oob_data  =   stu__mgr10__oob_data            ;

  assign   mgr_inst[11].stu__mgr__valid     =   stu__mgr11__valid               ;
  assign   mgr_inst[11].stu__mgr__cntl      =   stu__mgr11__cntl                ;
  assign   mgr__stu11__ready                =   mgr_inst[11].mgr__stu__ready    ;
  assign   mgr_inst[11].stu__mgr__type      =   stu__mgr11__type                ;
  assign   mgr_inst[11].stu__mgr__data      =   stu__mgr11__data                ;
  assign   mgr_inst[11].stu__mgr__oob_data  =   stu__mgr11__oob_data            ;

  assign   mgr_inst[12].stu__mgr__valid     =   stu__mgr12__valid               ;
  assign   mgr_inst[12].stu__mgr__cntl      =   stu__mgr12__cntl                ;
  assign   mgr__stu12__ready                =   mgr_inst[12].mgr__stu__ready    ;
  assign   mgr_inst[12].stu__mgr__type      =   stu__mgr12__type                ;
  assign   mgr_inst[12].stu__mgr__data      =   stu__mgr12__data                ;
  assign   mgr_inst[12].stu__mgr__oob_data  =   stu__mgr12__oob_data            ;

  assign   mgr_inst[13].stu__mgr__valid     =   stu__mgr13__valid               ;
  assign   mgr_inst[13].stu__mgr__cntl      =   stu__mgr13__cntl                ;
  assign   mgr__stu13__ready                =   mgr_inst[13].mgr__stu__ready    ;
  assign   mgr_inst[13].stu__mgr__type      =   stu__mgr13__type                ;
  assign   mgr_inst[13].stu__mgr__data      =   stu__mgr13__data                ;
  assign   mgr_inst[13].stu__mgr__oob_data  =   stu__mgr13__oob_data            ;

  assign   mgr_inst[14].stu__mgr__valid     =   stu__mgr14__valid               ;
  assign   mgr_inst[14].stu__mgr__cntl      =   stu__mgr14__cntl                ;
  assign   mgr__stu14__ready                =   mgr_inst[14].mgr__stu__ready    ;
  assign   mgr_inst[14].stu__mgr__type      =   stu__mgr14__type                ;
  assign   mgr_inst[14].stu__mgr__data      =   stu__mgr14__data                ;
  assign   mgr_inst[14].stu__mgr__oob_data  =   stu__mgr14__oob_data            ;

  assign   mgr_inst[15].stu__mgr__valid     =   stu__mgr15__valid               ;
  assign   mgr_inst[15].stu__mgr__cntl      =   stu__mgr15__cntl                ;
  assign   mgr__stu15__ready                =   mgr_inst[15].mgr__stu__ready    ;
  assign   mgr_inst[15].stu__mgr__type      =   stu__mgr15__type                ;
  assign   mgr_inst[15].stu__mgr__data      =   stu__mgr15__data                ;
  assign   mgr_inst[15].stu__mgr__oob_data  =   stu__mgr15__oob_data            ;

  assign   mgr_inst[16].stu__mgr__valid     =   stu__mgr16__valid               ;
  assign   mgr_inst[16].stu__mgr__cntl      =   stu__mgr16__cntl                ;
  assign   mgr__stu16__ready                =   mgr_inst[16].mgr__stu__ready    ;
  assign   mgr_inst[16].stu__mgr__type      =   stu__mgr16__type                ;
  assign   mgr_inst[16].stu__mgr__data      =   stu__mgr16__data                ;
  assign   mgr_inst[16].stu__mgr__oob_data  =   stu__mgr16__oob_data            ;

  assign   mgr_inst[17].stu__mgr__valid     =   stu__mgr17__valid               ;
  assign   mgr_inst[17].stu__mgr__cntl      =   stu__mgr17__cntl                ;
  assign   mgr__stu17__ready                =   mgr_inst[17].mgr__stu__ready    ;
  assign   mgr_inst[17].stu__mgr__type      =   stu__mgr17__type                ;
  assign   mgr_inst[17].stu__mgr__data      =   stu__mgr17__data                ;
  assign   mgr_inst[17].stu__mgr__oob_data  =   stu__mgr17__oob_data            ;

  assign   mgr_inst[18].stu__mgr__valid     =   stu__mgr18__valid               ;
  assign   mgr_inst[18].stu__mgr__cntl      =   stu__mgr18__cntl                ;
  assign   mgr__stu18__ready                =   mgr_inst[18].mgr__stu__ready    ;
  assign   mgr_inst[18].stu__mgr__type      =   stu__mgr18__type                ;
  assign   mgr_inst[18].stu__mgr__data      =   stu__mgr18__data                ;
  assign   mgr_inst[18].stu__mgr__oob_data  =   stu__mgr18__oob_data            ;

  assign   mgr_inst[19].stu__mgr__valid     =   stu__mgr19__valid               ;
  assign   mgr_inst[19].stu__mgr__cntl      =   stu__mgr19__cntl                ;
  assign   mgr__stu19__ready                =   mgr_inst[19].mgr__stu__ready    ;
  assign   mgr_inst[19].stu__mgr__type      =   stu__mgr19__type                ;
  assign   mgr_inst[19].stu__mgr__data      =   stu__mgr19__data                ;
  assign   mgr_inst[19].stu__mgr__oob_data  =   stu__mgr19__oob_data            ;

  assign   mgr_inst[20].stu__mgr__valid     =   stu__mgr20__valid               ;
  assign   mgr_inst[20].stu__mgr__cntl      =   stu__mgr20__cntl                ;
  assign   mgr__stu20__ready                =   mgr_inst[20].mgr__stu__ready    ;
  assign   mgr_inst[20].stu__mgr__type      =   stu__mgr20__type                ;
  assign   mgr_inst[20].stu__mgr__data      =   stu__mgr20__data                ;
  assign   mgr_inst[20].stu__mgr__oob_data  =   stu__mgr20__oob_data            ;

  assign   mgr_inst[21].stu__mgr__valid     =   stu__mgr21__valid               ;
  assign   mgr_inst[21].stu__mgr__cntl      =   stu__mgr21__cntl                ;
  assign   mgr__stu21__ready                =   mgr_inst[21].mgr__stu__ready    ;
  assign   mgr_inst[21].stu__mgr__type      =   stu__mgr21__type                ;
  assign   mgr_inst[21].stu__mgr__data      =   stu__mgr21__data                ;
  assign   mgr_inst[21].stu__mgr__oob_data  =   stu__mgr21__oob_data            ;

  assign   mgr_inst[22].stu__mgr__valid     =   stu__mgr22__valid               ;
  assign   mgr_inst[22].stu__mgr__cntl      =   stu__mgr22__cntl                ;
  assign   mgr__stu22__ready                =   mgr_inst[22].mgr__stu__ready    ;
  assign   mgr_inst[22].stu__mgr__type      =   stu__mgr22__type                ;
  assign   mgr_inst[22].stu__mgr__data      =   stu__mgr22__data                ;
  assign   mgr_inst[22].stu__mgr__oob_data  =   stu__mgr22__oob_data            ;

  assign   mgr_inst[23].stu__mgr__valid     =   stu__mgr23__valid               ;
  assign   mgr_inst[23].stu__mgr__cntl      =   stu__mgr23__cntl                ;
  assign   mgr__stu23__ready                =   mgr_inst[23].mgr__stu__ready    ;
  assign   mgr_inst[23].stu__mgr__type      =   stu__mgr23__type                ;
  assign   mgr_inst[23].stu__mgr__data      =   stu__mgr23__data                ;
  assign   mgr_inst[23].stu__mgr__oob_data  =   stu__mgr23__oob_data            ;

  assign   mgr_inst[24].stu__mgr__valid     =   stu__mgr24__valid               ;
  assign   mgr_inst[24].stu__mgr__cntl      =   stu__mgr24__cntl                ;
  assign   mgr__stu24__ready                =   mgr_inst[24].mgr__stu__ready    ;
  assign   mgr_inst[24].stu__mgr__type      =   stu__mgr24__type                ;
  assign   mgr_inst[24].stu__mgr__data      =   stu__mgr24__data                ;
  assign   mgr_inst[24].stu__mgr__oob_data  =   stu__mgr24__oob_data            ;

  assign   mgr_inst[25].stu__mgr__valid     =   stu__mgr25__valid               ;
  assign   mgr_inst[25].stu__mgr__cntl      =   stu__mgr25__cntl                ;
  assign   mgr__stu25__ready                =   mgr_inst[25].mgr__stu__ready    ;
  assign   mgr_inst[25].stu__mgr__type      =   stu__mgr25__type                ;
  assign   mgr_inst[25].stu__mgr__data      =   stu__mgr25__data                ;
  assign   mgr_inst[25].stu__mgr__oob_data  =   stu__mgr25__oob_data            ;

  assign   mgr_inst[26].stu__mgr__valid     =   stu__mgr26__valid               ;
  assign   mgr_inst[26].stu__mgr__cntl      =   stu__mgr26__cntl                ;
  assign   mgr__stu26__ready                =   mgr_inst[26].mgr__stu__ready    ;
  assign   mgr_inst[26].stu__mgr__type      =   stu__mgr26__type                ;
  assign   mgr_inst[26].stu__mgr__data      =   stu__mgr26__data                ;
  assign   mgr_inst[26].stu__mgr__oob_data  =   stu__mgr26__oob_data            ;

  assign   mgr_inst[27].stu__mgr__valid     =   stu__mgr27__valid               ;
  assign   mgr_inst[27].stu__mgr__cntl      =   stu__mgr27__cntl                ;
  assign   mgr__stu27__ready                =   mgr_inst[27].mgr__stu__ready    ;
  assign   mgr_inst[27].stu__mgr__type      =   stu__mgr27__type                ;
  assign   mgr_inst[27].stu__mgr__data      =   stu__mgr27__data                ;
  assign   mgr_inst[27].stu__mgr__oob_data  =   stu__mgr27__oob_data            ;

  assign   mgr_inst[28].stu__mgr__valid     =   stu__mgr28__valid               ;
  assign   mgr_inst[28].stu__mgr__cntl      =   stu__mgr28__cntl                ;
  assign   mgr__stu28__ready                =   mgr_inst[28].mgr__stu__ready    ;
  assign   mgr_inst[28].stu__mgr__type      =   stu__mgr28__type                ;
  assign   mgr_inst[28].stu__mgr__data      =   stu__mgr28__data                ;
  assign   mgr_inst[28].stu__mgr__oob_data  =   stu__mgr28__oob_data            ;

  assign   mgr_inst[29].stu__mgr__valid     =   stu__mgr29__valid               ;
  assign   mgr_inst[29].stu__mgr__cntl      =   stu__mgr29__cntl                ;
  assign   mgr__stu29__ready                =   mgr_inst[29].mgr__stu__ready    ;
  assign   mgr_inst[29].stu__mgr__type      =   stu__mgr29__type                ;
  assign   mgr_inst[29].stu__mgr__data      =   stu__mgr29__data                ;
  assign   mgr_inst[29].stu__mgr__oob_data  =   stu__mgr29__oob_data            ;

  assign   mgr_inst[30].stu__mgr__valid     =   stu__mgr30__valid               ;
  assign   mgr_inst[30].stu__mgr__cntl      =   stu__mgr30__cntl                ;
  assign   mgr__stu30__ready                =   mgr_inst[30].mgr__stu__ready    ;
  assign   mgr_inst[30].stu__mgr__type      =   stu__mgr30__type                ;
  assign   mgr_inst[30].stu__mgr__data      =   stu__mgr30__data                ;
  assign   mgr_inst[30].stu__mgr__oob_data  =   stu__mgr30__oob_data            ;

  assign   mgr_inst[31].stu__mgr__valid     =   stu__mgr31__valid               ;
  assign   mgr_inst[31].stu__mgr__cntl      =   stu__mgr31__cntl                ;
  assign   mgr__stu31__ready                =   mgr_inst[31].mgr__stu__ready    ;
  assign   mgr_inst[31].stu__mgr__type      =   stu__mgr31__type                ;
  assign   mgr_inst[31].stu__mgr__data      =   stu__mgr31__data                ;
  assign   mgr_inst[31].stu__mgr__oob_data  =   stu__mgr31__oob_data            ;

  assign   mgr_inst[32].stu__mgr__valid     =   stu__mgr32__valid               ;
  assign   mgr_inst[32].stu__mgr__cntl      =   stu__mgr32__cntl                ;
  assign   mgr__stu32__ready                =   mgr_inst[32].mgr__stu__ready    ;
  assign   mgr_inst[32].stu__mgr__type      =   stu__mgr32__type                ;
  assign   mgr_inst[32].stu__mgr__data      =   stu__mgr32__data                ;
  assign   mgr_inst[32].stu__mgr__oob_data  =   stu__mgr32__oob_data            ;

  assign   mgr_inst[33].stu__mgr__valid     =   stu__mgr33__valid               ;
  assign   mgr_inst[33].stu__mgr__cntl      =   stu__mgr33__cntl                ;
  assign   mgr__stu33__ready                =   mgr_inst[33].mgr__stu__ready    ;
  assign   mgr_inst[33].stu__mgr__type      =   stu__mgr33__type                ;
  assign   mgr_inst[33].stu__mgr__data      =   stu__mgr33__data                ;
  assign   mgr_inst[33].stu__mgr__oob_data  =   stu__mgr33__oob_data            ;

  assign   mgr_inst[34].stu__mgr__valid     =   stu__mgr34__valid               ;
  assign   mgr_inst[34].stu__mgr__cntl      =   stu__mgr34__cntl                ;
  assign   mgr__stu34__ready                =   mgr_inst[34].mgr__stu__ready    ;
  assign   mgr_inst[34].stu__mgr__type      =   stu__mgr34__type                ;
  assign   mgr_inst[34].stu__mgr__data      =   stu__mgr34__data                ;
  assign   mgr_inst[34].stu__mgr__oob_data  =   stu__mgr34__oob_data            ;

  assign   mgr_inst[35].stu__mgr__valid     =   stu__mgr35__valid               ;
  assign   mgr_inst[35].stu__mgr__cntl      =   stu__mgr35__cntl                ;
  assign   mgr__stu35__ready                =   mgr_inst[35].mgr__stu__ready    ;
  assign   mgr_inst[35].stu__mgr__type      =   stu__mgr35__type                ;
  assign   mgr_inst[35].stu__mgr__data      =   stu__mgr35__data                ;
  assign   mgr_inst[35].stu__mgr__oob_data  =   stu__mgr35__oob_data            ;

  assign   mgr_inst[36].stu__mgr__valid     =   stu__mgr36__valid               ;
  assign   mgr_inst[36].stu__mgr__cntl      =   stu__mgr36__cntl                ;
  assign   mgr__stu36__ready                =   mgr_inst[36].mgr__stu__ready    ;
  assign   mgr_inst[36].stu__mgr__type      =   stu__mgr36__type                ;
  assign   mgr_inst[36].stu__mgr__data      =   stu__mgr36__data                ;
  assign   mgr_inst[36].stu__mgr__oob_data  =   stu__mgr36__oob_data            ;

  assign   mgr_inst[37].stu__mgr__valid     =   stu__mgr37__valid               ;
  assign   mgr_inst[37].stu__mgr__cntl      =   stu__mgr37__cntl                ;
  assign   mgr__stu37__ready                =   mgr_inst[37].mgr__stu__ready    ;
  assign   mgr_inst[37].stu__mgr__type      =   stu__mgr37__type                ;
  assign   mgr_inst[37].stu__mgr__data      =   stu__mgr37__data                ;
  assign   mgr_inst[37].stu__mgr__oob_data  =   stu__mgr37__oob_data            ;

  assign   mgr_inst[38].stu__mgr__valid     =   stu__mgr38__valid               ;
  assign   mgr_inst[38].stu__mgr__cntl      =   stu__mgr38__cntl                ;
  assign   mgr__stu38__ready                =   mgr_inst[38].mgr__stu__ready    ;
  assign   mgr_inst[38].stu__mgr__type      =   stu__mgr38__type                ;
  assign   mgr_inst[38].stu__mgr__data      =   stu__mgr38__data                ;
  assign   mgr_inst[38].stu__mgr__oob_data  =   stu__mgr38__oob_data            ;

  assign   mgr_inst[39].stu__mgr__valid     =   stu__mgr39__valid               ;
  assign   mgr_inst[39].stu__mgr__cntl      =   stu__mgr39__cntl                ;
  assign   mgr__stu39__ready                =   mgr_inst[39].mgr__stu__ready    ;
  assign   mgr_inst[39].stu__mgr__type      =   stu__mgr39__type                ;
  assign   mgr_inst[39].stu__mgr__data      =   stu__mgr39__data                ;
  assign   mgr_inst[39].stu__mgr__oob_data  =   stu__mgr39__oob_data            ;

  assign   mgr_inst[40].stu__mgr__valid     =   stu__mgr40__valid               ;
  assign   mgr_inst[40].stu__mgr__cntl      =   stu__mgr40__cntl                ;
  assign   mgr__stu40__ready                =   mgr_inst[40].mgr__stu__ready    ;
  assign   mgr_inst[40].stu__mgr__type      =   stu__mgr40__type                ;
  assign   mgr_inst[40].stu__mgr__data      =   stu__mgr40__data                ;
  assign   mgr_inst[40].stu__mgr__oob_data  =   stu__mgr40__oob_data            ;

  assign   mgr_inst[41].stu__mgr__valid     =   stu__mgr41__valid               ;
  assign   mgr_inst[41].stu__mgr__cntl      =   stu__mgr41__cntl                ;
  assign   mgr__stu41__ready                =   mgr_inst[41].mgr__stu__ready    ;
  assign   mgr_inst[41].stu__mgr__type      =   stu__mgr41__type                ;
  assign   mgr_inst[41].stu__mgr__data      =   stu__mgr41__data                ;
  assign   mgr_inst[41].stu__mgr__oob_data  =   stu__mgr41__oob_data            ;

  assign   mgr_inst[42].stu__mgr__valid     =   stu__mgr42__valid               ;
  assign   mgr_inst[42].stu__mgr__cntl      =   stu__mgr42__cntl                ;
  assign   mgr__stu42__ready                =   mgr_inst[42].mgr__stu__ready    ;
  assign   mgr_inst[42].stu__mgr__type      =   stu__mgr42__type                ;
  assign   mgr_inst[42].stu__mgr__data      =   stu__mgr42__data                ;
  assign   mgr_inst[42].stu__mgr__oob_data  =   stu__mgr42__oob_data            ;

  assign   mgr_inst[43].stu__mgr__valid     =   stu__mgr43__valid               ;
  assign   mgr_inst[43].stu__mgr__cntl      =   stu__mgr43__cntl                ;
  assign   mgr__stu43__ready                =   mgr_inst[43].mgr__stu__ready    ;
  assign   mgr_inst[43].stu__mgr__type      =   stu__mgr43__type                ;
  assign   mgr_inst[43].stu__mgr__data      =   stu__mgr43__data                ;
  assign   mgr_inst[43].stu__mgr__oob_data  =   stu__mgr43__oob_data            ;

  assign   mgr_inst[44].stu__mgr__valid     =   stu__mgr44__valid               ;
  assign   mgr_inst[44].stu__mgr__cntl      =   stu__mgr44__cntl                ;
  assign   mgr__stu44__ready                =   mgr_inst[44].mgr__stu__ready    ;
  assign   mgr_inst[44].stu__mgr__type      =   stu__mgr44__type                ;
  assign   mgr_inst[44].stu__mgr__data      =   stu__mgr44__data                ;
  assign   mgr_inst[44].stu__mgr__oob_data  =   stu__mgr44__oob_data            ;

  assign   mgr_inst[45].stu__mgr__valid     =   stu__mgr45__valid               ;
  assign   mgr_inst[45].stu__mgr__cntl      =   stu__mgr45__cntl                ;
  assign   mgr__stu45__ready                =   mgr_inst[45].mgr__stu__ready    ;
  assign   mgr_inst[45].stu__mgr__type      =   stu__mgr45__type                ;
  assign   mgr_inst[45].stu__mgr__data      =   stu__mgr45__data                ;
  assign   mgr_inst[45].stu__mgr__oob_data  =   stu__mgr45__oob_data            ;

  assign   mgr_inst[46].stu__mgr__valid     =   stu__mgr46__valid               ;
  assign   mgr_inst[46].stu__mgr__cntl      =   stu__mgr46__cntl                ;
  assign   mgr__stu46__ready                =   mgr_inst[46].mgr__stu__ready    ;
  assign   mgr_inst[46].stu__mgr__type      =   stu__mgr46__type                ;
  assign   mgr_inst[46].stu__mgr__data      =   stu__mgr46__data                ;
  assign   mgr_inst[46].stu__mgr__oob_data  =   stu__mgr46__oob_data            ;

  assign   mgr_inst[47].stu__mgr__valid     =   stu__mgr47__valid               ;
  assign   mgr_inst[47].stu__mgr__cntl      =   stu__mgr47__cntl                ;
  assign   mgr__stu47__ready                =   mgr_inst[47].mgr__stu__ready    ;
  assign   mgr_inst[47].stu__mgr__type      =   stu__mgr47__type                ;
  assign   mgr_inst[47].stu__mgr__data      =   stu__mgr47__data                ;
  assign   mgr_inst[47].stu__mgr__oob_data  =   stu__mgr47__oob_data            ;

  assign   mgr_inst[48].stu__mgr__valid     =   stu__mgr48__valid               ;
  assign   mgr_inst[48].stu__mgr__cntl      =   stu__mgr48__cntl                ;
  assign   mgr__stu48__ready                =   mgr_inst[48].mgr__stu__ready    ;
  assign   mgr_inst[48].stu__mgr__type      =   stu__mgr48__type                ;
  assign   mgr_inst[48].stu__mgr__data      =   stu__mgr48__data                ;
  assign   mgr_inst[48].stu__mgr__oob_data  =   stu__mgr48__oob_data            ;

  assign   mgr_inst[49].stu__mgr__valid     =   stu__mgr49__valid               ;
  assign   mgr_inst[49].stu__mgr__cntl      =   stu__mgr49__cntl                ;
  assign   mgr__stu49__ready                =   mgr_inst[49].mgr__stu__ready    ;
  assign   mgr_inst[49].stu__mgr__type      =   stu__mgr49__type                ;
  assign   mgr_inst[49].stu__mgr__data      =   stu__mgr49__data                ;
  assign   mgr_inst[49].stu__mgr__oob_data  =   stu__mgr49__oob_data            ;

  assign   mgr_inst[50].stu__mgr__valid     =   stu__mgr50__valid               ;
  assign   mgr_inst[50].stu__mgr__cntl      =   stu__mgr50__cntl                ;
  assign   mgr__stu50__ready                =   mgr_inst[50].mgr__stu__ready    ;
  assign   mgr_inst[50].stu__mgr__type      =   stu__mgr50__type                ;
  assign   mgr_inst[50].stu__mgr__data      =   stu__mgr50__data                ;
  assign   mgr_inst[50].stu__mgr__oob_data  =   stu__mgr50__oob_data            ;

  assign   mgr_inst[51].stu__mgr__valid     =   stu__mgr51__valid               ;
  assign   mgr_inst[51].stu__mgr__cntl      =   stu__mgr51__cntl                ;
  assign   mgr__stu51__ready                =   mgr_inst[51].mgr__stu__ready    ;
  assign   mgr_inst[51].stu__mgr__type      =   stu__mgr51__type                ;
  assign   mgr_inst[51].stu__mgr__data      =   stu__mgr51__data                ;
  assign   mgr_inst[51].stu__mgr__oob_data  =   stu__mgr51__oob_data            ;

  assign   mgr_inst[52].stu__mgr__valid     =   stu__mgr52__valid               ;
  assign   mgr_inst[52].stu__mgr__cntl      =   stu__mgr52__cntl                ;
  assign   mgr__stu52__ready                =   mgr_inst[52].mgr__stu__ready    ;
  assign   mgr_inst[52].stu__mgr__type      =   stu__mgr52__type                ;
  assign   mgr_inst[52].stu__mgr__data      =   stu__mgr52__data                ;
  assign   mgr_inst[52].stu__mgr__oob_data  =   stu__mgr52__oob_data            ;

  assign   mgr_inst[53].stu__mgr__valid     =   stu__mgr53__valid               ;
  assign   mgr_inst[53].stu__mgr__cntl      =   stu__mgr53__cntl                ;
  assign   mgr__stu53__ready                =   mgr_inst[53].mgr__stu__ready    ;
  assign   mgr_inst[53].stu__mgr__type      =   stu__mgr53__type                ;
  assign   mgr_inst[53].stu__mgr__data      =   stu__mgr53__data                ;
  assign   mgr_inst[53].stu__mgr__oob_data  =   stu__mgr53__oob_data            ;

  assign   mgr_inst[54].stu__mgr__valid     =   stu__mgr54__valid               ;
  assign   mgr_inst[54].stu__mgr__cntl      =   stu__mgr54__cntl                ;
  assign   mgr__stu54__ready                =   mgr_inst[54].mgr__stu__ready    ;
  assign   mgr_inst[54].stu__mgr__type      =   stu__mgr54__type                ;
  assign   mgr_inst[54].stu__mgr__data      =   stu__mgr54__data                ;
  assign   mgr_inst[54].stu__mgr__oob_data  =   stu__mgr54__oob_data            ;

  assign   mgr_inst[55].stu__mgr__valid     =   stu__mgr55__valid               ;
  assign   mgr_inst[55].stu__mgr__cntl      =   stu__mgr55__cntl                ;
  assign   mgr__stu55__ready                =   mgr_inst[55].mgr__stu__ready    ;
  assign   mgr_inst[55].stu__mgr__type      =   stu__mgr55__type                ;
  assign   mgr_inst[55].stu__mgr__data      =   stu__mgr55__data                ;
  assign   mgr_inst[55].stu__mgr__oob_data  =   stu__mgr55__oob_data            ;

  assign   mgr_inst[56].stu__mgr__valid     =   stu__mgr56__valid               ;
  assign   mgr_inst[56].stu__mgr__cntl      =   stu__mgr56__cntl                ;
  assign   mgr__stu56__ready                =   mgr_inst[56].mgr__stu__ready    ;
  assign   mgr_inst[56].stu__mgr__type      =   stu__mgr56__type                ;
  assign   mgr_inst[56].stu__mgr__data      =   stu__mgr56__data                ;
  assign   mgr_inst[56].stu__mgr__oob_data  =   stu__mgr56__oob_data            ;

  assign   mgr_inst[57].stu__mgr__valid     =   stu__mgr57__valid               ;
  assign   mgr_inst[57].stu__mgr__cntl      =   stu__mgr57__cntl                ;
  assign   mgr__stu57__ready                =   mgr_inst[57].mgr__stu__ready    ;
  assign   mgr_inst[57].stu__mgr__type      =   stu__mgr57__type                ;
  assign   mgr_inst[57].stu__mgr__data      =   stu__mgr57__data                ;
  assign   mgr_inst[57].stu__mgr__oob_data  =   stu__mgr57__oob_data            ;

  assign   mgr_inst[58].stu__mgr__valid     =   stu__mgr58__valid               ;
  assign   mgr_inst[58].stu__mgr__cntl      =   stu__mgr58__cntl                ;
  assign   mgr__stu58__ready                =   mgr_inst[58].mgr__stu__ready    ;
  assign   mgr_inst[58].stu__mgr__type      =   stu__mgr58__type                ;
  assign   mgr_inst[58].stu__mgr__data      =   stu__mgr58__data                ;
  assign   mgr_inst[58].stu__mgr__oob_data  =   stu__mgr58__oob_data            ;

  assign   mgr_inst[59].stu__mgr__valid     =   stu__mgr59__valid               ;
  assign   mgr_inst[59].stu__mgr__cntl      =   stu__mgr59__cntl                ;
  assign   mgr__stu59__ready                =   mgr_inst[59].mgr__stu__ready    ;
  assign   mgr_inst[59].stu__mgr__type      =   stu__mgr59__type                ;
  assign   mgr_inst[59].stu__mgr__data      =   stu__mgr59__data                ;
  assign   mgr_inst[59].stu__mgr__oob_data  =   stu__mgr59__oob_data            ;

  assign   mgr_inst[60].stu__mgr__valid     =   stu__mgr60__valid               ;
  assign   mgr_inst[60].stu__mgr__cntl      =   stu__mgr60__cntl                ;
  assign   mgr__stu60__ready                =   mgr_inst[60].mgr__stu__ready    ;
  assign   mgr_inst[60].stu__mgr__type      =   stu__mgr60__type                ;
  assign   mgr_inst[60].stu__mgr__data      =   stu__mgr60__data                ;
  assign   mgr_inst[60].stu__mgr__oob_data  =   stu__mgr60__oob_data            ;

  assign   mgr_inst[61].stu__mgr__valid     =   stu__mgr61__valid               ;
  assign   mgr_inst[61].stu__mgr__cntl      =   stu__mgr61__cntl                ;
  assign   mgr__stu61__ready                =   mgr_inst[61].mgr__stu__ready    ;
  assign   mgr_inst[61].stu__mgr__type      =   stu__mgr61__type                ;
  assign   mgr_inst[61].stu__mgr__data      =   stu__mgr61__data                ;
  assign   mgr_inst[61].stu__mgr__oob_data  =   stu__mgr61__oob_data            ;

  assign   mgr_inst[62].stu__mgr__valid     =   stu__mgr62__valid               ;
  assign   mgr_inst[62].stu__mgr__cntl      =   stu__mgr62__cntl                ;
  assign   mgr__stu62__ready                =   mgr_inst[62].mgr__stu__ready    ;
  assign   mgr_inst[62].stu__mgr__type      =   stu__mgr62__type                ;
  assign   mgr_inst[62].stu__mgr__data      =   stu__mgr62__data                ;
  assign   mgr_inst[62].stu__mgr__oob_data  =   stu__mgr62__oob_data            ;

  assign   mgr_inst[63].stu__mgr__valid     =   stu__mgr63__valid               ;
  assign   mgr_inst[63].stu__mgr__cntl      =   stu__mgr63__cntl                ;
  assign   mgr__stu63__ready                =   mgr_inst[63].mgr__stu__ready    ;
  assign   mgr_inst[63].stu__mgr__type      =   stu__mgr63__type                ;
  assign   mgr_inst[63].stu__mgr__data      =   stu__mgr63__data                ;
  assign   mgr_inst[63].stu__mgr__oob_data  =   stu__mgr63__oob_data            ;

