
    wire                                           pe0__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe0__stu__cntl           ;
    wire                                           stu__pe0__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe0__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe0__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe0__stu__oob_data       ;

    wire                                           pe1__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe1__stu__cntl           ;
    wire                                           stu__pe1__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe1__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe1__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe1__stu__oob_data       ;

    wire                                           pe2__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe2__stu__cntl           ;
    wire                                           stu__pe2__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe2__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe2__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe2__stu__oob_data       ;

    wire                                           pe3__stu__valid          ;
    wire    [`COMMON_STD_INTF_CNTL_RANGE   ]       pe3__stu__cntl           ;
    wire                                           stu__pe3__ready          ;
    wire    [`STACK_UP_INTF_TYPE_RANGE     ]       pe3__stu__type           ;
    wire    [`STACK_UP_INTF_DATA_RANGE     ]       pe3__stu__data           ;
    wire    [`STACK_UP_INTF_OOB_DATA_RANGE ]       pe3__stu__oob_data       ;

