
            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            mgr0__std__oob_cntl                           ,
            mgr0__std__oob_valid                          ,
            std__mgr0__oob_ready                          ,
            mgr0__std__oob_type                           ,
            mgr0__std__oob_data                           ,

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            mgr1__std__oob_cntl                           ,
            mgr1__std__oob_valid                          ,
            std__mgr1__oob_ready                          ,
            mgr1__std__oob_type                           ,
            mgr1__std__oob_data                           ,

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            mgr2__std__oob_cntl                           ,
            mgr2__std__oob_valid                          ,
            std__mgr2__oob_ready                          ,
            mgr2__std__oob_type                           ,
            mgr2__std__oob_data                           ,

            // OOB controls the PE                          
            // For now assume OOB is separate to lanes      
            mgr3__std__oob_cntl                           ,
            mgr3__std__oob_valid                          ,
            std__mgr3__oob_ready                          ,
            mgr3__std__oob_type                           ,
            mgr3__std__oob_data                           ,
