
  // DMA port 0 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data0       ; 
  wire                                        memc__dma__read_data_valid0 ; 

  // DMA port 1 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data1       ; 
  wire                                        memc__dma__read_data_valid1 ; 

  // DMA port 2 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data2       ; 
  wire                                        memc__dma__read_data_valid2 ; 

  // DMA port 3 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data3       ; 
  wire                                        memc__dma__read_data_valid3 ; 

  // DMA port 4 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data4       ; 
  wire                                        memc__dma__read_data_valid4 ; 

  // DMA port 5 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data5       ; 
  wire                                        memc__dma__read_data_valid5 ; 

  // DMA port 6 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data6       ; 
  wire                                        memc__dma__read_data_valid6 ; 

  // DMA port 7 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data7       ; 
  wire                                        memc__dma__read_data_valid7 ; 

  // DMA port 8 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data8       ; 
  wire                                        memc__dma__read_data_valid8 ; 

  // DMA port 9 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data9       ; 
  wire                                        memc__dma__read_data_valid9 ; 

  // DMA port 10 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data10       ; 
  wire                                        memc__dma__read_data_valid10 ; 

  // DMA port 11 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data11       ; 
  wire                                        memc__dma__read_data_valid11 ; 

  // DMA port 12 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data12       ; 
  wire                                        memc__dma__read_data_valid12 ; 

  // DMA port 13 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data13       ; 
  wire                                        memc__dma__read_data_valid13 ; 

  // DMA port 14 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data14       ; 
  wire                                        memc__dma__read_data_valid14 ; 

  // DMA port 15 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data15       ; 
  wire                                        memc__dma__read_data_valid15 ; 

  // DMA port 16 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data16       ; 
  wire                                        memc__dma__read_data_valid16 ; 

  // DMA port 17 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data17       ; 
  wire                                        memc__dma__read_data_valid17 ; 

  // DMA port 18 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data18       ; 
  wire                                        memc__dma__read_data_valid18 ; 

  // DMA port 19 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data19       ; 
  wire                                        memc__dma__read_data_valid19 ; 

  // DMA port 20 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data20       ; 
  wire                                        memc__dma__read_data_valid20 ; 

  // DMA port 21 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data21       ; 
  wire                                        memc__dma__read_data_valid21 ; 

  // DMA port 22 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data22       ; 
  wire                                        memc__dma__read_data_valid22 ; 

  // DMA port 23 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data23       ; 
  wire                                        memc__dma__read_data_valid23 ; 

  // DMA port 24 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data24       ; 
  wire                                        memc__dma__read_data_valid24 ; 

  // DMA port 25 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data25       ; 
  wire                                        memc__dma__read_data_valid25 ; 

  // DMA port 26 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data26       ; 
  wire                                        memc__dma__read_data_valid26 ; 

  // DMA port 27 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data27       ; 
  wire                                        memc__dma__read_data_valid27 ; 

  // DMA port 28 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data28       ; 
  wire                                        memc__dma__read_data_valid28 ; 

  // DMA port 29 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data29       ; 
  wire                                        memc__dma__read_data_valid29 ; 

  // DMA port 30 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data30       ; 
  wire                                        memc__dma__read_data_valid30 ; 

  // DMA port 31 Read datapath signals
  wire [`MEM_ACC_CONT_MEMORY_DATA_RANGE    ]  memc__dma__read_data31       ; 
  wire                                        memc__dma__read_data_valid31 ; 


  // What bank is the LDST accessing
  // Bank0
  wire ldst_write_addr_to_bank0      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire ldst_read_addr_to_bank0       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd0)  ;
  wire ldst_write_request_to_bank0   =  ldst_write_addr_to_bank0    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank0    =  ldst_write_request_to_bank0 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank0    =  ldst_read_addr_to_bank0      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank0     =  ldst_read_request_to_bank0   & memc__ldst__read_ready   ;                                         
  // Bank1
  wire ldst_write_addr_to_bank1      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire ldst_read_addr_to_bank1       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd1)  ;
  wire ldst_write_request_to_bank1   =  ldst_write_addr_to_bank1    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank1    =  ldst_write_request_to_bank1 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank1    =  ldst_read_addr_to_bank1      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank1     =  ldst_read_request_to_bank1   & memc__ldst__read_ready   ;                                         
  // Bank2
  wire ldst_write_addr_to_bank2      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire ldst_read_addr_to_bank2       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd2)  ;
  wire ldst_write_request_to_bank2   =  ldst_write_addr_to_bank2    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank2    =  ldst_write_request_to_bank2 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank2    =  ldst_read_addr_to_bank2      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank2     =  ldst_read_request_to_bank2   & memc__ldst__read_ready   ;                                         
  // Bank3
  wire ldst_write_addr_to_bank3      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire ldst_read_addr_to_bank3       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd3)  ;
  wire ldst_write_request_to_bank3   =  ldst_write_addr_to_bank3    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank3    =  ldst_write_request_to_bank3 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank3    =  ldst_read_addr_to_bank3      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank3     =  ldst_read_request_to_bank3   & memc__ldst__read_ready   ;                                         
  // Bank4
  wire ldst_write_addr_to_bank4      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire ldst_read_addr_to_bank4       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd4)  ;
  wire ldst_write_request_to_bank4   =  ldst_write_addr_to_bank4    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank4    =  ldst_write_request_to_bank4 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank4    =  ldst_read_addr_to_bank4      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank4     =  ldst_read_request_to_bank4   & memc__ldst__read_ready   ;                                         
  // Bank5
  wire ldst_write_addr_to_bank5      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire ldst_read_addr_to_bank5       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd5)  ;
  wire ldst_write_request_to_bank5   =  ldst_write_addr_to_bank5    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank5    =  ldst_write_request_to_bank5 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank5    =  ldst_read_addr_to_bank5      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank5     =  ldst_read_request_to_bank5   & memc__ldst__read_ready   ;                                         
  // Bank6
  wire ldst_write_addr_to_bank6      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire ldst_read_addr_to_bank6       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd6)  ;
  wire ldst_write_request_to_bank6   =  ldst_write_addr_to_bank6    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank6    =  ldst_write_request_to_bank6 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank6    =  ldst_read_addr_to_bank6      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank6     =  ldst_read_request_to_bank6   & memc__ldst__read_ready   ;                                         
  // Bank7
  wire ldst_write_addr_to_bank7      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire ldst_read_addr_to_bank7       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd7)  ;
  wire ldst_write_request_to_bank7   =  ldst_write_addr_to_bank7    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank7    =  ldst_write_request_to_bank7 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank7    =  ldst_read_addr_to_bank7      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank7     =  ldst_read_request_to_bank7   & memc__ldst__read_ready   ;                                         
  // Bank8
  wire ldst_write_addr_to_bank8      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire ldst_read_addr_to_bank8       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd8)  ;
  wire ldst_write_request_to_bank8   =  ldst_write_addr_to_bank8    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank8    =  ldst_write_request_to_bank8 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank8    =  ldst_read_addr_to_bank8      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank8     =  ldst_read_request_to_bank8   & memc__ldst__read_ready   ;                                         
  // Bank9
  wire ldst_write_addr_to_bank9      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire ldst_read_addr_to_bank9       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd9)  ;
  wire ldst_write_request_to_bank9   =  ldst_write_addr_to_bank9    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank9    =  ldst_write_request_to_bank9 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank9    =  ldst_read_addr_to_bank9      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank9     =  ldst_read_request_to_bank9   & memc__ldst__read_ready   ;                                         
  // Bank10
  wire ldst_write_addr_to_bank10      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire ldst_read_addr_to_bank10       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd10)  ;
  wire ldst_write_request_to_bank10   =  ldst_write_addr_to_bank10    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank10    =  ldst_write_request_to_bank10 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank10    =  ldst_read_addr_to_bank10      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank10     =  ldst_read_request_to_bank10   & memc__ldst__read_ready   ;                                         
  // Bank11
  wire ldst_write_addr_to_bank11      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire ldst_read_addr_to_bank11       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd11)  ;
  wire ldst_write_request_to_bank11   =  ldst_write_addr_to_bank11    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank11    =  ldst_write_request_to_bank11 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank11    =  ldst_read_addr_to_bank11      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank11     =  ldst_read_request_to_bank11   & memc__ldst__read_ready   ;                                         
  // Bank12
  wire ldst_write_addr_to_bank12      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire ldst_read_addr_to_bank12       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd12)  ;
  wire ldst_write_request_to_bank12   =  ldst_write_addr_to_bank12    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank12    =  ldst_write_request_to_bank12 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank12    =  ldst_read_addr_to_bank12      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank12     =  ldst_read_request_to_bank12   & memc__ldst__read_ready   ;                                         
  // Bank13
  wire ldst_write_addr_to_bank13      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire ldst_read_addr_to_bank13       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd13)  ;
  wire ldst_write_request_to_bank13   =  ldst_write_addr_to_bank13    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank13    =  ldst_write_request_to_bank13 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank13    =  ldst_read_addr_to_bank13      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank13     =  ldst_read_request_to_bank13   & memc__ldst__read_ready   ;                                         
  // Bank14
  wire ldst_write_addr_to_bank14      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire ldst_read_addr_to_bank14       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd14)  ;
  wire ldst_write_request_to_bank14   =  ldst_write_addr_to_bank14    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank14    =  ldst_write_request_to_bank14 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank14    =  ldst_read_addr_to_bank14      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank14     =  ldst_read_request_to_bank14   & memc__ldst__read_ready   ;                                         
  // Bank15
  wire ldst_write_addr_to_bank15      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire ldst_read_addr_to_bank15       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd15)  ;
  wire ldst_write_request_to_bank15   =  ldst_write_addr_to_bank15    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank15    =  ldst_write_request_to_bank15 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank15    =  ldst_read_addr_to_bank15      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank15     =  ldst_read_request_to_bank15   & memc__ldst__read_ready   ;                                         
  // Bank16
  wire ldst_write_addr_to_bank16      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire ldst_read_addr_to_bank16       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd16)  ;
  wire ldst_write_request_to_bank16   =  ldst_write_addr_to_bank16    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank16    =  ldst_write_request_to_bank16 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank16    =  ldst_read_addr_to_bank16      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank16     =  ldst_read_request_to_bank16   & memc__ldst__read_ready   ;                                         
  // Bank17
  wire ldst_write_addr_to_bank17      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire ldst_read_addr_to_bank17       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd17)  ;
  wire ldst_write_request_to_bank17   =  ldst_write_addr_to_bank17    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank17    =  ldst_write_request_to_bank17 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank17    =  ldst_read_addr_to_bank17      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank17     =  ldst_read_request_to_bank17   & memc__ldst__read_ready   ;                                         
  // Bank18
  wire ldst_write_addr_to_bank18      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire ldst_read_addr_to_bank18       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd18)  ;
  wire ldst_write_request_to_bank18   =  ldst_write_addr_to_bank18    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank18    =  ldst_write_request_to_bank18 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank18    =  ldst_read_addr_to_bank18      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank18     =  ldst_read_request_to_bank18   & memc__ldst__read_ready   ;                                         
  // Bank19
  wire ldst_write_addr_to_bank19      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire ldst_read_addr_to_bank19       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd19)  ;
  wire ldst_write_request_to_bank19   =  ldst_write_addr_to_bank19    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank19    =  ldst_write_request_to_bank19 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank19    =  ldst_read_addr_to_bank19      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank19     =  ldst_read_request_to_bank19   & memc__ldst__read_ready   ;                                         
  // Bank20
  wire ldst_write_addr_to_bank20      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire ldst_read_addr_to_bank20       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd20)  ;
  wire ldst_write_request_to_bank20   =  ldst_write_addr_to_bank20    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank20    =  ldst_write_request_to_bank20 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank20    =  ldst_read_addr_to_bank20      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank20     =  ldst_read_request_to_bank20   & memc__ldst__read_ready   ;                                         
  // Bank21
  wire ldst_write_addr_to_bank21      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire ldst_read_addr_to_bank21       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd21)  ;
  wire ldst_write_request_to_bank21   =  ldst_write_addr_to_bank21    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank21    =  ldst_write_request_to_bank21 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank21    =  ldst_read_addr_to_bank21      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank21     =  ldst_read_request_to_bank21   & memc__ldst__read_ready   ;                                         
  // Bank22
  wire ldst_write_addr_to_bank22      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire ldst_read_addr_to_bank22       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd22)  ;
  wire ldst_write_request_to_bank22   =  ldst_write_addr_to_bank22    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank22    =  ldst_write_request_to_bank22 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank22    =  ldst_read_addr_to_bank22      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank22     =  ldst_read_request_to_bank22   & memc__ldst__read_ready   ;                                         
  // Bank23
  wire ldst_write_addr_to_bank23      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire ldst_read_addr_to_bank23       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd23)  ;
  wire ldst_write_request_to_bank23   =  ldst_write_addr_to_bank23    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank23    =  ldst_write_request_to_bank23 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank23    =  ldst_read_addr_to_bank23      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank23     =  ldst_read_request_to_bank23   & memc__ldst__read_ready   ;                                         
  // Bank24
  wire ldst_write_addr_to_bank24      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire ldst_read_addr_to_bank24       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd24)  ;
  wire ldst_write_request_to_bank24   =  ldst_write_addr_to_bank24    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank24    =  ldst_write_request_to_bank24 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank24    =  ldst_read_addr_to_bank24      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank24     =  ldst_read_request_to_bank24   & memc__ldst__read_ready   ;                                         
  // Bank25
  wire ldst_write_addr_to_bank25      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire ldst_read_addr_to_bank25       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd25)  ;
  wire ldst_write_request_to_bank25   =  ldst_write_addr_to_bank25    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank25    =  ldst_write_request_to_bank25 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank25    =  ldst_read_addr_to_bank25      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank25     =  ldst_read_request_to_bank25   & memc__ldst__read_ready   ;                                         
  // Bank26
  wire ldst_write_addr_to_bank26      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire ldst_read_addr_to_bank26       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd26)  ;
  wire ldst_write_request_to_bank26   =  ldst_write_addr_to_bank26    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank26    =  ldst_write_request_to_bank26 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank26    =  ldst_read_addr_to_bank26      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank26     =  ldst_read_request_to_bank26   & memc__ldst__read_ready   ;                                         
  // Bank27
  wire ldst_write_addr_to_bank27      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire ldst_read_addr_to_bank27       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd27)  ;
  wire ldst_write_request_to_bank27   =  ldst_write_addr_to_bank27    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank27    =  ldst_write_request_to_bank27 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank27    =  ldst_read_addr_to_bank27      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank27     =  ldst_read_request_to_bank27   & memc__ldst__read_ready   ;                                         
  // Bank28
  wire ldst_write_addr_to_bank28      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire ldst_read_addr_to_bank28       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd28)  ;
  wire ldst_write_request_to_bank28   =  ldst_write_addr_to_bank28    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank28    =  ldst_write_request_to_bank28 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank28    =  ldst_read_addr_to_bank28      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank28     =  ldst_read_request_to_bank28   & memc__ldst__read_ready   ;                                         
  // Bank29
  wire ldst_write_addr_to_bank29      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire ldst_read_addr_to_bank29       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd29)  ;
  wire ldst_write_request_to_bank29   =  ldst_write_addr_to_bank29    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank29    =  ldst_write_request_to_bank29 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank29    =  ldst_read_addr_to_bank29      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank29     =  ldst_read_request_to_bank29   & memc__ldst__read_ready   ;                                         
  // Bank30
  wire ldst_write_addr_to_bank30      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire ldst_read_addr_to_bank30       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd30)  ;
  wire ldst_write_request_to_bank30   =  ldst_write_addr_to_bank30    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank30    =  ldst_write_request_to_bank30 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank30    =  ldst_read_addr_to_bank30      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank30     =  ldst_read_request_to_bank30   & memc__ldst__read_ready   ;                                         
  // Bank31
  wire ldst_write_addr_to_bank31      =  (ldst__memc__write_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire ldst_read_addr_to_bank31       =  (ldst__memc__read_address[`MEM_ACC_CONT_MEMORY_ADDRESS_MSB  : `MEM_ACC_CONT_MEMORY_ADDRESS_MSB-4] == 5'd31)  ;
  wire ldst_write_request_to_bank31   =  ldst_write_addr_to_bank31    & ldst__memc__write_valid   ;                                         
  wire ldst_write_access_to_bank31    =  ldst_write_request_to_bank31 & memc__ldst__write_ready   ;  // request and ready to accept request 
  wire ldst_read_request_to_bank31    =  ldst_read_addr_to_bank31      & ldst__memc__read_valid   ;                                         
  wire ldst_read_access_to_bank31     =  ldst_read_request_to_bank31   & memc__ldst__read_ready   ;                                         

  // What banks are the DMA's accessing
  // DMA 0
  wire read_pause0     =  dma__memc__read_pause0   ;  
  // DMA/Bank 0
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request0_to_bank0   =  dma__memc__write_valid0  ;                                         
  wire write_access0_to_bank0    =  write_request0_to_bank0   & memc__dma__write_ready0  ;  // request and ready to accept request 
  wire read_request0_to_bank0    =  dma__memc__read_valid0   ;                                         
  wire read_access0_to_bank0     =  read_request0_to_bank0    & memc__dma__read_ready0   ;                                         
  // DMA 1
  wire read_pause1     =  dma__memc__read_pause1   ;  
  // DMA/Bank 1
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request1_to_bank1   =  dma__memc__write_valid1  ;                                         
  wire write_access1_to_bank1    =  write_request1_to_bank1   & memc__dma__write_ready1  ;  // request and ready to accept request 
  wire read_request1_to_bank1    =  dma__memc__read_valid1   ;                                         
  wire read_access1_to_bank1     =  read_request1_to_bank1    & memc__dma__read_ready1   ;                                         
  // DMA 2
  wire read_pause2     =  dma__memc__read_pause2   ;  
  // DMA/Bank 2
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request2_to_bank2   =  dma__memc__write_valid2  ;                                         
  wire write_access2_to_bank2    =  write_request2_to_bank2   & memc__dma__write_ready2  ;  // request and ready to accept request 
  wire read_request2_to_bank2    =  dma__memc__read_valid2   ;                                         
  wire read_access2_to_bank2     =  read_request2_to_bank2    & memc__dma__read_ready2   ;                                         
  // DMA 3
  wire read_pause3     =  dma__memc__read_pause3   ;  
  // DMA/Bank 3
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request3_to_bank3   =  dma__memc__write_valid3  ;                                         
  wire write_access3_to_bank3    =  write_request3_to_bank3   & memc__dma__write_ready3  ;  // request and ready to accept request 
  wire read_request3_to_bank3    =  dma__memc__read_valid3   ;                                         
  wire read_access3_to_bank3     =  read_request3_to_bank3    & memc__dma__read_ready3   ;                                         
  // DMA 4
  wire read_pause4     =  dma__memc__read_pause4   ;  
  // DMA/Bank 4
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request4_to_bank4   =  dma__memc__write_valid4  ;                                         
  wire write_access4_to_bank4    =  write_request4_to_bank4   & memc__dma__write_ready4  ;  // request and ready to accept request 
  wire read_request4_to_bank4    =  dma__memc__read_valid4   ;                                         
  wire read_access4_to_bank4     =  read_request4_to_bank4    & memc__dma__read_ready4   ;                                         
  // DMA 5
  wire read_pause5     =  dma__memc__read_pause5   ;  
  // DMA/Bank 5
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request5_to_bank5   =  dma__memc__write_valid5  ;                                         
  wire write_access5_to_bank5    =  write_request5_to_bank5   & memc__dma__write_ready5  ;  // request and ready to accept request 
  wire read_request5_to_bank5    =  dma__memc__read_valid5   ;                                         
  wire read_access5_to_bank5     =  read_request5_to_bank5    & memc__dma__read_ready5   ;                                         
  // DMA 6
  wire read_pause6     =  dma__memc__read_pause6   ;  
  // DMA/Bank 6
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request6_to_bank6   =  dma__memc__write_valid6  ;                                         
  wire write_access6_to_bank6    =  write_request6_to_bank6   & memc__dma__write_ready6  ;  // request and ready to accept request 
  wire read_request6_to_bank6    =  dma__memc__read_valid6   ;                                         
  wire read_access6_to_bank6     =  read_request6_to_bank6    & memc__dma__read_ready6   ;                                         
  // DMA 7
  wire read_pause7     =  dma__memc__read_pause7   ;  
  // DMA/Bank 7
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request7_to_bank7   =  dma__memc__write_valid7  ;                                         
  wire write_access7_to_bank7    =  write_request7_to_bank7   & memc__dma__write_ready7  ;  // request and ready to accept request 
  wire read_request7_to_bank7    =  dma__memc__read_valid7   ;                                         
  wire read_access7_to_bank7     =  read_request7_to_bank7    & memc__dma__read_ready7   ;                                         
  // DMA 8
  wire read_pause8     =  dma__memc__read_pause8   ;  
  // DMA/Bank 8
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request8_to_bank8   =  dma__memc__write_valid8  ;                                         
  wire write_access8_to_bank8    =  write_request8_to_bank8   & memc__dma__write_ready8  ;  // request and ready to accept request 
  wire read_request8_to_bank8    =  dma__memc__read_valid8   ;                                         
  wire read_access8_to_bank8     =  read_request8_to_bank8    & memc__dma__read_ready8   ;                                         
  // DMA 9
  wire read_pause9     =  dma__memc__read_pause9   ;  
  // DMA/Bank 9
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request9_to_bank9   =  dma__memc__write_valid9  ;                                         
  wire write_access9_to_bank9    =  write_request9_to_bank9   & memc__dma__write_ready9  ;  // request and ready to accept request 
  wire read_request9_to_bank9    =  dma__memc__read_valid9   ;                                         
  wire read_access9_to_bank9     =  read_request9_to_bank9    & memc__dma__read_ready9   ;                                         
  // DMA 10
  wire read_pause10     =  dma__memc__read_pause10   ;  
  // DMA/Bank 10
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request10_to_bank10   =  dma__memc__write_valid10  ;                                         
  wire write_access10_to_bank10    =  write_request10_to_bank10   & memc__dma__write_ready10  ;  // request and ready to accept request 
  wire read_request10_to_bank10    =  dma__memc__read_valid10   ;                                         
  wire read_access10_to_bank10     =  read_request10_to_bank10    & memc__dma__read_ready10   ;                                         
  // DMA 11
  wire read_pause11     =  dma__memc__read_pause11   ;  
  // DMA/Bank 11
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request11_to_bank11   =  dma__memc__write_valid11  ;                                         
  wire write_access11_to_bank11    =  write_request11_to_bank11   & memc__dma__write_ready11  ;  // request and ready to accept request 
  wire read_request11_to_bank11    =  dma__memc__read_valid11   ;                                         
  wire read_access11_to_bank11     =  read_request11_to_bank11    & memc__dma__read_ready11   ;                                         
  // DMA 12
  wire read_pause12     =  dma__memc__read_pause12   ;  
  // DMA/Bank 12
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request12_to_bank12   =  dma__memc__write_valid12  ;                                         
  wire write_access12_to_bank12    =  write_request12_to_bank12   & memc__dma__write_ready12  ;  // request and ready to accept request 
  wire read_request12_to_bank12    =  dma__memc__read_valid12   ;                                         
  wire read_access12_to_bank12     =  read_request12_to_bank12    & memc__dma__read_ready12   ;                                         
  // DMA 13
  wire read_pause13     =  dma__memc__read_pause13   ;  
  // DMA/Bank 13
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request13_to_bank13   =  dma__memc__write_valid13  ;                                         
  wire write_access13_to_bank13    =  write_request13_to_bank13   & memc__dma__write_ready13  ;  // request and ready to accept request 
  wire read_request13_to_bank13    =  dma__memc__read_valid13   ;                                         
  wire read_access13_to_bank13     =  read_request13_to_bank13    & memc__dma__read_ready13   ;                                         
  // DMA 14
  wire read_pause14     =  dma__memc__read_pause14   ;  
  // DMA/Bank 14
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request14_to_bank14   =  dma__memc__write_valid14  ;                                         
  wire write_access14_to_bank14    =  write_request14_to_bank14   & memc__dma__write_ready14  ;  // request and ready to accept request 
  wire read_request14_to_bank14    =  dma__memc__read_valid14   ;                                         
  wire read_access14_to_bank14     =  read_request14_to_bank14    & memc__dma__read_ready14   ;                                         
  // DMA 15
  wire read_pause15     =  dma__memc__read_pause15   ;  
  // DMA/Bank 15
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request15_to_bank15   =  dma__memc__write_valid15  ;                                         
  wire write_access15_to_bank15    =  write_request15_to_bank15   & memc__dma__write_ready15  ;  // request and ready to accept request 
  wire read_request15_to_bank15    =  dma__memc__read_valid15   ;                                         
  wire read_access15_to_bank15     =  read_request15_to_bank15    & memc__dma__read_ready15   ;                                         
  // DMA 16
  wire read_pause16     =  dma__memc__read_pause16   ;  
  // DMA/Bank 16
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request16_to_bank16   =  dma__memc__write_valid16  ;                                         
  wire write_access16_to_bank16    =  write_request16_to_bank16   & memc__dma__write_ready16  ;  // request and ready to accept request 
  wire read_request16_to_bank16    =  dma__memc__read_valid16   ;                                         
  wire read_access16_to_bank16     =  read_request16_to_bank16    & memc__dma__read_ready16   ;                                         
  // DMA 17
  wire read_pause17     =  dma__memc__read_pause17   ;  
  // DMA/Bank 17
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request17_to_bank17   =  dma__memc__write_valid17  ;                                         
  wire write_access17_to_bank17    =  write_request17_to_bank17   & memc__dma__write_ready17  ;  // request and ready to accept request 
  wire read_request17_to_bank17    =  dma__memc__read_valid17   ;                                         
  wire read_access17_to_bank17     =  read_request17_to_bank17    & memc__dma__read_ready17   ;                                         
  // DMA 18
  wire read_pause18     =  dma__memc__read_pause18   ;  
  // DMA/Bank 18
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request18_to_bank18   =  dma__memc__write_valid18  ;                                         
  wire write_access18_to_bank18    =  write_request18_to_bank18   & memc__dma__write_ready18  ;  // request and ready to accept request 
  wire read_request18_to_bank18    =  dma__memc__read_valid18   ;                                         
  wire read_access18_to_bank18     =  read_request18_to_bank18    & memc__dma__read_ready18   ;                                         
  // DMA 19
  wire read_pause19     =  dma__memc__read_pause19   ;  
  // DMA/Bank 19
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request19_to_bank19   =  dma__memc__write_valid19  ;                                         
  wire write_access19_to_bank19    =  write_request19_to_bank19   & memc__dma__write_ready19  ;  // request and ready to accept request 
  wire read_request19_to_bank19    =  dma__memc__read_valid19   ;                                         
  wire read_access19_to_bank19     =  read_request19_to_bank19    & memc__dma__read_ready19   ;                                         
  // DMA 20
  wire read_pause20     =  dma__memc__read_pause20   ;  
  // DMA/Bank 20
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request20_to_bank20   =  dma__memc__write_valid20  ;                                         
  wire write_access20_to_bank20    =  write_request20_to_bank20   & memc__dma__write_ready20  ;  // request and ready to accept request 
  wire read_request20_to_bank20    =  dma__memc__read_valid20   ;                                         
  wire read_access20_to_bank20     =  read_request20_to_bank20    & memc__dma__read_ready20   ;                                         
  // DMA 21
  wire read_pause21     =  dma__memc__read_pause21   ;  
  // DMA/Bank 21
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request21_to_bank21   =  dma__memc__write_valid21  ;                                         
  wire write_access21_to_bank21    =  write_request21_to_bank21   & memc__dma__write_ready21  ;  // request and ready to accept request 
  wire read_request21_to_bank21    =  dma__memc__read_valid21   ;                                         
  wire read_access21_to_bank21     =  read_request21_to_bank21    & memc__dma__read_ready21   ;                                         
  // DMA 22
  wire read_pause22     =  dma__memc__read_pause22   ;  
  // DMA/Bank 22
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request22_to_bank22   =  dma__memc__write_valid22  ;                                         
  wire write_access22_to_bank22    =  write_request22_to_bank22   & memc__dma__write_ready22  ;  // request and ready to accept request 
  wire read_request22_to_bank22    =  dma__memc__read_valid22   ;                                         
  wire read_access22_to_bank22     =  read_request22_to_bank22    & memc__dma__read_ready22   ;                                         
  // DMA 23
  wire read_pause23     =  dma__memc__read_pause23   ;  
  // DMA/Bank 23
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request23_to_bank23   =  dma__memc__write_valid23  ;                                         
  wire write_access23_to_bank23    =  write_request23_to_bank23   & memc__dma__write_ready23  ;  // request and ready to accept request 
  wire read_request23_to_bank23    =  dma__memc__read_valid23   ;                                         
  wire read_access23_to_bank23     =  read_request23_to_bank23    & memc__dma__read_ready23   ;                                         
  // DMA 24
  wire read_pause24     =  dma__memc__read_pause24   ;  
  // DMA/Bank 24
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request24_to_bank24   =  dma__memc__write_valid24  ;                                         
  wire write_access24_to_bank24    =  write_request24_to_bank24   & memc__dma__write_ready24  ;  // request and ready to accept request 
  wire read_request24_to_bank24    =  dma__memc__read_valid24   ;                                         
  wire read_access24_to_bank24     =  read_request24_to_bank24    & memc__dma__read_ready24   ;                                         
  // DMA 25
  wire read_pause25     =  dma__memc__read_pause25   ;  
  // DMA/Bank 25
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request25_to_bank25   =  dma__memc__write_valid25  ;                                         
  wire write_access25_to_bank25    =  write_request25_to_bank25   & memc__dma__write_ready25  ;  // request and ready to accept request 
  wire read_request25_to_bank25    =  dma__memc__read_valid25   ;                                         
  wire read_access25_to_bank25     =  read_request25_to_bank25    & memc__dma__read_ready25   ;                                         
  // DMA 26
  wire read_pause26     =  dma__memc__read_pause26   ;  
  // DMA/Bank 26
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request26_to_bank26   =  dma__memc__write_valid26  ;                                         
  wire write_access26_to_bank26    =  write_request26_to_bank26   & memc__dma__write_ready26  ;  // request and ready to accept request 
  wire read_request26_to_bank26    =  dma__memc__read_valid26   ;                                         
  wire read_access26_to_bank26     =  read_request26_to_bank26    & memc__dma__read_ready26   ;                                         
  // DMA 27
  wire read_pause27     =  dma__memc__read_pause27   ;  
  // DMA/Bank 27
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request27_to_bank27   =  dma__memc__write_valid27  ;                                         
  wire write_access27_to_bank27    =  write_request27_to_bank27   & memc__dma__write_ready27  ;  // request and ready to accept request 
  wire read_request27_to_bank27    =  dma__memc__read_valid27   ;                                         
  wire read_access27_to_bank27     =  read_request27_to_bank27    & memc__dma__read_ready27   ;                                         
  // DMA 28
  wire read_pause28     =  dma__memc__read_pause28   ;  
  // DMA/Bank 28
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request28_to_bank28   =  dma__memc__write_valid28  ;                                         
  wire write_access28_to_bank28    =  write_request28_to_bank28   & memc__dma__write_ready28  ;  // request and ready to accept request 
  wire read_request28_to_bank28    =  dma__memc__read_valid28   ;                                         
  wire read_access28_to_bank28     =  read_request28_to_bank28    & memc__dma__read_ready28   ;                                         
  // DMA 29
  wire read_pause29     =  dma__memc__read_pause29   ;  
  // DMA/Bank 29
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request29_to_bank29   =  dma__memc__write_valid29  ;                                         
  wire write_access29_to_bank29    =  write_request29_to_bank29   & memc__dma__write_ready29  ;  // request and ready to accept request 
  wire read_request29_to_bank29    =  dma__memc__read_valid29   ;                                         
  wire read_access29_to_bank29     =  read_request29_to_bank29    & memc__dma__read_ready29   ;                                         
  // DMA 30
  wire read_pause30     =  dma__memc__read_pause30   ;  
  // DMA/Bank 30
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request30_to_bank30   =  dma__memc__write_valid30  ;                                         
  wire write_access30_to_bank30    =  write_request30_to_bank30   & memc__dma__write_ready30  ;  // request and ready to accept request 
  wire read_request30_to_bank30    =  dma__memc__read_valid30   ;                                         
  wire read_access30_to_bank30     =  read_request30_to_bank30    & memc__dma__read_ready30   ;                                         
  // DMA 31
  wire read_pause31     =  dma__memc__read_pause31   ;  
  // DMA/Bank 31
  // Signals indicating whether a request is being made and if the request is accepted
  wire write_request31_to_bank31   =  dma__memc__write_valid31  ;                                         
  wire write_access31_to_bank31    =  write_request31_to_bank31   & memc__dma__write_ready31  ;  // request and ready to accept request 
  wire read_request31_to_bank31    =  dma__memc__read_valid31   ;                                         
  wire read_access31_to_bank31     =  read_request31_to_bank31    & memc__dma__read_ready31   ;                                         