
  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe0__allSynchronized    ( GenStackBus[0].sys__pe__allSynchronized           ), 
        .pe0__sys__thisSynchronized   ( GenStackBus[0].pe__sys__thisSynchronized          ), 
        .pe0__sys__ready              ( GenStackBus[0].pe__sys__ready                     ), 
        .pe0__sys__complete           ( GenStackBus[0].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe1__allSynchronized    ( GenStackBus[1].sys__pe__allSynchronized           ), 
        .pe1__sys__thisSynchronized   ( GenStackBus[1].pe__sys__thisSynchronized          ), 
        .pe1__sys__ready              ( GenStackBus[1].pe__sys__ready                     ), 
        .pe1__sys__complete           ( GenStackBus[1].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe2__allSynchronized    ( GenStackBus[2].sys__pe__allSynchronized           ), 
        .pe2__sys__thisSynchronized   ( GenStackBus[2].pe__sys__thisSynchronized          ), 
        .pe2__sys__ready              ( GenStackBus[2].pe__sys__ready                     ), 
        .pe2__sys__complete           ( GenStackBus[2].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe3__allSynchronized    ( GenStackBus[3].sys__pe__allSynchronized           ), 
        .pe3__sys__thisSynchronized   ( GenStackBus[3].pe__sys__thisSynchronized          ), 
        .pe3__sys__ready              ( GenStackBus[3].pe__sys__ready                     ), 
        .pe3__sys__complete           ( GenStackBus[3].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe4__allSynchronized    ( GenStackBus[4].sys__pe__allSynchronized           ), 
        .pe4__sys__thisSynchronized   ( GenStackBus[4].pe__sys__thisSynchronized          ), 
        .pe4__sys__ready              ( GenStackBus[4].pe__sys__ready                     ), 
        .pe4__sys__complete           ( GenStackBus[4].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe5__allSynchronized    ( GenStackBus[5].sys__pe__allSynchronized           ), 
        .pe5__sys__thisSynchronized   ( GenStackBus[5].pe__sys__thisSynchronized          ), 
        .pe5__sys__ready              ( GenStackBus[5].pe__sys__ready                     ), 
        .pe5__sys__complete           ( GenStackBus[5].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe6__allSynchronized    ( GenStackBus[6].sys__pe__allSynchronized           ), 
        .pe6__sys__thisSynchronized   ( GenStackBus[6].pe__sys__thisSynchronized          ), 
        .pe6__sys__ready              ( GenStackBus[6].pe__sys__ready                     ), 
        .pe6__sys__complete           ( GenStackBus[6].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe7__allSynchronized    ( GenStackBus[7].sys__pe__allSynchronized           ), 
        .pe7__sys__thisSynchronized   ( GenStackBus[7].pe__sys__thisSynchronized          ), 
        .pe7__sys__ready              ( GenStackBus[7].pe__sys__ready                     ), 
        .pe7__sys__complete           ( GenStackBus[7].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe8__allSynchronized    ( GenStackBus[8].sys__pe__allSynchronized           ), 
        .pe8__sys__thisSynchronized   ( GenStackBus[8].pe__sys__thisSynchronized          ), 
        .pe8__sys__ready              ( GenStackBus[8].pe__sys__ready                     ), 
        .pe8__sys__complete           ( GenStackBus[8].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe9__allSynchronized    ( GenStackBus[9].sys__pe__allSynchronized           ), 
        .pe9__sys__thisSynchronized   ( GenStackBus[9].pe__sys__thisSynchronized          ), 
        .pe9__sys__ready              ( GenStackBus[9].pe__sys__ready                     ), 
        .pe9__sys__complete           ( GenStackBus[9].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe10__allSynchronized    ( GenStackBus[10].sys__pe__allSynchronized           ), 
        .pe10__sys__thisSynchronized   ( GenStackBus[10].pe__sys__thisSynchronized          ), 
        .pe10__sys__ready              ( GenStackBus[10].pe__sys__ready                     ), 
        .pe10__sys__complete           ( GenStackBus[10].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe11__allSynchronized    ( GenStackBus[11].sys__pe__allSynchronized           ), 
        .pe11__sys__thisSynchronized   ( GenStackBus[11].pe__sys__thisSynchronized          ), 
        .pe11__sys__ready              ( GenStackBus[11].pe__sys__ready                     ), 
        .pe11__sys__complete           ( GenStackBus[11].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe12__allSynchronized    ( GenStackBus[12].sys__pe__allSynchronized           ), 
        .pe12__sys__thisSynchronized   ( GenStackBus[12].pe__sys__thisSynchronized          ), 
        .pe12__sys__ready              ( GenStackBus[12].pe__sys__ready                     ), 
        .pe12__sys__complete           ( GenStackBus[12].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe13__allSynchronized    ( GenStackBus[13].sys__pe__allSynchronized           ), 
        .pe13__sys__thisSynchronized   ( GenStackBus[13].pe__sys__thisSynchronized          ), 
        .pe13__sys__ready              ( GenStackBus[13].pe__sys__ready                     ), 
        .pe13__sys__complete           ( GenStackBus[13].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe14__allSynchronized    ( GenStackBus[14].sys__pe__allSynchronized           ), 
        .pe14__sys__thisSynchronized   ( GenStackBus[14].pe__sys__thisSynchronized          ), 
        .pe14__sys__ready              ( GenStackBus[14].pe__sys__ready                     ), 
        .pe14__sys__complete           ( GenStackBus[14].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe15__allSynchronized    ( GenStackBus[15].sys__pe__allSynchronized           ), 
        .pe15__sys__thisSynchronized   ( GenStackBus[15].pe__sys__thisSynchronized          ), 
        .pe15__sys__ready              ( GenStackBus[15].pe__sys__ready                     ), 
        .pe15__sys__complete           ( GenStackBus[15].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe16__allSynchronized    ( GenStackBus[16].sys__pe__allSynchronized           ), 
        .pe16__sys__thisSynchronized   ( GenStackBus[16].pe__sys__thisSynchronized          ), 
        .pe16__sys__ready              ( GenStackBus[16].pe__sys__ready                     ), 
        .pe16__sys__complete           ( GenStackBus[16].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe17__allSynchronized    ( GenStackBus[17].sys__pe__allSynchronized           ), 
        .pe17__sys__thisSynchronized   ( GenStackBus[17].pe__sys__thisSynchronized          ), 
        .pe17__sys__ready              ( GenStackBus[17].pe__sys__ready                     ), 
        .pe17__sys__complete           ( GenStackBus[17].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe18__allSynchronized    ( GenStackBus[18].sys__pe__allSynchronized           ), 
        .pe18__sys__thisSynchronized   ( GenStackBus[18].pe__sys__thisSynchronized          ), 
        .pe18__sys__ready              ( GenStackBus[18].pe__sys__ready                     ), 
        .pe18__sys__complete           ( GenStackBus[18].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe19__allSynchronized    ( GenStackBus[19].sys__pe__allSynchronized           ), 
        .pe19__sys__thisSynchronized   ( GenStackBus[19].pe__sys__thisSynchronized          ), 
        .pe19__sys__ready              ( GenStackBus[19].pe__sys__ready                     ), 
        .pe19__sys__complete           ( GenStackBus[19].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe20__allSynchronized    ( GenStackBus[20].sys__pe__allSynchronized           ), 
        .pe20__sys__thisSynchronized   ( GenStackBus[20].pe__sys__thisSynchronized          ), 
        .pe20__sys__ready              ( GenStackBus[20].pe__sys__ready                     ), 
        .pe20__sys__complete           ( GenStackBus[20].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe21__allSynchronized    ( GenStackBus[21].sys__pe__allSynchronized           ), 
        .pe21__sys__thisSynchronized   ( GenStackBus[21].pe__sys__thisSynchronized          ), 
        .pe21__sys__ready              ( GenStackBus[21].pe__sys__ready                     ), 
        .pe21__sys__complete           ( GenStackBus[21].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe22__allSynchronized    ( GenStackBus[22].sys__pe__allSynchronized           ), 
        .pe22__sys__thisSynchronized   ( GenStackBus[22].pe__sys__thisSynchronized          ), 
        .pe22__sys__ready              ( GenStackBus[22].pe__sys__ready                     ), 
        .pe22__sys__complete           ( GenStackBus[22].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe23__allSynchronized    ( GenStackBus[23].sys__pe__allSynchronized           ), 
        .pe23__sys__thisSynchronized   ( GenStackBus[23].pe__sys__thisSynchronized          ), 
        .pe23__sys__ready              ( GenStackBus[23].pe__sys__ready                     ), 
        .pe23__sys__complete           ( GenStackBus[23].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe24__allSynchronized    ( GenStackBus[24].sys__pe__allSynchronized           ), 
        .pe24__sys__thisSynchronized   ( GenStackBus[24].pe__sys__thisSynchronized          ), 
        .pe24__sys__ready              ( GenStackBus[24].pe__sys__ready                     ), 
        .pe24__sys__complete           ( GenStackBus[24].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe25__allSynchronized    ( GenStackBus[25].sys__pe__allSynchronized           ), 
        .pe25__sys__thisSynchronized   ( GenStackBus[25].pe__sys__thisSynchronized          ), 
        .pe25__sys__ready              ( GenStackBus[25].pe__sys__ready                     ), 
        .pe25__sys__complete           ( GenStackBus[25].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe26__allSynchronized    ( GenStackBus[26].sys__pe__allSynchronized           ), 
        .pe26__sys__thisSynchronized   ( GenStackBus[26].pe__sys__thisSynchronized          ), 
        .pe26__sys__ready              ( GenStackBus[26].pe__sys__ready                     ), 
        .pe26__sys__complete           ( GenStackBus[26].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe27__allSynchronized    ( GenStackBus[27].sys__pe__allSynchronized           ), 
        .pe27__sys__thisSynchronized   ( GenStackBus[27].pe__sys__thisSynchronized          ), 
        .pe27__sys__ready              ( GenStackBus[27].pe__sys__ready                     ), 
        .pe27__sys__complete           ( GenStackBus[27].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe28__allSynchronized    ( GenStackBus[28].sys__pe__allSynchronized           ), 
        .pe28__sys__thisSynchronized   ( GenStackBus[28].pe__sys__thisSynchronized          ), 
        .pe28__sys__ready              ( GenStackBus[28].pe__sys__ready                     ), 
        .pe28__sys__complete           ( GenStackBus[28].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe29__allSynchronized    ( GenStackBus[29].sys__pe__allSynchronized           ), 
        .pe29__sys__thisSynchronized   ( GenStackBus[29].pe__sys__thisSynchronized          ), 
        .pe29__sys__ready              ( GenStackBus[29].pe__sys__ready                     ), 
        .pe29__sys__complete           ( GenStackBus[29].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe30__allSynchronized    ( GenStackBus[30].sys__pe__allSynchronized           ), 
        .pe30__sys__thisSynchronized   ( GenStackBus[30].pe__sys__thisSynchronized          ), 
        .pe30__sys__ready              ( GenStackBus[30].pe__sys__ready                     ), 
        .pe30__sys__complete           ( GenStackBus[30].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe31__allSynchronized    ( GenStackBus[31].sys__pe__allSynchronized           ), 
        .pe31__sys__thisSynchronized   ( GenStackBus[31].pe__sys__thisSynchronized          ), 
        .pe31__sys__ready              ( GenStackBus[31].pe__sys__ready                     ), 
        .pe31__sys__complete           ( GenStackBus[31].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe32__allSynchronized    ( GenStackBus[32].sys__pe__allSynchronized           ), 
        .pe32__sys__thisSynchronized   ( GenStackBus[32].pe__sys__thisSynchronized          ), 
        .pe32__sys__ready              ( GenStackBus[32].pe__sys__ready                     ), 
        .pe32__sys__complete           ( GenStackBus[32].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe33__allSynchronized    ( GenStackBus[33].sys__pe__allSynchronized           ), 
        .pe33__sys__thisSynchronized   ( GenStackBus[33].pe__sys__thisSynchronized          ), 
        .pe33__sys__ready              ( GenStackBus[33].pe__sys__ready                     ), 
        .pe33__sys__complete           ( GenStackBus[33].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe34__allSynchronized    ( GenStackBus[34].sys__pe__allSynchronized           ), 
        .pe34__sys__thisSynchronized   ( GenStackBus[34].pe__sys__thisSynchronized          ), 
        .pe34__sys__ready              ( GenStackBus[34].pe__sys__ready                     ), 
        .pe34__sys__complete           ( GenStackBus[34].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe35__allSynchronized    ( GenStackBus[35].sys__pe__allSynchronized           ), 
        .pe35__sys__thisSynchronized   ( GenStackBus[35].pe__sys__thisSynchronized          ), 
        .pe35__sys__ready              ( GenStackBus[35].pe__sys__ready                     ), 
        .pe35__sys__complete           ( GenStackBus[35].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe36__allSynchronized    ( GenStackBus[36].sys__pe__allSynchronized           ), 
        .pe36__sys__thisSynchronized   ( GenStackBus[36].pe__sys__thisSynchronized          ), 
        .pe36__sys__ready              ( GenStackBus[36].pe__sys__ready                     ), 
        .pe36__sys__complete           ( GenStackBus[36].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe37__allSynchronized    ( GenStackBus[37].sys__pe__allSynchronized           ), 
        .pe37__sys__thisSynchronized   ( GenStackBus[37].pe__sys__thisSynchronized          ), 
        .pe37__sys__ready              ( GenStackBus[37].pe__sys__ready                     ), 
        .pe37__sys__complete           ( GenStackBus[37].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe38__allSynchronized    ( GenStackBus[38].sys__pe__allSynchronized           ), 
        .pe38__sys__thisSynchronized   ( GenStackBus[38].pe__sys__thisSynchronized          ), 
        .pe38__sys__ready              ( GenStackBus[38].pe__sys__ready                     ), 
        .pe38__sys__complete           ( GenStackBus[38].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe39__allSynchronized    ( GenStackBus[39].sys__pe__allSynchronized           ), 
        .pe39__sys__thisSynchronized   ( GenStackBus[39].pe__sys__thisSynchronized          ), 
        .pe39__sys__ready              ( GenStackBus[39].pe__sys__ready                     ), 
        .pe39__sys__complete           ( GenStackBus[39].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe40__allSynchronized    ( GenStackBus[40].sys__pe__allSynchronized           ), 
        .pe40__sys__thisSynchronized   ( GenStackBus[40].pe__sys__thisSynchronized          ), 
        .pe40__sys__ready              ( GenStackBus[40].pe__sys__ready                     ), 
        .pe40__sys__complete           ( GenStackBus[40].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe41__allSynchronized    ( GenStackBus[41].sys__pe__allSynchronized           ), 
        .pe41__sys__thisSynchronized   ( GenStackBus[41].pe__sys__thisSynchronized          ), 
        .pe41__sys__ready              ( GenStackBus[41].pe__sys__ready                     ), 
        .pe41__sys__complete           ( GenStackBus[41].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe42__allSynchronized    ( GenStackBus[42].sys__pe__allSynchronized           ), 
        .pe42__sys__thisSynchronized   ( GenStackBus[42].pe__sys__thisSynchronized          ), 
        .pe42__sys__ready              ( GenStackBus[42].pe__sys__ready                     ), 
        .pe42__sys__complete           ( GenStackBus[42].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe43__allSynchronized    ( GenStackBus[43].sys__pe__allSynchronized           ), 
        .pe43__sys__thisSynchronized   ( GenStackBus[43].pe__sys__thisSynchronized          ), 
        .pe43__sys__ready              ( GenStackBus[43].pe__sys__ready                     ), 
        .pe43__sys__complete           ( GenStackBus[43].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe44__allSynchronized    ( GenStackBus[44].sys__pe__allSynchronized           ), 
        .pe44__sys__thisSynchronized   ( GenStackBus[44].pe__sys__thisSynchronized          ), 
        .pe44__sys__ready              ( GenStackBus[44].pe__sys__ready                     ), 
        .pe44__sys__complete           ( GenStackBus[44].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe45__allSynchronized    ( GenStackBus[45].sys__pe__allSynchronized           ), 
        .pe45__sys__thisSynchronized   ( GenStackBus[45].pe__sys__thisSynchronized          ), 
        .pe45__sys__ready              ( GenStackBus[45].pe__sys__ready                     ), 
        .pe45__sys__complete           ( GenStackBus[45].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe46__allSynchronized    ( GenStackBus[46].sys__pe__allSynchronized           ), 
        .pe46__sys__thisSynchronized   ( GenStackBus[46].pe__sys__thisSynchronized          ), 
        .pe46__sys__ready              ( GenStackBus[46].pe__sys__ready                     ), 
        .pe46__sys__complete           ( GenStackBus[46].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe47__allSynchronized    ( GenStackBus[47].sys__pe__allSynchronized           ), 
        .pe47__sys__thisSynchronized   ( GenStackBus[47].pe__sys__thisSynchronized          ), 
        .pe47__sys__ready              ( GenStackBus[47].pe__sys__ready                     ), 
        .pe47__sys__complete           ( GenStackBus[47].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe48__allSynchronized    ( GenStackBus[48].sys__pe__allSynchronized           ), 
        .pe48__sys__thisSynchronized   ( GenStackBus[48].pe__sys__thisSynchronized          ), 
        .pe48__sys__ready              ( GenStackBus[48].pe__sys__ready                     ), 
        .pe48__sys__complete           ( GenStackBus[48].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe49__allSynchronized    ( GenStackBus[49].sys__pe__allSynchronized           ), 
        .pe49__sys__thisSynchronized   ( GenStackBus[49].pe__sys__thisSynchronized          ), 
        .pe49__sys__ready              ( GenStackBus[49].pe__sys__ready                     ), 
        .pe49__sys__complete           ( GenStackBus[49].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe50__allSynchronized    ( GenStackBus[50].sys__pe__allSynchronized           ), 
        .pe50__sys__thisSynchronized   ( GenStackBus[50].pe__sys__thisSynchronized          ), 
        .pe50__sys__ready              ( GenStackBus[50].pe__sys__ready                     ), 
        .pe50__sys__complete           ( GenStackBus[50].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe51__allSynchronized    ( GenStackBus[51].sys__pe__allSynchronized           ), 
        .pe51__sys__thisSynchronized   ( GenStackBus[51].pe__sys__thisSynchronized          ), 
        .pe51__sys__ready              ( GenStackBus[51].pe__sys__ready                     ), 
        .pe51__sys__complete           ( GenStackBus[51].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe52__allSynchronized    ( GenStackBus[52].sys__pe__allSynchronized           ), 
        .pe52__sys__thisSynchronized   ( GenStackBus[52].pe__sys__thisSynchronized          ), 
        .pe52__sys__ready              ( GenStackBus[52].pe__sys__ready                     ), 
        .pe52__sys__complete           ( GenStackBus[52].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe53__allSynchronized    ( GenStackBus[53].sys__pe__allSynchronized           ), 
        .pe53__sys__thisSynchronized   ( GenStackBus[53].pe__sys__thisSynchronized          ), 
        .pe53__sys__ready              ( GenStackBus[53].pe__sys__ready                     ), 
        .pe53__sys__complete           ( GenStackBus[53].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe54__allSynchronized    ( GenStackBus[54].sys__pe__allSynchronized           ), 
        .pe54__sys__thisSynchronized   ( GenStackBus[54].pe__sys__thisSynchronized          ), 
        .pe54__sys__ready              ( GenStackBus[54].pe__sys__ready                     ), 
        .pe54__sys__complete           ( GenStackBus[54].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe55__allSynchronized    ( GenStackBus[55].sys__pe__allSynchronized           ), 
        .pe55__sys__thisSynchronized   ( GenStackBus[55].pe__sys__thisSynchronized          ), 
        .pe55__sys__ready              ( GenStackBus[55].pe__sys__ready                     ), 
        .pe55__sys__complete           ( GenStackBus[55].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe56__allSynchronized    ( GenStackBus[56].sys__pe__allSynchronized           ), 
        .pe56__sys__thisSynchronized   ( GenStackBus[56].pe__sys__thisSynchronized          ), 
        .pe56__sys__ready              ( GenStackBus[56].pe__sys__ready                     ), 
        .pe56__sys__complete           ( GenStackBus[56].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe57__allSynchronized    ( GenStackBus[57].sys__pe__allSynchronized           ), 
        .pe57__sys__thisSynchronized   ( GenStackBus[57].pe__sys__thisSynchronized          ), 
        .pe57__sys__ready              ( GenStackBus[57].pe__sys__ready                     ), 
        .pe57__sys__complete           ( GenStackBus[57].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe58__allSynchronized    ( GenStackBus[58].sys__pe__allSynchronized           ), 
        .pe58__sys__thisSynchronized   ( GenStackBus[58].pe__sys__thisSynchronized          ), 
        .pe58__sys__ready              ( GenStackBus[58].pe__sys__ready                     ), 
        .pe58__sys__complete           ( GenStackBus[58].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe59__allSynchronized    ( GenStackBus[59].sys__pe__allSynchronized           ), 
        .pe59__sys__thisSynchronized   ( GenStackBus[59].pe__sys__thisSynchronized          ), 
        .pe59__sys__ready              ( GenStackBus[59].pe__sys__ready                     ), 
        .pe59__sys__complete           ( GenStackBus[59].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe60__allSynchronized    ( GenStackBus[60].sys__pe__allSynchronized           ), 
        .pe60__sys__thisSynchronized   ( GenStackBus[60].pe__sys__thisSynchronized          ), 
        .pe60__sys__ready              ( GenStackBus[60].pe__sys__ready                     ), 
        .pe60__sys__complete           ( GenStackBus[60].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe61__allSynchronized    ( GenStackBus[61].sys__pe__allSynchronized           ), 
        .pe61__sys__thisSynchronized   ( GenStackBus[61].pe__sys__thisSynchronized          ), 
        .pe61__sys__ready              ( GenStackBus[61].pe__sys__ready                     ), 
        .pe61__sys__complete           ( GenStackBus[61].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe62__allSynchronized    ( GenStackBus[62].sys__pe__allSynchronized           ), 
        .pe62__sys__thisSynchronized   ( GenStackBus[62].pe__sys__thisSynchronized          ), 
        .pe62__sys__ready              ( GenStackBus[62].pe__sys__ready                     ), 
        .pe62__sys__complete           ( GenStackBus[62].pe__sys__complete                  ), 

  // General control and status                                                                     
  //  - doesnt seem to work if you use cb_test for observed signals                                 
  //  - tried all combinations, e.g. cb_test to grab the signal and no cb for checking etc.         
        .sys__pe63__allSynchronized    ( GenStackBus[63].sys__pe__allSynchronized           ), 
        .pe63__sys__thisSynchronized   ( GenStackBus[63].pe__sys__thisSynchronized          ), 
        .pe63__sys__ready              ( GenStackBus[63].pe__sys__ready                     ), 
        .pe63__sys__complete           ( GenStackBus[63].pe__sys__complete                  ), 
