
    input                                         stu__mgr0__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr0__cntl           ;
    output                                        mgr0__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr0__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr0__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr0__oob_data       ;

    input                                         stu__mgr1__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr1__cntl           ;
    output                                        mgr1__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr1__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr1__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr1__oob_data       ;

    input                                         stu__mgr2__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr2__cntl           ;
    output                                        mgr2__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr2__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr2__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr2__oob_data       ;

    input                                         stu__mgr3__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr3__cntl           ;
    output                                        mgr3__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr3__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr3__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr3__oob_data       ;

    input                                         stu__mgr4__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr4__cntl           ;
    output                                        mgr4__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr4__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr4__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr4__oob_data       ;

    input                                         stu__mgr5__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr5__cntl           ;
    output                                        mgr5__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr5__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr5__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr5__oob_data       ;

    input                                         stu__mgr6__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr6__cntl           ;
    output                                        mgr6__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr6__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr6__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr6__oob_data       ;

    input                                         stu__mgr7__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr7__cntl           ;
    output                                        mgr7__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr7__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr7__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr7__oob_data       ;

    input                                         stu__mgr8__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr8__cntl           ;
    output                                        mgr8__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr8__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr8__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr8__oob_data       ;

    input                                         stu__mgr9__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr9__cntl           ;
    output                                        mgr9__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr9__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr9__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr9__oob_data       ;

    input                                         stu__mgr10__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr10__cntl           ;
    output                                        mgr10__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr10__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr10__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr10__oob_data       ;

    input                                         stu__mgr11__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr11__cntl           ;
    output                                        mgr11__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr11__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr11__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr11__oob_data       ;

    input                                         stu__mgr12__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr12__cntl           ;
    output                                        mgr12__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr12__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr12__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr12__oob_data       ;

    input                                         stu__mgr13__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr13__cntl           ;
    output                                        mgr13__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr13__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr13__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr13__oob_data       ;

    input                                         stu__mgr14__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr14__cntl           ;
    output                                        mgr14__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr14__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr14__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr14__oob_data       ;

    input                                         stu__mgr15__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr15__cntl           ;
    output                                        mgr15__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr15__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr15__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr15__oob_data       ;

    input                                         stu__mgr16__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr16__cntl           ;
    output                                        mgr16__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr16__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr16__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr16__oob_data       ;

    input                                         stu__mgr17__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr17__cntl           ;
    output                                        mgr17__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr17__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr17__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr17__oob_data       ;

    input                                         stu__mgr18__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr18__cntl           ;
    output                                        mgr18__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr18__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr18__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr18__oob_data       ;

    input                                         stu__mgr19__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr19__cntl           ;
    output                                        mgr19__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr19__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr19__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr19__oob_data       ;

    input                                         stu__mgr20__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr20__cntl           ;
    output                                        mgr20__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr20__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr20__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr20__oob_data       ;

    input                                         stu__mgr21__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr21__cntl           ;
    output                                        mgr21__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr21__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr21__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr21__oob_data       ;

    input                                         stu__mgr22__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr22__cntl           ;
    output                                        mgr22__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr22__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr22__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr22__oob_data       ;

    input                                         stu__mgr23__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr23__cntl           ;
    output                                        mgr23__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr23__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr23__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr23__oob_data       ;

    input                                         stu__mgr24__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr24__cntl           ;
    output                                        mgr24__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr24__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr24__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr24__oob_data       ;

    input                                         stu__mgr25__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr25__cntl           ;
    output                                        mgr25__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr25__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr25__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr25__oob_data       ;

    input                                         stu__mgr26__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr26__cntl           ;
    output                                        mgr26__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr26__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr26__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr26__oob_data       ;

    input                                         stu__mgr27__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr27__cntl           ;
    output                                        mgr27__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr27__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr27__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr27__oob_data       ;

    input                                         stu__mgr28__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr28__cntl           ;
    output                                        mgr28__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr28__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr28__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr28__oob_data       ;

    input                                         stu__mgr29__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr29__cntl           ;
    output                                        mgr29__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr29__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr29__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr29__oob_data       ;

    input                                         stu__mgr30__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr30__cntl           ;
    output                                        mgr30__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr30__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr30__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr30__oob_data       ;

    input                                         stu__mgr31__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr31__cntl           ;
    output                                        mgr31__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr31__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr31__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr31__oob_data       ;

    input                                         stu__mgr32__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr32__cntl           ;
    output                                        mgr32__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr32__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr32__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr32__oob_data       ;

    input                                         stu__mgr33__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr33__cntl           ;
    output                                        mgr33__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr33__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr33__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr33__oob_data       ;

    input                                         stu__mgr34__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr34__cntl           ;
    output                                        mgr34__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr34__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr34__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr34__oob_data       ;

    input                                         stu__mgr35__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr35__cntl           ;
    output                                        mgr35__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr35__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr35__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr35__oob_data       ;

    input                                         stu__mgr36__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr36__cntl           ;
    output                                        mgr36__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr36__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr36__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr36__oob_data       ;

    input                                         stu__mgr37__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr37__cntl           ;
    output                                        mgr37__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr37__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr37__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr37__oob_data       ;

    input                                         stu__mgr38__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr38__cntl           ;
    output                                        mgr38__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr38__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr38__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr38__oob_data       ;

    input                                         stu__mgr39__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr39__cntl           ;
    output                                        mgr39__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr39__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr39__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr39__oob_data       ;

    input                                         stu__mgr40__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr40__cntl           ;
    output                                        mgr40__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr40__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr40__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr40__oob_data       ;

    input                                         stu__mgr41__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr41__cntl           ;
    output                                        mgr41__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr41__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr41__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr41__oob_data       ;

    input                                         stu__mgr42__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr42__cntl           ;
    output                                        mgr42__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr42__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr42__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr42__oob_data       ;

    input                                         stu__mgr43__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr43__cntl           ;
    output                                        mgr43__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr43__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr43__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr43__oob_data       ;

    input                                         stu__mgr44__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr44__cntl           ;
    output                                        mgr44__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr44__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr44__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr44__oob_data       ;

    input                                         stu__mgr45__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr45__cntl           ;
    output                                        mgr45__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr45__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr45__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr45__oob_data       ;

    input                                         stu__mgr46__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr46__cntl           ;
    output                                        mgr46__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr46__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr46__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr46__oob_data       ;

    input                                         stu__mgr47__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr47__cntl           ;
    output                                        mgr47__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr47__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr47__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr47__oob_data       ;

    input                                         stu__mgr48__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr48__cntl           ;
    output                                        mgr48__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr48__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr48__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr48__oob_data       ;

    input                                         stu__mgr49__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr49__cntl           ;
    output                                        mgr49__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr49__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr49__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr49__oob_data       ;

    input                                         stu__mgr50__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr50__cntl           ;
    output                                        mgr50__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr50__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr50__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr50__oob_data       ;

    input                                         stu__mgr51__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr51__cntl           ;
    output                                        mgr51__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr51__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr51__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr51__oob_data       ;

    input                                         stu__mgr52__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr52__cntl           ;
    output                                        mgr52__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr52__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr52__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr52__oob_data       ;

    input                                         stu__mgr53__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr53__cntl           ;
    output                                        mgr53__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr53__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr53__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr53__oob_data       ;

    input                                         stu__mgr54__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr54__cntl           ;
    output                                        mgr54__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr54__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr54__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr54__oob_data       ;

    input                                         stu__mgr55__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr55__cntl           ;
    output                                        mgr55__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr55__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr55__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr55__oob_data       ;

    input                                         stu__mgr56__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr56__cntl           ;
    output                                        mgr56__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr56__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr56__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr56__oob_data       ;

    input                                         stu__mgr57__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr57__cntl           ;
    output                                        mgr57__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr57__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr57__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr57__oob_data       ;

    input                                         stu__mgr58__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr58__cntl           ;
    output                                        mgr58__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr58__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr58__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr58__oob_data       ;

    input                                         stu__mgr59__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr59__cntl           ;
    output                                        mgr59__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr59__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr59__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr59__oob_data       ;

    input                                         stu__mgr60__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr60__cntl           ;
    output                                        mgr60__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr60__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr60__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr60__oob_data       ;

    input                                         stu__mgr61__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr61__cntl           ;
    output                                        mgr61__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr61__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr61__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr61__oob_data       ;

    input                                         stu__mgr62__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr62__cntl           ;
    output                                        mgr62__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr62__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr62__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr62__oob_data       ;

    input                                         stu__mgr63__valid          ;
    input  [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr63__cntl           ;
    output                                        mgr63__stu__ready          ;
    input  [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr63__type           ;
    input  [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr63__data           ;
    input  [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr63__oob_data       ;

