
        wire                                      read_data_strm0_valid_next  ;  
        reg                                       read_data_strm0_valid       ;  
        wire                                      dma_read_addr0_to_bank        ;  
        wire                                      dma_write_addr0_to_bank       ;  
        wire                                      read_data_strm1_valid_next  ;  
        reg                                       read_data_strm1_valid       ;  
        wire                                      dma_read_addr1_to_bank        ;  
        wire                                      dma_write_addr1_to_bank       ;  
        wire                                      read_data_strm2_valid_next  ;  
        reg                                       read_data_strm2_valid       ;  
        wire                                      dma_read_addr2_to_bank        ;  
        wire                                      dma_write_addr2_to_bank       ;  
        wire                                      read_data_strm3_valid_next  ;  
        reg                                       read_data_strm3_valid       ;  
        wire                                      dma_read_addr3_to_bank        ;  
        wire                                      dma_write_addr3_to_bank       ;  
        wire                                      read_data_strm4_valid_next  ;  
        reg                                       read_data_strm4_valid       ;  
        wire                                      dma_read_addr4_to_bank        ;  
        wire                                      dma_write_addr4_to_bank       ;  
        wire                                      read_data_strm5_valid_next  ;  
        reg                                       read_data_strm5_valid       ;  
        wire                                      dma_read_addr5_to_bank        ;  
        wire                                      dma_write_addr5_to_bank       ;  
        wire                                      read_data_strm6_valid_next  ;  
        reg                                       read_data_strm6_valid       ;  
        wire                                      dma_read_addr6_to_bank        ;  
        wire                                      dma_write_addr6_to_bank       ;  
        wire                                      read_data_strm7_valid_next  ;  
        reg                                       read_data_strm7_valid       ;  
        wire                                      dma_read_addr7_to_bank        ;  
        wire                                      dma_write_addr7_to_bank       ;  
        wire                                      read_data_strm8_valid_next  ;  
        reg                                       read_data_strm8_valid       ;  
        wire                                      dma_read_addr8_to_bank        ;  
        wire                                      dma_write_addr8_to_bank       ;  
        wire                                      read_data_strm9_valid_next  ;  
        reg                                       read_data_strm9_valid       ;  
        wire                                      dma_read_addr9_to_bank        ;  
        wire                                      dma_write_addr9_to_bank       ;  
        wire                                      read_data_strm10_valid_next  ;  
        reg                                       read_data_strm10_valid       ;  
        wire                                      dma_read_addr10_to_bank        ;  
        wire                                      dma_write_addr10_to_bank       ;  
        wire                                      read_data_strm11_valid_next  ;  
        reg                                       read_data_strm11_valid       ;  
        wire                                      dma_read_addr11_to_bank        ;  
        wire                                      dma_write_addr11_to_bank       ;  
        wire                                      read_data_strm12_valid_next  ;  
        reg                                       read_data_strm12_valid       ;  
        wire                                      dma_read_addr12_to_bank        ;  
        wire                                      dma_write_addr12_to_bank       ;  
        wire                                      read_data_strm13_valid_next  ;  
        reg                                       read_data_strm13_valid       ;  
        wire                                      dma_read_addr13_to_bank        ;  
        wire                                      dma_write_addr13_to_bank       ;  
        wire                                      read_data_strm14_valid_next  ;  
        reg                                       read_data_strm14_valid       ;  
        wire                                      dma_read_addr14_to_bank        ;  
        wire                                      dma_write_addr14_to_bank       ;  
        wire                                      read_data_strm15_valid_next  ;  
        reg                                       read_data_strm15_valid       ;  
        wire                                      dma_read_addr15_to_bank        ;  
        wire                                      dma_write_addr15_to_bank       ;  
        wire                                      read_data_strm16_valid_next  ;  
        reg                                       read_data_strm16_valid       ;  
        wire                                      dma_read_addr16_to_bank        ;  
        wire                                      dma_write_addr16_to_bank       ;  
        wire                                      read_data_strm17_valid_next  ;  
        reg                                       read_data_strm17_valid       ;  
        wire                                      dma_read_addr17_to_bank        ;  
        wire                                      dma_write_addr17_to_bank       ;  
        wire                                      read_data_strm18_valid_next  ;  
        reg                                       read_data_strm18_valid       ;  
        wire                                      dma_read_addr18_to_bank        ;  
        wire                                      dma_write_addr18_to_bank       ;  
        wire                                      read_data_strm19_valid_next  ;  
        reg                                       read_data_strm19_valid       ;  
        wire                                      dma_read_addr19_to_bank        ;  
        wire                                      dma_write_addr19_to_bank       ;  
        wire                                      read_data_strm20_valid_next  ;  
        reg                                       read_data_strm20_valid       ;  
        wire                                      dma_read_addr20_to_bank        ;  
        wire                                      dma_write_addr20_to_bank       ;  
        wire                                      read_data_strm21_valid_next  ;  
        reg                                       read_data_strm21_valid       ;  
        wire                                      dma_read_addr21_to_bank        ;  
        wire                                      dma_write_addr21_to_bank       ;  
        wire                                      read_data_strm22_valid_next  ;  
        reg                                       read_data_strm22_valid       ;  
        wire                                      dma_read_addr22_to_bank        ;  
        wire                                      dma_write_addr22_to_bank       ;  
        wire                                      read_data_strm23_valid_next  ;  
        reg                                       read_data_strm23_valid       ;  
        wire                                      dma_read_addr23_to_bank        ;  
        wire                                      dma_write_addr23_to_bank       ;  
        wire                                      read_data_strm24_valid_next  ;  
        reg                                       read_data_strm24_valid       ;  
        wire                                      dma_read_addr24_to_bank        ;  
        wire                                      dma_write_addr24_to_bank       ;  
        wire                                      read_data_strm25_valid_next  ;  
        reg                                       read_data_strm25_valid       ;  
        wire                                      dma_read_addr25_to_bank        ;  
        wire                                      dma_write_addr25_to_bank       ;  
        wire                                      read_data_strm26_valid_next  ;  
        reg                                       read_data_strm26_valid       ;  
        wire                                      dma_read_addr26_to_bank        ;  
        wire                                      dma_write_addr26_to_bank       ;  
        wire                                      read_data_strm27_valid_next  ;  
        reg                                       read_data_strm27_valid       ;  
        wire                                      dma_read_addr27_to_bank        ;  
        wire                                      dma_write_addr27_to_bank       ;  
        wire                                      read_data_strm28_valid_next  ;  
        reg                                       read_data_strm28_valid       ;  
        wire                                      dma_read_addr28_to_bank        ;  
        wire                                      dma_write_addr28_to_bank       ;  
        wire                                      read_data_strm29_valid_next  ;  
        reg                                       read_data_strm29_valid       ;  
        wire                                      dma_read_addr29_to_bank        ;  
        wire                                      dma_write_addr29_to_bank       ;  
        wire                                      read_data_strm30_valid_next  ;  
        reg                                       read_data_strm30_valid       ;  
        wire                                      dma_read_addr30_to_bank        ;  
        wire                                      dma_write_addr30_to_bank       ;  
        wire                                      read_data_strm31_valid_next  ;  
        reg                                       read_data_strm31_valid       ;  
        wire                                      dma_read_addr31_to_bank        ;  
        wire                                      dma_write_addr31_to_bank       ;  