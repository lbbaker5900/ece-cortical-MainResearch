`ifndef _TB_common_vh_
`define _TB_common_vh_

//----------------------------------------------------------------------------------------------------
// Define what drives SIMD registers into streamingOps_cntl
//
//`define TB_ENABLE_REGFILE_DRIVER
//`undef  TB_ENABLE_REGFILE_DRIVER

`endif
