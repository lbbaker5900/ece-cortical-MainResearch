`ifndef _wu_memory_vh
`define _wu_memory_vh

/*****************************************************************

    File name   : wu_memory.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : Mar 2017
    email       : lbbaker@ncsu.edu

*****************************************************************/


//--------------------------------------------------------
  
//------------------------------------------------------------------------------------------------------------


`endif
