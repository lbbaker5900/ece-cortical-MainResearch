
    input                                          stu__mgr0__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr0__cntl           ;
    output                                         mgr0__stu__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr0__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr0__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr0__oob_data       ;

    input                                          stu__mgr1__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr1__cntl           ;
    output                                         mgr1__stu__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr1__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr1__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr1__oob_data       ;

    input                                          stu__mgr2__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr2__cntl           ;
    output                                         mgr2__stu__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr2__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr2__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr2__oob_data       ;

    input                                          stu__mgr3__valid          ;
    input   [`COMMON_STD_INTF_CNTL_RANGE   ]       stu__mgr3__cntl           ;
    output                                         mgr3__stu__ready          ;
    input   [`STACK_UP_INTF_TYPE_RANGE     ]       stu__mgr3__type           ;
    input   [`STACK_UP_INTF_DATA_RANGE     ]       stu__mgr3__data           ;
    input   [`STACK_UP_INTF_OOB_DATA_RANGE ]       stu__mgr3__oob_data       ;

