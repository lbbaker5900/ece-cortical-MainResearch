
                // Memory Port 0                 
                .dma__memc__write_valid0       ( dma__memc__lane0_write_valid0     ),
                .dma__memc__write_address0     ( dma__memc__lane0_write_address0   ),
                .dma__memc__write_data0        ( dma__memc__lane0_write_data0      ),
                .memc__dma__write_ready0       ( memc__dma__lane0_write_ready0     ),
                .dma__memc__read_valid0        ( dma__memc__lane0_read_valid0      ),
                .dma__memc__read_address0      ( dma__memc__lane0_read_address0    ),
                .memc__dma__read_data0         ( memc__dma__lane0_read_data0       ),
                .memc__dma__read_data_valid0   ( memc__dma__lane0_read_data_valid0 ),
                .memc__dma__read_ready0        ( memc__dma__lane0_read_ready0      ),
                .dma__memc__read_pause0        ( dma__memc__lane0_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid1       ( dma__memc__lane1_write_valid0     ),
                .dma__memc__write_address1     ( dma__memc__lane1_write_address0   ),
                .dma__memc__write_data1        ( dma__memc__lane1_write_data0      ),
                .memc__dma__write_ready1       ( memc__dma__lane1_write_ready0     ),
                .dma__memc__read_valid1        ( dma__memc__lane1_read_valid0      ),
                .dma__memc__read_address1      ( dma__memc__lane1_read_address0    ),
                .memc__dma__read_data1         ( memc__dma__lane1_read_data0       ),
                .memc__dma__read_data_valid1   ( memc__dma__lane1_read_data_valid0 ),
                .memc__dma__read_ready1        ( memc__dma__lane1_read_ready0      ),
                .dma__memc__read_pause1        ( dma__memc__lane1_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid2       ( dma__memc__lane2_write_valid0     ),
                .dma__memc__write_address2     ( dma__memc__lane2_write_address0   ),
                .dma__memc__write_data2        ( dma__memc__lane2_write_data0      ),
                .memc__dma__write_ready2       ( memc__dma__lane2_write_ready0     ),
                .dma__memc__read_valid2        ( dma__memc__lane2_read_valid0      ),
                .dma__memc__read_address2      ( dma__memc__lane2_read_address0    ),
                .memc__dma__read_data2         ( memc__dma__lane2_read_data0       ),
                .memc__dma__read_data_valid2   ( memc__dma__lane2_read_data_valid0 ),
                .memc__dma__read_ready2        ( memc__dma__lane2_read_ready0      ),
                .dma__memc__read_pause2        ( dma__memc__lane2_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid3       ( dma__memc__lane3_write_valid0     ),
                .dma__memc__write_address3     ( dma__memc__lane3_write_address0   ),
                .dma__memc__write_data3        ( dma__memc__lane3_write_data0      ),
                .memc__dma__write_ready3       ( memc__dma__lane3_write_ready0     ),
                .dma__memc__read_valid3        ( dma__memc__lane3_read_valid0      ),
                .dma__memc__read_address3      ( dma__memc__lane3_read_address0    ),
                .memc__dma__read_data3         ( memc__dma__lane3_read_data0       ),
                .memc__dma__read_data_valid3   ( memc__dma__lane3_read_data_valid0 ),
                .memc__dma__read_ready3        ( memc__dma__lane3_read_ready0      ),
                .dma__memc__read_pause3        ( dma__memc__lane3_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid4       ( dma__memc__lane4_write_valid0     ),
                .dma__memc__write_address4     ( dma__memc__lane4_write_address0   ),
                .dma__memc__write_data4        ( dma__memc__lane4_write_data0      ),
                .memc__dma__write_ready4       ( memc__dma__lane4_write_ready0     ),
                .dma__memc__read_valid4        ( dma__memc__lane4_read_valid0      ),
                .dma__memc__read_address4      ( dma__memc__lane4_read_address0    ),
                .memc__dma__read_data4         ( memc__dma__lane4_read_data0       ),
                .memc__dma__read_data_valid4   ( memc__dma__lane4_read_data_valid0 ),
                .memc__dma__read_ready4        ( memc__dma__lane4_read_ready0      ),
                .dma__memc__read_pause4        ( dma__memc__lane4_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid5       ( dma__memc__lane5_write_valid0     ),
                .dma__memc__write_address5     ( dma__memc__lane5_write_address0   ),
                .dma__memc__write_data5        ( dma__memc__lane5_write_data0      ),
                .memc__dma__write_ready5       ( memc__dma__lane5_write_ready0     ),
                .dma__memc__read_valid5        ( dma__memc__lane5_read_valid0      ),
                .dma__memc__read_address5      ( dma__memc__lane5_read_address0    ),
                .memc__dma__read_data5         ( memc__dma__lane5_read_data0       ),
                .memc__dma__read_data_valid5   ( memc__dma__lane5_read_data_valid0 ),
                .memc__dma__read_ready5        ( memc__dma__lane5_read_ready0      ),
                .dma__memc__read_pause5        ( dma__memc__lane5_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid6       ( dma__memc__lane6_write_valid0     ),
                .dma__memc__write_address6     ( dma__memc__lane6_write_address0   ),
                .dma__memc__write_data6        ( dma__memc__lane6_write_data0      ),
                .memc__dma__write_ready6       ( memc__dma__lane6_write_ready0     ),
                .dma__memc__read_valid6        ( dma__memc__lane6_read_valid0      ),
                .dma__memc__read_address6      ( dma__memc__lane6_read_address0    ),
                .memc__dma__read_data6         ( memc__dma__lane6_read_data0       ),
                .memc__dma__read_data_valid6   ( memc__dma__lane6_read_data_valid0 ),
                .memc__dma__read_ready6        ( memc__dma__lane6_read_ready0      ),
                .dma__memc__read_pause6        ( dma__memc__lane6_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid7       ( dma__memc__lane7_write_valid0     ),
                .dma__memc__write_address7     ( dma__memc__lane7_write_address0   ),
                .dma__memc__write_data7        ( dma__memc__lane7_write_data0      ),
                .memc__dma__write_ready7       ( memc__dma__lane7_write_ready0     ),
                .dma__memc__read_valid7        ( dma__memc__lane7_read_valid0      ),
                .dma__memc__read_address7      ( dma__memc__lane7_read_address0    ),
                .memc__dma__read_data7         ( memc__dma__lane7_read_data0       ),
                .memc__dma__read_data_valid7   ( memc__dma__lane7_read_data_valid0 ),
                .memc__dma__read_ready7        ( memc__dma__lane7_read_ready0      ),
                .dma__memc__read_pause7        ( dma__memc__lane7_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid8       ( dma__memc__lane8_write_valid0     ),
                .dma__memc__write_address8     ( dma__memc__lane8_write_address0   ),
                .dma__memc__write_data8        ( dma__memc__lane8_write_data0      ),
                .memc__dma__write_ready8       ( memc__dma__lane8_write_ready0     ),
                .dma__memc__read_valid8        ( dma__memc__lane8_read_valid0      ),
                .dma__memc__read_address8      ( dma__memc__lane8_read_address0    ),
                .memc__dma__read_data8         ( memc__dma__lane8_read_data0       ),
                .memc__dma__read_data_valid8   ( memc__dma__lane8_read_data_valid0 ),
                .memc__dma__read_ready8        ( memc__dma__lane8_read_ready0      ),
                .dma__memc__read_pause8        ( dma__memc__lane8_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid9       ( dma__memc__lane9_write_valid0     ),
                .dma__memc__write_address9     ( dma__memc__lane9_write_address0   ),
                .dma__memc__write_data9        ( dma__memc__lane9_write_data0      ),
                .memc__dma__write_ready9       ( memc__dma__lane9_write_ready0     ),
                .dma__memc__read_valid9        ( dma__memc__lane9_read_valid0      ),
                .dma__memc__read_address9      ( dma__memc__lane9_read_address0    ),
                .memc__dma__read_data9         ( memc__dma__lane9_read_data0       ),
                .memc__dma__read_data_valid9   ( memc__dma__lane9_read_data_valid0 ),
                .memc__dma__read_ready9        ( memc__dma__lane9_read_ready0      ),
                .dma__memc__read_pause9        ( dma__memc__lane9_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid10       ( dma__memc__lane10_write_valid0     ),
                .dma__memc__write_address10     ( dma__memc__lane10_write_address0   ),
                .dma__memc__write_data10        ( dma__memc__lane10_write_data0      ),
                .memc__dma__write_ready10       ( memc__dma__lane10_write_ready0     ),
                .dma__memc__read_valid10        ( dma__memc__lane10_read_valid0      ),
                .dma__memc__read_address10      ( dma__memc__lane10_read_address0    ),
                .memc__dma__read_data10         ( memc__dma__lane10_read_data0       ),
                .memc__dma__read_data_valid10   ( memc__dma__lane10_read_data_valid0 ),
                .memc__dma__read_ready10        ( memc__dma__lane10_read_ready0      ),
                .dma__memc__read_pause10        ( dma__memc__lane10_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid11       ( dma__memc__lane11_write_valid0     ),
                .dma__memc__write_address11     ( dma__memc__lane11_write_address0   ),
                .dma__memc__write_data11        ( dma__memc__lane11_write_data0      ),
                .memc__dma__write_ready11       ( memc__dma__lane11_write_ready0     ),
                .dma__memc__read_valid11        ( dma__memc__lane11_read_valid0      ),
                .dma__memc__read_address11      ( dma__memc__lane11_read_address0    ),
                .memc__dma__read_data11         ( memc__dma__lane11_read_data0       ),
                .memc__dma__read_data_valid11   ( memc__dma__lane11_read_data_valid0 ),
                .memc__dma__read_ready11        ( memc__dma__lane11_read_ready0      ),
                .dma__memc__read_pause11        ( dma__memc__lane11_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid12       ( dma__memc__lane12_write_valid0     ),
                .dma__memc__write_address12     ( dma__memc__lane12_write_address0   ),
                .dma__memc__write_data12        ( dma__memc__lane12_write_data0      ),
                .memc__dma__write_ready12       ( memc__dma__lane12_write_ready0     ),
                .dma__memc__read_valid12        ( dma__memc__lane12_read_valid0      ),
                .dma__memc__read_address12      ( dma__memc__lane12_read_address0    ),
                .memc__dma__read_data12         ( memc__dma__lane12_read_data0       ),
                .memc__dma__read_data_valid12   ( memc__dma__lane12_read_data_valid0 ),
                .memc__dma__read_ready12        ( memc__dma__lane12_read_ready0      ),
                .dma__memc__read_pause12        ( dma__memc__lane12_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid13       ( dma__memc__lane13_write_valid0     ),
                .dma__memc__write_address13     ( dma__memc__lane13_write_address0   ),
                .dma__memc__write_data13        ( dma__memc__lane13_write_data0      ),
                .memc__dma__write_ready13       ( memc__dma__lane13_write_ready0     ),
                .dma__memc__read_valid13        ( dma__memc__lane13_read_valid0      ),
                .dma__memc__read_address13      ( dma__memc__lane13_read_address0    ),
                .memc__dma__read_data13         ( memc__dma__lane13_read_data0       ),
                .memc__dma__read_data_valid13   ( memc__dma__lane13_read_data_valid0 ),
                .memc__dma__read_ready13        ( memc__dma__lane13_read_ready0      ),
                .dma__memc__read_pause13        ( dma__memc__lane13_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid14       ( dma__memc__lane14_write_valid0     ),
                .dma__memc__write_address14     ( dma__memc__lane14_write_address0   ),
                .dma__memc__write_data14        ( dma__memc__lane14_write_data0      ),
                .memc__dma__write_ready14       ( memc__dma__lane14_write_ready0     ),
                .dma__memc__read_valid14        ( dma__memc__lane14_read_valid0      ),
                .dma__memc__read_address14      ( dma__memc__lane14_read_address0    ),
                .memc__dma__read_data14         ( memc__dma__lane14_read_data0       ),
                .memc__dma__read_data_valid14   ( memc__dma__lane14_read_data_valid0 ),
                .memc__dma__read_ready14        ( memc__dma__lane14_read_ready0      ),
                .dma__memc__read_pause14        ( dma__memc__lane14_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid15       ( dma__memc__lane15_write_valid0     ),
                .dma__memc__write_address15     ( dma__memc__lane15_write_address0   ),
                .dma__memc__write_data15        ( dma__memc__lane15_write_data0      ),
                .memc__dma__write_ready15       ( memc__dma__lane15_write_ready0     ),
                .dma__memc__read_valid15        ( dma__memc__lane15_read_valid0      ),
                .dma__memc__read_address15      ( dma__memc__lane15_read_address0    ),
                .memc__dma__read_data15         ( memc__dma__lane15_read_data0       ),
                .memc__dma__read_data_valid15   ( memc__dma__lane15_read_data_valid0 ),
                .memc__dma__read_ready15        ( memc__dma__lane15_read_ready0      ),
                .dma__memc__read_pause15        ( dma__memc__lane15_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid16       ( dma__memc__lane16_write_valid0     ),
                .dma__memc__write_address16     ( dma__memc__lane16_write_address0   ),
                .dma__memc__write_data16        ( dma__memc__lane16_write_data0      ),
                .memc__dma__write_ready16       ( memc__dma__lane16_write_ready0     ),
                .dma__memc__read_valid16        ( dma__memc__lane16_read_valid0      ),
                .dma__memc__read_address16      ( dma__memc__lane16_read_address0    ),
                .memc__dma__read_data16         ( memc__dma__lane16_read_data0       ),
                .memc__dma__read_data_valid16   ( memc__dma__lane16_read_data_valid0 ),
                .memc__dma__read_ready16        ( memc__dma__lane16_read_ready0      ),
                .dma__memc__read_pause16        ( dma__memc__lane16_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid17       ( dma__memc__lane17_write_valid0     ),
                .dma__memc__write_address17     ( dma__memc__lane17_write_address0   ),
                .dma__memc__write_data17        ( dma__memc__lane17_write_data0      ),
                .memc__dma__write_ready17       ( memc__dma__lane17_write_ready0     ),
                .dma__memc__read_valid17        ( dma__memc__lane17_read_valid0      ),
                .dma__memc__read_address17      ( dma__memc__lane17_read_address0    ),
                .memc__dma__read_data17         ( memc__dma__lane17_read_data0       ),
                .memc__dma__read_data_valid17   ( memc__dma__lane17_read_data_valid0 ),
                .memc__dma__read_ready17        ( memc__dma__lane17_read_ready0      ),
                .dma__memc__read_pause17        ( dma__memc__lane17_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid18       ( dma__memc__lane18_write_valid0     ),
                .dma__memc__write_address18     ( dma__memc__lane18_write_address0   ),
                .dma__memc__write_data18        ( dma__memc__lane18_write_data0      ),
                .memc__dma__write_ready18       ( memc__dma__lane18_write_ready0     ),
                .dma__memc__read_valid18        ( dma__memc__lane18_read_valid0      ),
                .dma__memc__read_address18      ( dma__memc__lane18_read_address0    ),
                .memc__dma__read_data18         ( memc__dma__lane18_read_data0       ),
                .memc__dma__read_data_valid18   ( memc__dma__lane18_read_data_valid0 ),
                .memc__dma__read_ready18        ( memc__dma__lane18_read_ready0      ),
                .dma__memc__read_pause18        ( dma__memc__lane18_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid19       ( dma__memc__lane19_write_valid0     ),
                .dma__memc__write_address19     ( dma__memc__lane19_write_address0   ),
                .dma__memc__write_data19        ( dma__memc__lane19_write_data0      ),
                .memc__dma__write_ready19       ( memc__dma__lane19_write_ready0     ),
                .dma__memc__read_valid19        ( dma__memc__lane19_read_valid0      ),
                .dma__memc__read_address19      ( dma__memc__lane19_read_address0    ),
                .memc__dma__read_data19         ( memc__dma__lane19_read_data0       ),
                .memc__dma__read_data_valid19   ( memc__dma__lane19_read_data_valid0 ),
                .memc__dma__read_ready19        ( memc__dma__lane19_read_ready0      ),
                .dma__memc__read_pause19        ( dma__memc__lane19_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid20       ( dma__memc__lane20_write_valid0     ),
                .dma__memc__write_address20     ( dma__memc__lane20_write_address0   ),
                .dma__memc__write_data20        ( dma__memc__lane20_write_data0      ),
                .memc__dma__write_ready20       ( memc__dma__lane20_write_ready0     ),
                .dma__memc__read_valid20        ( dma__memc__lane20_read_valid0      ),
                .dma__memc__read_address20      ( dma__memc__lane20_read_address0    ),
                .memc__dma__read_data20         ( memc__dma__lane20_read_data0       ),
                .memc__dma__read_data_valid20   ( memc__dma__lane20_read_data_valid0 ),
                .memc__dma__read_ready20        ( memc__dma__lane20_read_ready0      ),
                .dma__memc__read_pause20        ( dma__memc__lane20_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid21       ( dma__memc__lane21_write_valid0     ),
                .dma__memc__write_address21     ( dma__memc__lane21_write_address0   ),
                .dma__memc__write_data21        ( dma__memc__lane21_write_data0      ),
                .memc__dma__write_ready21       ( memc__dma__lane21_write_ready0     ),
                .dma__memc__read_valid21        ( dma__memc__lane21_read_valid0      ),
                .dma__memc__read_address21      ( dma__memc__lane21_read_address0    ),
                .memc__dma__read_data21         ( memc__dma__lane21_read_data0       ),
                .memc__dma__read_data_valid21   ( memc__dma__lane21_read_data_valid0 ),
                .memc__dma__read_ready21        ( memc__dma__lane21_read_ready0      ),
                .dma__memc__read_pause21        ( dma__memc__lane21_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid22       ( dma__memc__lane22_write_valid0     ),
                .dma__memc__write_address22     ( dma__memc__lane22_write_address0   ),
                .dma__memc__write_data22        ( dma__memc__lane22_write_data0      ),
                .memc__dma__write_ready22       ( memc__dma__lane22_write_ready0     ),
                .dma__memc__read_valid22        ( dma__memc__lane22_read_valid0      ),
                .dma__memc__read_address22      ( dma__memc__lane22_read_address0    ),
                .memc__dma__read_data22         ( memc__dma__lane22_read_data0       ),
                .memc__dma__read_data_valid22   ( memc__dma__lane22_read_data_valid0 ),
                .memc__dma__read_ready22        ( memc__dma__lane22_read_ready0      ),
                .dma__memc__read_pause22        ( dma__memc__lane22_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid23       ( dma__memc__lane23_write_valid0     ),
                .dma__memc__write_address23     ( dma__memc__lane23_write_address0   ),
                .dma__memc__write_data23        ( dma__memc__lane23_write_data0      ),
                .memc__dma__write_ready23       ( memc__dma__lane23_write_ready0     ),
                .dma__memc__read_valid23        ( dma__memc__lane23_read_valid0      ),
                .dma__memc__read_address23      ( dma__memc__lane23_read_address0    ),
                .memc__dma__read_data23         ( memc__dma__lane23_read_data0       ),
                .memc__dma__read_data_valid23   ( memc__dma__lane23_read_data_valid0 ),
                .memc__dma__read_ready23        ( memc__dma__lane23_read_ready0      ),
                .dma__memc__read_pause23        ( dma__memc__lane23_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid24       ( dma__memc__lane24_write_valid0     ),
                .dma__memc__write_address24     ( dma__memc__lane24_write_address0   ),
                .dma__memc__write_data24        ( dma__memc__lane24_write_data0      ),
                .memc__dma__write_ready24       ( memc__dma__lane24_write_ready0     ),
                .dma__memc__read_valid24        ( dma__memc__lane24_read_valid0      ),
                .dma__memc__read_address24      ( dma__memc__lane24_read_address0    ),
                .memc__dma__read_data24         ( memc__dma__lane24_read_data0       ),
                .memc__dma__read_data_valid24   ( memc__dma__lane24_read_data_valid0 ),
                .memc__dma__read_ready24        ( memc__dma__lane24_read_ready0      ),
                .dma__memc__read_pause24        ( dma__memc__lane24_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid25       ( dma__memc__lane25_write_valid0     ),
                .dma__memc__write_address25     ( dma__memc__lane25_write_address0   ),
                .dma__memc__write_data25        ( dma__memc__lane25_write_data0      ),
                .memc__dma__write_ready25       ( memc__dma__lane25_write_ready0     ),
                .dma__memc__read_valid25        ( dma__memc__lane25_read_valid0      ),
                .dma__memc__read_address25      ( dma__memc__lane25_read_address0    ),
                .memc__dma__read_data25         ( memc__dma__lane25_read_data0       ),
                .memc__dma__read_data_valid25   ( memc__dma__lane25_read_data_valid0 ),
                .memc__dma__read_ready25        ( memc__dma__lane25_read_ready0      ),
                .dma__memc__read_pause25        ( dma__memc__lane25_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid26       ( dma__memc__lane26_write_valid0     ),
                .dma__memc__write_address26     ( dma__memc__lane26_write_address0   ),
                .dma__memc__write_data26        ( dma__memc__lane26_write_data0      ),
                .memc__dma__write_ready26       ( memc__dma__lane26_write_ready0     ),
                .dma__memc__read_valid26        ( dma__memc__lane26_read_valid0      ),
                .dma__memc__read_address26      ( dma__memc__lane26_read_address0    ),
                .memc__dma__read_data26         ( memc__dma__lane26_read_data0       ),
                .memc__dma__read_data_valid26   ( memc__dma__lane26_read_data_valid0 ),
                .memc__dma__read_ready26        ( memc__dma__lane26_read_ready0      ),
                .dma__memc__read_pause26        ( dma__memc__lane26_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid27       ( dma__memc__lane27_write_valid0     ),
                .dma__memc__write_address27     ( dma__memc__lane27_write_address0   ),
                .dma__memc__write_data27        ( dma__memc__lane27_write_data0      ),
                .memc__dma__write_ready27       ( memc__dma__lane27_write_ready0     ),
                .dma__memc__read_valid27        ( dma__memc__lane27_read_valid0      ),
                .dma__memc__read_address27      ( dma__memc__lane27_read_address0    ),
                .memc__dma__read_data27         ( memc__dma__lane27_read_data0       ),
                .memc__dma__read_data_valid27   ( memc__dma__lane27_read_data_valid0 ),
                .memc__dma__read_ready27        ( memc__dma__lane27_read_ready0      ),
                .dma__memc__read_pause27        ( dma__memc__lane27_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid28       ( dma__memc__lane28_write_valid0     ),
                .dma__memc__write_address28     ( dma__memc__lane28_write_address0   ),
                .dma__memc__write_data28        ( dma__memc__lane28_write_data0      ),
                .memc__dma__write_ready28       ( memc__dma__lane28_write_ready0     ),
                .dma__memc__read_valid28        ( dma__memc__lane28_read_valid0      ),
                .dma__memc__read_address28      ( dma__memc__lane28_read_address0    ),
                .memc__dma__read_data28         ( memc__dma__lane28_read_data0       ),
                .memc__dma__read_data_valid28   ( memc__dma__lane28_read_data_valid0 ),
                .memc__dma__read_ready28        ( memc__dma__lane28_read_ready0      ),
                .dma__memc__read_pause28        ( dma__memc__lane28_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid29       ( dma__memc__lane29_write_valid0     ),
                .dma__memc__write_address29     ( dma__memc__lane29_write_address0   ),
                .dma__memc__write_data29        ( dma__memc__lane29_write_data0      ),
                .memc__dma__write_ready29       ( memc__dma__lane29_write_ready0     ),
                .dma__memc__read_valid29        ( dma__memc__lane29_read_valid0      ),
                .dma__memc__read_address29      ( dma__memc__lane29_read_address0    ),
                .memc__dma__read_data29         ( memc__dma__lane29_read_data0       ),
                .memc__dma__read_data_valid29   ( memc__dma__lane29_read_data_valid0 ),
                .memc__dma__read_ready29        ( memc__dma__lane29_read_ready0      ),
                .dma__memc__read_pause29        ( dma__memc__lane29_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid30       ( dma__memc__lane30_write_valid0     ),
                .dma__memc__write_address30     ( dma__memc__lane30_write_address0   ),
                .dma__memc__write_data30        ( dma__memc__lane30_write_data0      ),
                .memc__dma__write_ready30       ( memc__dma__lane30_write_ready0     ),
                .dma__memc__read_valid30        ( dma__memc__lane30_read_valid0      ),
                .dma__memc__read_address30      ( dma__memc__lane30_read_address0    ),
                .memc__dma__read_data30         ( memc__dma__lane30_read_data0       ),
                .memc__dma__read_data_valid30   ( memc__dma__lane30_read_data_valid0 ),
                .memc__dma__read_ready30        ( memc__dma__lane30_read_ready0      ),
                .dma__memc__read_pause30        ( dma__memc__lane30_read_pause0      ),
                // Memory Port 0                 
                .dma__memc__write_valid31       ( dma__memc__lane31_write_valid0     ),
                .dma__memc__write_address31     ( dma__memc__lane31_write_address0   ),
                .dma__memc__write_data31        ( dma__memc__lane31_write_data0      ),
                .memc__dma__write_ready31       ( memc__dma__lane31_write_ready0     ),
                .dma__memc__read_valid31        ( dma__memc__lane31_read_valid0      ),
                .dma__memc__read_address31      ( dma__memc__lane31_read_address0    ),
                .memc__dma__read_data31         ( memc__dma__lane31_read_data0       ),
                .memc__dma__read_data_valid31   ( memc__dma__lane31_read_data_valid0 ),
                .memc__dma__read_ready31        ( memc__dma__lane31_read_ready0      ),
                .dma__memc__read_pause31        ( dma__memc__lane31_read_pause0      ),