`ifndef _dfi_vh
`define _dfi_vh

/*****************************************************************

    File name   : dfi.vh
    Author      : Lee Baker
    Affiliation : North Carolina State University, Raleigh, NC
    Date        : June 2017
    email       : lbbaker@ncsu.edu

      Note: leveraged from https://github.ncsu.edu/ECE-Memory-Controller-IS/ece-diram4-memory-controller/blob/master/HDL/run_s/dfi

*****************************************************************/


//---------------------------------------------------------------------------------------------------------------------



`endif
