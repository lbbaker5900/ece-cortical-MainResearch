
                  //----------------------------------------------------------------------------------------------------
                  // PE 0
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[0][0].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[0][0].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[0][0].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[0][0].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[0][0].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[0][0].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[0][0].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[0][0].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[0][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[0][0].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[0][1].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[0][1].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[0][1].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[0][1].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[0][1].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[0][1].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[0][1].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[0][1].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[0][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[0][1].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[0][2].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[0][2].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[0][2].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[0][2].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[0][2].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[0][2].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[0][2].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[0][2].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[0][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[0][2].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[0][3].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[0][3].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[0][3].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[0][3].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[0][3].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[0][3].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[0][3].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[0][3].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[0][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[0][3].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[0][4].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[0][4].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[0][4].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[0][4].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[0][4].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[0][4].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[0][4].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[0][4].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[0][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[0][4].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[0][5].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[0][5].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[0][5].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[0][5].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[0][5].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[0][5].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[0][5].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[0][5].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[0][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[0][5].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[0][6].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[0][6].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[0][6].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[0][6].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[0][6].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[0][6].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[0][6].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[0][6].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[0][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[0][6].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[0][7].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[0][7].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[0][7].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[0][7].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[0][7].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[0][7].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[0][7].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[0][7].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[0][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[0][7].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[0][8].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[0][8].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[0][8].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[0][8].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[0][8].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[0][8].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[0][8].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[0][8].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[0][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[0][8].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[0][9].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[0][9].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[0][9].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[0][9].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[0][9].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[0][9].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[0][9].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[0][9].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[0][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[0][9].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[0][10].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[0][10].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[0][10].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[0][10].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[0][10].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[0][10].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[0][10].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[0][10].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[0][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[0][10].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[0][11].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[0][11].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[0][11].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[0][11].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[0][11].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[0][11].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[0][11].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[0][11].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[0][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[0][11].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[0][12].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[0][12].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[0][12].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[0][12].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[0][12].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[0][12].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[0][12].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[0][12].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[0][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[0][12].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[0][13].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[0][13].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[0][13].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[0][13].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[0][13].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[0][13].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[0][13].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[0][13].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[0][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[0][13].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[0][14].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[0][14].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[0][14].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[0][14].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[0][14].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[0][14].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[0][14].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[0][14].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[0][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[0][14].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[0][15].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[0][15].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[0][15].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[0][15].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[0][15].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[0][15].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[0][15].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[0][15].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[0][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[0][15].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[0][16].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[0][16].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[0][16].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[0][16].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[0][16].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[0][16].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[0][16].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[0][16].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[0][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[0][16].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[0][17].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[0][17].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[0][17].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[0][17].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[0][17].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[0][17].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[0][17].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[0][17].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[0][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[0][17].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[0][18].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[0][18].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[0][18].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[0][18].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[0][18].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[0][18].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[0][18].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[0][18].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[0][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[0][18].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[0][19].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[0][19].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[0][19].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[0][19].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[0][19].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[0][19].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[0][19].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[0][19].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[0][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[0][19].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[0][20].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[0][20].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[0][20].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[0][20].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[0][20].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[0][20].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[0][20].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[0][20].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[0][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[0][20].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[0][21].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[0][21].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[0][21].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[0][21].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[0][21].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[0][21].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[0][21].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[0][21].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[0][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[0][21].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[0][22].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[0][22].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[0][22].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[0][22].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[0][22].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[0][22].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[0][22].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[0][22].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[0][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[0][22].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[0][23].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[0][23].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[0][23].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[0][23].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[0][23].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[0][23].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[0][23].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[0][23].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[0][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[0][23].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[0][24].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[0][24].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[0][24].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[0][24].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[0][24].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[0][24].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[0][24].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[0][24].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[0][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[0][24].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[0][25].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[0][25].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[0][25].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[0][25].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[0][25].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[0][25].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[0][25].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[0][25].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[0][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[0][25].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[0][26].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[0][26].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[0][26].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[0][26].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[0][26].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[0][26].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[0][26].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[0][26].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[0][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[0][26].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[0][27].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[0][27].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[0][27].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[0][27].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[0][27].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[0][27].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[0][27].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[0][27].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[0][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[0][27].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[0][28].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[0][28].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[0][28].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[0][28].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[0][28].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[0][28].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[0][28].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[0][28].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[0][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[0][28].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[0][29].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[0][29].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[0][29].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[0][29].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[0][29].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[0][29].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[0][29].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[0][29].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[0][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[0][29].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[0][30].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[0][30].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[0][30].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[0][30].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[0][30].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[0][30].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[0][30].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[0][30].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[0][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[0][30].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[0][31].dma__memc__write_valid      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[0][31].dma__memc__write_address    = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[0][31].dma__memc__write_data       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[0][31].dma__memc__read_valid       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[0][31].dma__memc__read_address     = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[0][31].dma__memc__read_pause       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[0][31].memc__dma__write_ready      = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[0][31].memc__dma__read_data        = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[0][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[0][31].memc__dma__read_ready       = pe_array_inst.pe_inst[0].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 1
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[1][0].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[1][0].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[1][0].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[1][0].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[1][0].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[1][0].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[1][0].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[1][0].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[1][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[1][0].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[1][1].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[1][1].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[1][1].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[1][1].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[1][1].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[1][1].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[1][1].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[1][1].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[1][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[1][1].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[1][2].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[1][2].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[1][2].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[1][2].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[1][2].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[1][2].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[1][2].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[1][2].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[1][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[1][2].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[1][3].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[1][3].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[1][3].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[1][3].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[1][3].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[1][3].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[1][3].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[1][3].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[1][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[1][3].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[1][4].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[1][4].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[1][4].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[1][4].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[1][4].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[1][4].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[1][4].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[1][4].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[1][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[1][4].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[1][5].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[1][5].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[1][5].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[1][5].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[1][5].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[1][5].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[1][5].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[1][5].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[1][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[1][5].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[1][6].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[1][6].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[1][6].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[1][6].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[1][6].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[1][6].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[1][6].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[1][6].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[1][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[1][6].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[1][7].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[1][7].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[1][7].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[1][7].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[1][7].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[1][7].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[1][7].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[1][7].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[1][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[1][7].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[1][8].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[1][8].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[1][8].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[1][8].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[1][8].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[1][8].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[1][8].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[1][8].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[1][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[1][8].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[1][9].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[1][9].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[1][9].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[1][9].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[1][9].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[1][9].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[1][9].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[1][9].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[1][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[1][9].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[1][10].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[1][10].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[1][10].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[1][10].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[1][10].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[1][10].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[1][10].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[1][10].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[1][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[1][10].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[1][11].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[1][11].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[1][11].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[1][11].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[1][11].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[1][11].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[1][11].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[1][11].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[1][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[1][11].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[1][12].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[1][12].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[1][12].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[1][12].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[1][12].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[1][12].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[1][12].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[1][12].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[1][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[1][12].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[1][13].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[1][13].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[1][13].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[1][13].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[1][13].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[1][13].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[1][13].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[1][13].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[1][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[1][13].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[1][14].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[1][14].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[1][14].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[1][14].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[1][14].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[1][14].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[1][14].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[1][14].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[1][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[1][14].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[1][15].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[1][15].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[1][15].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[1][15].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[1][15].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[1][15].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[1][15].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[1][15].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[1][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[1][15].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[1][16].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[1][16].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[1][16].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[1][16].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[1][16].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[1][16].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[1][16].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[1][16].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[1][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[1][16].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[1][17].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[1][17].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[1][17].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[1][17].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[1][17].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[1][17].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[1][17].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[1][17].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[1][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[1][17].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[1][18].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[1][18].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[1][18].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[1][18].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[1][18].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[1][18].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[1][18].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[1][18].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[1][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[1][18].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[1][19].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[1][19].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[1][19].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[1][19].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[1][19].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[1][19].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[1][19].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[1][19].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[1][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[1][19].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[1][20].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[1][20].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[1][20].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[1][20].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[1][20].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[1][20].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[1][20].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[1][20].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[1][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[1][20].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[1][21].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[1][21].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[1][21].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[1][21].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[1][21].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[1][21].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[1][21].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[1][21].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[1][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[1][21].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[1][22].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[1][22].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[1][22].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[1][22].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[1][22].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[1][22].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[1][22].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[1][22].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[1][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[1][22].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[1][23].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[1][23].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[1][23].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[1][23].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[1][23].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[1][23].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[1][23].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[1][23].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[1][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[1][23].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[1][24].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[1][24].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[1][24].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[1][24].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[1][24].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[1][24].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[1][24].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[1][24].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[1][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[1][24].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[1][25].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[1][25].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[1][25].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[1][25].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[1][25].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[1][25].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[1][25].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[1][25].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[1][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[1][25].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[1][26].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[1][26].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[1][26].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[1][26].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[1][26].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[1][26].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[1][26].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[1][26].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[1][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[1][26].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[1][27].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[1][27].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[1][27].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[1][27].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[1][27].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[1][27].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[1][27].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[1][27].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[1][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[1][27].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[1][28].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[1][28].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[1][28].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[1][28].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[1][28].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[1][28].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[1][28].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[1][28].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[1][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[1][28].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[1][29].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[1][29].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[1][29].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[1][29].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[1][29].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[1][29].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[1][29].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[1][29].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[1][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[1][29].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[1][30].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[1][30].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[1][30].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[1][30].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[1][30].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[1][30].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[1][30].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[1][30].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[1][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[1][30].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[1][31].dma__memc__write_valid      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[1][31].dma__memc__write_address    = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[1][31].dma__memc__write_data       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[1][31].dma__memc__read_valid       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[1][31].dma__memc__read_address     = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[1][31].dma__memc__read_pause       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[1][31].memc__dma__write_ready      = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[1][31].memc__dma__read_data        = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[1][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[1][31].memc__dma__read_ready       = pe_array_inst.pe_inst[1].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 2
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[2][0].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[2][0].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[2][0].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[2][0].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[2][0].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[2][0].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[2][0].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[2][0].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[2][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[2][0].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[2][1].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[2][1].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[2][1].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[2][1].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[2][1].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[2][1].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[2][1].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[2][1].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[2][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[2][1].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[2][2].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[2][2].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[2][2].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[2][2].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[2][2].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[2][2].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[2][2].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[2][2].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[2][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[2][2].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[2][3].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[2][3].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[2][3].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[2][3].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[2][3].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[2][3].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[2][3].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[2][3].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[2][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[2][3].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[2][4].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[2][4].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[2][4].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[2][4].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[2][4].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[2][4].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[2][4].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[2][4].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[2][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[2][4].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[2][5].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[2][5].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[2][5].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[2][5].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[2][5].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[2][5].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[2][5].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[2][5].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[2][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[2][5].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[2][6].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[2][6].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[2][6].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[2][6].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[2][6].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[2][6].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[2][6].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[2][6].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[2][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[2][6].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[2][7].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[2][7].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[2][7].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[2][7].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[2][7].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[2][7].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[2][7].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[2][7].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[2][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[2][7].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[2][8].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[2][8].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[2][8].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[2][8].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[2][8].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[2][8].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[2][8].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[2][8].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[2][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[2][8].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[2][9].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[2][9].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[2][9].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[2][9].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[2][9].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[2][9].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[2][9].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[2][9].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[2][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[2][9].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[2][10].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[2][10].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[2][10].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[2][10].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[2][10].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[2][10].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[2][10].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[2][10].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[2][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[2][10].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[2][11].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[2][11].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[2][11].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[2][11].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[2][11].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[2][11].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[2][11].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[2][11].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[2][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[2][11].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[2][12].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[2][12].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[2][12].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[2][12].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[2][12].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[2][12].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[2][12].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[2][12].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[2][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[2][12].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[2][13].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[2][13].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[2][13].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[2][13].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[2][13].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[2][13].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[2][13].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[2][13].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[2][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[2][13].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[2][14].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[2][14].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[2][14].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[2][14].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[2][14].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[2][14].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[2][14].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[2][14].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[2][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[2][14].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[2][15].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[2][15].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[2][15].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[2][15].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[2][15].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[2][15].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[2][15].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[2][15].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[2][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[2][15].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[2][16].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[2][16].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[2][16].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[2][16].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[2][16].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[2][16].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[2][16].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[2][16].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[2][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[2][16].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[2][17].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[2][17].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[2][17].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[2][17].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[2][17].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[2][17].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[2][17].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[2][17].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[2][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[2][17].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[2][18].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[2][18].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[2][18].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[2][18].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[2][18].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[2][18].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[2][18].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[2][18].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[2][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[2][18].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[2][19].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[2][19].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[2][19].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[2][19].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[2][19].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[2][19].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[2][19].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[2][19].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[2][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[2][19].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[2][20].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[2][20].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[2][20].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[2][20].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[2][20].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[2][20].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[2][20].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[2][20].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[2][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[2][20].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[2][21].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[2][21].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[2][21].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[2][21].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[2][21].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[2][21].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[2][21].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[2][21].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[2][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[2][21].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[2][22].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[2][22].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[2][22].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[2][22].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[2][22].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[2][22].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[2][22].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[2][22].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[2][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[2][22].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[2][23].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[2][23].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[2][23].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[2][23].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[2][23].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[2][23].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[2][23].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[2][23].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[2][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[2][23].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[2][24].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[2][24].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[2][24].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[2][24].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[2][24].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[2][24].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[2][24].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[2][24].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[2][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[2][24].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[2][25].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[2][25].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[2][25].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[2][25].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[2][25].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[2][25].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[2][25].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[2][25].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[2][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[2][25].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[2][26].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[2][26].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[2][26].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[2][26].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[2][26].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[2][26].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[2][26].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[2][26].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[2][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[2][26].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[2][27].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[2][27].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[2][27].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[2][27].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[2][27].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[2][27].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[2][27].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[2][27].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[2][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[2][27].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[2][28].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[2][28].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[2][28].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[2][28].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[2][28].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[2][28].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[2][28].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[2][28].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[2][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[2][28].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[2][29].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[2][29].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[2][29].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[2][29].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[2][29].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[2][29].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[2][29].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[2][29].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[2][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[2][29].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[2][30].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[2][30].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[2][30].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[2][30].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[2][30].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[2][30].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[2][30].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[2][30].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[2][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[2][30].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[2][31].dma__memc__write_valid      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[2][31].dma__memc__write_address    = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[2][31].dma__memc__write_data       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[2][31].dma__memc__read_valid       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[2][31].dma__memc__read_address     = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[2][31].dma__memc__read_pause       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[2][31].memc__dma__write_ready      = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[2][31].memc__dma__read_data        = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[2][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[2][31].memc__dma__read_ready       = pe_array_inst.pe_inst[2].pe.mem_acc_cont.memc__dma__read_ready31         ;

                  //----------------------------------------------------------------------------------------------------
                  // PE 3
                  // 
                  //--------------------------------------------------
                  // Lane 0
                  assign Dma2Mem[3][0].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid0        ;
                  assign Dma2Mem[3][0].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address0      ;
                  assign Dma2Mem[3][0].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data0         ;
                  assign Dma2Mem[3][0].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid0         ;
                  assign Dma2Mem[3][0].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address0       ;
                  assign Dma2Mem[3][0].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause0         ;

                  assign Dma2Mem[3][0].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready0        ;
                  assign Dma2Mem[3][0].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data0          ;
                  assign Dma2Mem[3][0].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid0    ;
                  assign Dma2Mem[3][0].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready0         ;

                  //--------------------------------------------------
                  // Lane 1
                  assign Dma2Mem[3][1].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid1        ;
                  assign Dma2Mem[3][1].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address1      ;
                  assign Dma2Mem[3][1].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data1         ;
                  assign Dma2Mem[3][1].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid1         ;
                  assign Dma2Mem[3][1].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address1       ;
                  assign Dma2Mem[3][1].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause1         ;

                  assign Dma2Mem[3][1].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready1        ;
                  assign Dma2Mem[3][1].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data1          ;
                  assign Dma2Mem[3][1].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid1    ;
                  assign Dma2Mem[3][1].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready1         ;

                  //--------------------------------------------------
                  // Lane 2
                  assign Dma2Mem[3][2].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid2        ;
                  assign Dma2Mem[3][2].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address2      ;
                  assign Dma2Mem[3][2].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data2         ;
                  assign Dma2Mem[3][2].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid2         ;
                  assign Dma2Mem[3][2].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address2       ;
                  assign Dma2Mem[3][2].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause2         ;

                  assign Dma2Mem[3][2].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready2        ;
                  assign Dma2Mem[3][2].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data2          ;
                  assign Dma2Mem[3][2].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid2    ;
                  assign Dma2Mem[3][2].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready2         ;

                  //--------------------------------------------------
                  // Lane 3
                  assign Dma2Mem[3][3].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid3        ;
                  assign Dma2Mem[3][3].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address3      ;
                  assign Dma2Mem[3][3].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data3         ;
                  assign Dma2Mem[3][3].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid3         ;
                  assign Dma2Mem[3][3].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address3       ;
                  assign Dma2Mem[3][3].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause3         ;

                  assign Dma2Mem[3][3].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready3        ;
                  assign Dma2Mem[3][3].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data3          ;
                  assign Dma2Mem[3][3].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid3    ;
                  assign Dma2Mem[3][3].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready3         ;

                  //--------------------------------------------------
                  // Lane 4
                  assign Dma2Mem[3][4].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid4        ;
                  assign Dma2Mem[3][4].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address4      ;
                  assign Dma2Mem[3][4].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data4         ;
                  assign Dma2Mem[3][4].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid4         ;
                  assign Dma2Mem[3][4].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address4       ;
                  assign Dma2Mem[3][4].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause4         ;

                  assign Dma2Mem[3][4].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready4        ;
                  assign Dma2Mem[3][4].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data4          ;
                  assign Dma2Mem[3][4].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid4    ;
                  assign Dma2Mem[3][4].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready4         ;

                  //--------------------------------------------------
                  // Lane 5
                  assign Dma2Mem[3][5].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid5        ;
                  assign Dma2Mem[3][5].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address5      ;
                  assign Dma2Mem[3][5].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data5         ;
                  assign Dma2Mem[3][5].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid5         ;
                  assign Dma2Mem[3][5].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address5       ;
                  assign Dma2Mem[3][5].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause5         ;

                  assign Dma2Mem[3][5].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready5        ;
                  assign Dma2Mem[3][5].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data5          ;
                  assign Dma2Mem[3][5].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid5    ;
                  assign Dma2Mem[3][5].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready5         ;

                  //--------------------------------------------------
                  // Lane 6
                  assign Dma2Mem[3][6].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid6        ;
                  assign Dma2Mem[3][6].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address6      ;
                  assign Dma2Mem[3][6].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data6         ;
                  assign Dma2Mem[3][6].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid6         ;
                  assign Dma2Mem[3][6].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address6       ;
                  assign Dma2Mem[3][6].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause6         ;

                  assign Dma2Mem[3][6].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready6        ;
                  assign Dma2Mem[3][6].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data6          ;
                  assign Dma2Mem[3][6].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid6    ;
                  assign Dma2Mem[3][6].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready6         ;

                  //--------------------------------------------------
                  // Lane 7
                  assign Dma2Mem[3][7].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid7        ;
                  assign Dma2Mem[3][7].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address7      ;
                  assign Dma2Mem[3][7].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data7         ;
                  assign Dma2Mem[3][7].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid7         ;
                  assign Dma2Mem[3][7].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address7       ;
                  assign Dma2Mem[3][7].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause7         ;

                  assign Dma2Mem[3][7].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready7        ;
                  assign Dma2Mem[3][7].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data7          ;
                  assign Dma2Mem[3][7].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid7    ;
                  assign Dma2Mem[3][7].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready7         ;

                  //--------------------------------------------------
                  // Lane 8
                  assign Dma2Mem[3][8].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid8        ;
                  assign Dma2Mem[3][8].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address8      ;
                  assign Dma2Mem[3][8].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data8         ;
                  assign Dma2Mem[3][8].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid8         ;
                  assign Dma2Mem[3][8].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address8       ;
                  assign Dma2Mem[3][8].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause8         ;

                  assign Dma2Mem[3][8].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready8        ;
                  assign Dma2Mem[3][8].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data8          ;
                  assign Dma2Mem[3][8].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid8    ;
                  assign Dma2Mem[3][8].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready8         ;

                  //--------------------------------------------------
                  // Lane 9
                  assign Dma2Mem[3][9].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid9        ;
                  assign Dma2Mem[3][9].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address9      ;
                  assign Dma2Mem[3][9].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data9         ;
                  assign Dma2Mem[3][9].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid9         ;
                  assign Dma2Mem[3][9].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address9       ;
                  assign Dma2Mem[3][9].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause9         ;

                  assign Dma2Mem[3][9].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready9        ;
                  assign Dma2Mem[3][9].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data9          ;
                  assign Dma2Mem[3][9].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid9    ;
                  assign Dma2Mem[3][9].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready9         ;

                  //--------------------------------------------------
                  // Lane 10
                  assign Dma2Mem[3][10].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid10        ;
                  assign Dma2Mem[3][10].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address10      ;
                  assign Dma2Mem[3][10].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data10         ;
                  assign Dma2Mem[3][10].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid10         ;
                  assign Dma2Mem[3][10].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address10       ;
                  assign Dma2Mem[3][10].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause10         ;

                  assign Dma2Mem[3][10].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready10        ;
                  assign Dma2Mem[3][10].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data10          ;
                  assign Dma2Mem[3][10].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid10    ;
                  assign Dma2Mem[3][10].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready10         ;

                  //--------------------------------------------------
                  // Lane 11
                  assign Dma2Mem[3][11].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid11        ;
                  assign Dma2Mem[3][11].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address11      ;
                  assign Dma2Mem[3][11].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data11         ;
                  assign Dma2Mem[3][11].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid11         ;
                  assign Dma2Mem[3][11].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address11       ;
                  assign Dma2Mem[3][11].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause11         ;

                  assign Dma2Mem[3][11].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready11        ;
                  assign Dma2Mem[3][11].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data11          ;
                  assign Dma2Mem[3][11].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid11    ;
                  assign Dma2Mem[3][11].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready11         ;

                  //--------------------------------------------------
                  // Lane 12
                  assign Dma2Mem[3][12].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid12        ;
                  assign Dma2Mem[3][12].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address12      ;
                  assign Dma2Mem[3][12].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data12         ;
                  assign Dma2Mem[3][12].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid12         ;
                  assign Dma2Mem[3][12].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address12       ;
                  assign Dma2Mem[3][12].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause12         ;

                  assign Dma2Mem[3][12].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready12        ;
                  assign Dma2Mem[3][12].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data12          ;
                  assign Dma2Mem[3][12].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid12    ;
                  assign Dma2Mem[3][12].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready12         ;

                  //--------------------------------------------------
                  // Lane 13
                  assign Dma2Mem[3][13].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid13        ;
                  assign Dma2Mem[3][13].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address13      ;
                  assign Dma2Mem[3][13].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data13         ;
                  assign Dma2Mem[3][13].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid13         ;
                  assign Dma2Mem[3][13].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address13       ;
                  assign Dma2Mem[3][13].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause13         ;

                  assign Dma2Mem[3][13].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready13        ;
                  assign Dma2Mem[3][13].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data13          ;
                  assign Dma2Mem[3][13].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid13    ;
                  assign Dma2Mem[3][13].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready13         ;

                  //--------------------------------------------------
                  // Lane 14
                  assign Dma2Mem[3][14].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid14        ;
                  assign Dma2Mem[3][14].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address14      ;
                  assign Dma2Mem[3][14].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data14         ;
                  assign Dma2Mem[3][14].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid14         ;
                  assign Dma2Mem[3][14].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address14       ;
                  assign Dma2Mem[3][14].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause14         ;

                  assign Dma2Mem[3][14].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready14        ;
                  assign Dma2Mem[3][14].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data14          ;
                  assign Dma2Mem[3][14].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid14    ;
                  assign Dma2Mem[3][14].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready14         ;

                  //--------------------------------------------------
                  // Lane 15
                  assign Dma2Mem[3][15].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid15        ;
                  assign Dma2Mem[3][15].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address15      ;
                  assign Dma2Mem[3][15].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data15         ;
                  assign Dma2Mem[3][15].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid15         ;
                  assign Dma2Mem[3][15].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address15       ;
                  assign Dma2Mem[3][15].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause15         ;

                  assign Dma2Mem[3][15].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready15        ;
                  assign Dma2Mem[3][15].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data15          ;
                  assign Dma2Mem[3][15].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid15    ;
                  assign Dma2Mem[3][15].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready15         ;

                  //--------------------------------------------------
                  // Lane 16
                  assign Dma2Mem[3][16].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid16        ;
                  assign Dma2Mem[3][16].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address16      ;
                  assign Dma2Mem[3][16].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data16         ;
                  assign Dma2Mem[3][16].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid16         ;
                  assign Dma2Mem[3][16].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address16       ;
                  assign Dma2Mem[3][16].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause16         ;

                  assign Dma2Mem[3][16].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready16        ;
                  assign Dma2Mem[3][16].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data16          ;
                  assign Dma2Mem[3][16].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid16    ;
                  assign Dma2Mem[3][16].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready16         ;

                  //--------------------------------------------------
                  // Lane 17
                  assign Dma2Mem[3][17].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid17        ;
                  assign Dma2Mem[3][17].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address17      ;
                  assign Dma2Mem[3][17].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data17         ;
                  assign Dma2Mem[3][17].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid17         ;
                  assign Dma2Mem[3][17].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address17       ;
                  assign Dma2Mem[3][17].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause17         ;

                  assign Dma2Mem[3][17].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready17        ;
                  assign Dma2Mem[3][17].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data17          ;
                  assign Dma2Mem[3][17].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid17    ;
                  assign Dma2Mem[3][17].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready17         ;

                  //--------------------------------------------------
                  // Lane 18
                  assign Dma2Mem[3][18].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid18        ;
                  assign Dma2Mem[3][18].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address18      ;
                  assign Dma2Mem[3][18].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data18         ;
                  assign Dma2Mem[3][18].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid18         ;
                  assign Dma2Mem[3][18].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address18       ;
                  assign Dma2Mem[3][18].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause18         ;

                  assign Dma2Mem[3][18].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready18        ;
                  assign Dma2Mem[3][18].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data18          ;
                  assign Dma2Mem[3][18].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid18    ;
                  assign Dma2Mem[3][18].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready18         ;

                  //--------------------------------------------------
                  // Lane 19
                  assign Dma2Mem[3][19].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid19        ;
                  assign Dma2Mem[3][19].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address19      ;
                  assign Dma2Mem[3][19].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data19         ;
                  assign Dma2Mem[3][19].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid19         ;
                  assign Dma2Mem[3][19].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address19       ;
                  assign Dma2Mem[3][19].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause19         ;

                  assign Dma2Mem[3][19].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready19        ;
                  assign Dma2Mem[3][19].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data19          ;
                  assign Dma2Mem[3][19].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid19    ;
                  assign Dma2Mem[3][19].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready19         ;

                  //--------------------------------------------------
                  // Lane 20
                  assign Dma2Mem[3][20].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid20        ;
                  assign Dma2Mem[3][20].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address20      ;
                  assign Dma2Mem[3][20].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data20         ;
                  assign Dma2Mem[3][20].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid20         ;
                  assign Dma2Mem[3][20].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address20       ;
                  assign Dma2Mem[3][20].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause20         ;

                  assign Dma2Mem[3][20].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready20        ;
                  assign Dma2Mem[3][20].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data20          ;
                  assign Dma2Mem[3][20].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid20    ;
                  assign Dma2Mem[3][20].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready20         ;

                  //--------------------------------------------------
                  // Lane 21
                  assign Dma2Mem[3][21].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid21        ;
                  assign Dma2Mem[3][21].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address21      ;
                  assign Dma2Mem[3][21].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data21         ;
                  assign Dma2Mem[3][21].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid21         ;
                  assign Dma2Mem[3][21].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address21       ;
                  assign Dma2Mem[3][21].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause21         ;

                  assign Dma2Mem[3][21].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready21        ;
                  assign Dma2Mem[3][21].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data21          ;
                  assign Dma2Mem[3][21].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid21    ;
                  assign Dma2Mem[3][21].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready21         ;

                  //--------------------------------------------------
                  // Lane 22
                  assign Dma2Mem[3][22].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid22        ;
                  assign Dma2Mem[3][22].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address22      ;
                  assign Dma2Mem[3][22].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data22         ;
                  assign Dma2Mem[3][22].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid22         ;
                  assign Dma2Mem[3][22].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address22       ;
                  assign Dma2Mem[3][22].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause22         ;

                  assign Dma2Mem[3][22].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready22        ;
                  assign Dma2Mem[3][22].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data22          ;
                  assign Dma2Mem[3][22].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid22    ;
                  assign Dma2Mem[3][22].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready22         ;

                  //--------------------------------------------------
                  // Lane 23
                  assign Dma2Mem[3][23].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid23        ;
                  assign Dma2Mem[3][23].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address23      ;
                  assign Dma2Mem[3][23].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data23         ;
                  assign Dma2Mem[3][23].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid23         ;
                  assign Dma2Mem[3][23].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address23       ;
                  assign Dma2Mem[3][23].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause23         ;

                  assign Dma2Mem[3][23].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready23        ;
                  assign Dma2Mem[3][23].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data23          ;
                  assign Dma2Mem[3][23].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid23    ;
                  assign Dma2Mem[3][23].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready23         ;

                  //--------------------------------------------------
                  // Lane 24
                  assign Dma2Mem[3][24].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid24        ;
                  assign Dma2Mem[3][24].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address24      ;
                  assign Dma2Mem[3][24].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data24         ;
                  assign Dma2Mem[3][24].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid24         ;
                  assign Dma2Mem[3][24].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address24       ;
                  assign Dma2Mem[3][24].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause24         ;

                  assign Dma2Mem[3][24].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready24        ;
                  assign Dma2Mem[3][24].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data24          ;
                  assign Dma2Mem[3][24].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid24    ;
                  assign Dma2Mem[3][24].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready24         ;

                  //--------------------------------------------------
                  // Lane 25
                  assign Dma2Mem[3][25].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid25        ;
                  assign Dma2Mem[3][25].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address25      ;
                  assign Dma2Mem[3][25].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data25         ;
                  assign Dma2Mem[3][25].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid25         ;
                  assign Dma2Mem[3][25].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address25       ;
                  assign Dma2Mem[3][25].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause25         ;

                  assign Dma2Mem[3][25].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready25        ;
                  assign Dma2Mem[3][25].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data25          ;
                  assign Dma2Mem[3][25].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid25    ;
                  assign Dma2Mem[3][25].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready25         ;

                  //--------------------------------------------------
                  // Lane 26
                  assign Dma2Mem[3][26].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid26        ;
                  assign Dma2Mem[3][26].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address26      ;
                  assign Dma2Mem[3][26].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data26         ;
                  assign Dma2Mem[3][26].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid26         ;
                  assign Dma2Mem[3][26].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address26       ;
                  assign Dma2Mem[3][26].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause26         ;

                  assign Dma2Mem[3][26].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready26        ;
                  assign Dma2Mem[3][26].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data26          ;
                  assign Dma2Mem[3][26].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid26    ;
                  assign Dma2Mem[3][26].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready26         ;

                  //--------------------------------------------------
                  // Lane 27
                  assign Dma2Mem[3][27].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid27        ;
                  assign Dma2Mem[3][27].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address27      ;
                  assign Dma2Mem[3][27].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data27         ;
                  assign Dma2Mem[3][27].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid27         ;
                  assign Dma2Mem[3][27].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address27       ;
                  assign Dma2Mem[3][27].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause27         ;

                  assign Dma2Mem[3][27].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready27        ;
                  assign Dma2Mem[3][27].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data27          ;
                  assign Dma2Mem[3][27].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid27    ;
                  assign Dma2Mem[3][27].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready27         ;

                  //--------------------------------------------------
                  // Lane 28
                  assign Dma2Mem[3][28].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid28        ;
                  assign Dma2Mem[3][28].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address28      ;
                  assign Dma2Mem[3][28].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data28         ;
                  assign Dma2Mem[3][28].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid28         ;
                  assign Dma2Mem[3][28].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address28       ;
                  assign Dma2Mem[3][28].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause28         ;

                  assign Dma2Mem[3][28].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready28        ;
                  assign Dma2Mem[3][28].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data28          ;
                  assign Dma2Mem[3][28].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid28    ;
                  assign Dma2Mem[3][28].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready28         ;

                  //--------------------------------------------------
                  // Lane 29
                  assign Dma2Mem[3][29].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid29        ;
                  assign Dma2Mem[3][29].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address29      ;
                  assign Dma2Mem[3][29].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data29         ;
                  assign Dma2Mem[3][29].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid29         ;
                  assign Dma2Mem[3][29].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address29       ;
                  assign Dma2Mem[3][29].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause29         ;

                  assign Dma2Mem[3][29].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready29        ;
                  assign Dma2Mem[3][29].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data29          ;
                  assign Dma2Mem[3][29].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid29    ;
                  assign Dma2Mem[3][29].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready29         ;

                  //--------------------------------------------------
                  // Lane 30
                  assign Dma2Mem[3][30].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid30        ;
                  assign Dma2Mem[3][30].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address30      ;
                  assign Dma2Mem[3][30].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data30         ;
                  assign Dma2Mem[3][30].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid30         ;
                  assign Dma2Mem[3][30].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address30       ;
                  assign Dma2Mem[3][30].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause30         ;

                  assign Dma2Mem[3][30].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready30        ;
                  assign Dma2Mem[3][30].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data30          ;
                  assign Dma2Mem[3][30].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid30    ;
                  assign Dma2Mem[3][30].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready30         ;

                  //--------------------------------------------------
                  // Lane 31
                  assign Dma2Mem[3][31].dma__memc__write_valid      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_valid31        ;
                  assign Dma2Mem[3][31].dma__memc__write_address    = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_address31      ;
                  assign Dma2Mem[3][31].dma__memc__write_data       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__write_data31         ;
                  assign Dma2Mem[3][31].dma__memc__read_valid       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_valid31         ;
                  assign Dma2Mem[3][31].dma__memc__read_address     = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_address31       ;
                  assign Dma2Mem[3][31].dma__memc__read_pause       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.dma__memc__read_pause31         ;

                  assign Dma2Mem[3][31].memc__dma__write_ready      = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__write_ready31        ;
                  assign Dma2Mem[3][31].memc__dma__read_data        = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data31          ;
                  assign Dma2Mem[3][31].memc__dma__read_data_valid  = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_data_valid31    ;
                  assign Dma2Mem[3][31].memc__dma__read_ready       = pe_array_inst.pe_inst[3].pe.mem_acc_cont.memc__dma__read_ready31         ;
