
  // NoC port 0
  output                                   pe__noc__port0_valid           ;
  output [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port0_cntl            ;
  output [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port0_data            ;
  input                                    noc__pe__port0_fc              ;
  input                                    noc__pe__port0_valid           ;
  input  [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port0_cntl            ;
  input  [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port0_data            ;
  output                                   pe__noc__port0_fc              ;
  input  [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port0_destinationMask ;

  // NoC port 1
  output                                   pe__noc__port1_valid           ;
  output [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port1_cntl            ;
  output [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port1_data            ;
  input                                    noc__pe__port1_fc              ;
  input                                    noc__pe__port1_valid           ;
  input  [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port1_cntl            ;
  input  [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port1_data            ;
  output                                   pe__noc__port1_fc              ;
  input  [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port1_destinationMask ;

  // NoC port 2
  output                                   pe__noc__port2_valid           ;
  output [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port2_cntl            ;
  output [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port2_data            ;
  input                                    noc__pe__port2_fc              ;
  input                                    noc__pe__port2_valid           ;
  input  [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port2_cntl            ;
  input  [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port2_data            ;
  output                                   pe__noc__port2_fc              ;
  input  [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port2_destinationMask ;

  // NoC port 3
  output                                   pe__noc__port3_valid           ;
  output [`COMMON_STD_INTF_CNTL_RANGE ]  pe__noc__port3_cntl            ;
  output [`NOC_CONT_NOC_PORT_DATA_RANGE ]  pe__noc__port3_data            ;
  input                                    noc__pe__port3_fc              ;
  input                                    noc__pe__port3_valid           ;
  input  [`COMMON_STD_INTF_CNTL_RANGE ]  noc__pe__port3_cntl            ;
  input  [`NOC_CONT_NOC_PORT_DATA_RANGE ]  noc__pe__port3_data            ;
  output                                   pe__noc__port3_fc              ;
  input  [`PE_PE_ID_BITMASK_RANGE       ]  sys__pe__port3_destinationMask ;

