
            // NoC port 0
            pe__noc__port0_valid            ,
            pe__noc__port0_cntl             ,
            pe__noc__port0_data             ,
            noc__pe__port0_fc               ,
            noc__pe__port0_valid            ,
            noc__pe__port0_cntl             ,
            noc__pe__port0_data             ,
            pe__noc__port0_fc               ,
            sys__pe__port0_destinationMask  ,

            // NoC port 1
            pe__noc__port1_valid            ,
            pe__noc__port1_cntl             ,
            pe__noc__port1_data             ,
            noc__pe__port1_fc               ,
            noc__pe__port1_valid            ,
            noc__pe__port1_cntl             ,
            noc__pe__port1_data             ,
            pe__noc__port1_fc               ,
            sys__pe__port1_destinationMask  ,

            // NoC port 2
            pe__noc__port2_valid            ,
            pe__noc__port2_cntl             ,
            pe__noc__port2_data             ,
            noc__pe__port2_fc               ,
            noc__pe__port2_valid            ,
            noc__pe__port2_cntl             ,
            noc__pe__port2_data             ,
            pe__noc__port2_fc               ,
            sys__pe__port2_destinationMask  ,

            // NoC port 3
            pe__noc__port3_valid            ,
            pe__noc__port3_cntl             ,
            pe__noc__port3_data             ,
            noc__pe__port3_fc               ,
            noc__pe__port3_valid            ,
            noc__pe__port3_cntl             ,
            noc__pe__port3_data             ,
            pe__noc__port3_fc               ,
            sys__pe__port3_destinationMask  ,

